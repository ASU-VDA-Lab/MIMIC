module fake_netlist_5_45_n_4086 (n_137, n_294, n_431, n_318, n_380, n_419, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_422, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_420, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_4086);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_422;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_4086;

wire n_924;
wire n_1263;
wire n_3304;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_2771;
wire n_785;
wire n_3241;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3863;
wire n_3795;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_3906;
wire n_880;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_3641;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4038;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_3445;
wire n_447;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_625;
wire n_854;
wire n_1462;
wire n_2069;
wire n_2396;
wire n_1799;
wire n_3621;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4033;
wire n_877;
wire n_2538;
wire n_2105;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_556;
wire n_3036;
wire n_2482;
wire n_3891;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4061;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2193;
wire n_2052;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_2091;
wire n_1517;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_2651;
wire n_3947;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_2099;
wire n_2408;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1071;
wire n_496;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_521;
wire n_3744;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_680;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_553;
wire n_901;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3550;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3542;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_446;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_464;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_477;
wire n_3191;
wire n_571;
wire n_1585;
wire n_461;
wire n_2684;
wire n_2712;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3837;
wire n_1971;
wire n_1599;
wire n_3936;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2700;
wire n_2644;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_907;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_3915;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_3714;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_3651;
wire n_3310;
wire n_593;
wire n_3487;
wire n_2258;
wire n_4069;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_3781;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_884;
wire n_3328;
wire n_944;
wire n_1754;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_647;
wire n_3433;
wire n_4024;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_857;
wire n_832;
wire n_2305;
wire n_3430;
wire n_3392;
wire n_3975;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_561;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_686;
wire n_3989;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_558;
wire n_3655;
wire n_2808;
wire n_702;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_822;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_728;
wire n_2930;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_809;
wire n_3923;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_3895;
wire n_3643;
wire n_2222;
wire n_1892;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_747;
wire n_2064;
wire n_784;
wire n_3978;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_776;
wire n_1798;
wire n_2022;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_3416;
wire n_452;
wire n_525;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_498;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3113;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_524;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_456;
wire n_959;
wire n_2459;
wire n_3031;
wire n_535;
wire n_3396;
wire n_3701;
wire n_940;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2320;
wire n_2473;
wire n_2038;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_442;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3820;
wire n_636;
wire n_3741;
wire n_660;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_459;
wire n_2312;
wire n_3990;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_473;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_3149;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_2897;
wire n_2077;
wire n_1416;
wire n_3614;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_3466;
wire n_3458;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_761;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_2110;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_582;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_2367;
wire n_512;
wire n_1870;
wire n_1591;
wire n_2033;
wire n_4071;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3929;
wire n_3077;
wire n_3838;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_3675;
wire n_2424;
wire n_2255;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_441;
wire n_860;
wire n_3229;
wire n_450;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_513;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3618;
wire n_3592;
wire n_4031;
wire n_495;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_824;
wire n_3808;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3824;
wire n_2662;
wire n_2740;
wire n_3890;
wire n_3751;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_1630;
wire n_716;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_531;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_950;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_444;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_912;
wire n_968;
wire n_3548;
wire n_451;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_3953;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_1357;
wire n_483;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_455;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3299;
wire n_3041;
wire n_3274;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2685;
wire n_2037;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_3913;
wire n_3737;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_3866;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_943;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_543;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_4029;
wire n_3400;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_918;
wire n_3854;
wire n_3529;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_540;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_1511;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2393;
wire n_833;
wire n_2318;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2793;
wire n_2707;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_3998;
wire n_2285;
wire n_1446;
wire n_3147;
wire n_2758;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_3869;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_4010;
wire n_1204;
wire n_3708;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_1722;
wire n_3957;
wire n_661;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_510;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_3697;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_836;
wire n_990;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_458;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_601;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2722;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1335;
wire n_1777;
wire n_1514;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_3967;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_1584;
wire n_487;
wire n_1726;
wire n_665;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_3972;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_3639;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_3308;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_791;
wire n_732;
wire n_1533;
wire n_1979;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_808;
wire n_2484;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_500;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_766;
wire n_3928;
wire n_541;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_536;
wire n_3438;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_827;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_3968;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_703;
wire n_698;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3239;
wire n_3139;
wire n_2773;
wire n_3172;
wire n_3292;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1530;
wire n_1497;
wire n_4075;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_867;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_760;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_622;
wire n_1962;
wire n_3996;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_3391;
wire n_682;
wire n_1567;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_4015;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_479;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_3903;
wire n_3551;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3859;
wire n_3865;
wire n_3722;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_3251;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_462;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_722;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_471;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_474;
wire n_2940;
wire n_542;
wire n_3435;
wire n_3521;
wire n_463;
wire n_3575;
wire n_1546;
wire n_595;
wire n_502;
wire n_3562;
wire n_3948;
wire n_466;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2505;
wire n_2438;
wire n_2427;
wire n_1673;
wire n_465;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_3250;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3921;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_2196;
wire n_3591;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_494;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_3930;
wire n_730;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_3772;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_453;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_491;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_3225;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_206),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_357),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_316),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_247),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_89),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_29),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_84),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_49),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_270),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_327),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_191),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_173),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_300),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_272),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_235),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_258),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_265),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_10),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_237),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_3),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_208),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_137),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_118),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_410),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_135),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_190),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_433),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_121),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_124),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_135),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_5),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_250),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_368),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_27),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_175),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_260),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_95),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_170),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_128),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_235),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_105),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_14),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_196),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_405),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_156),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_427),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_118),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_308),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_65),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_249),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_41),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_146),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_146),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_263),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_191),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_8),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_208),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_366),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_311),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_258),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_22),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_215),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_206),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_277),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_26),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_271),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_40),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_401),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_388),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_223),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_83),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_257),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_425),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_156),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_173),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_119),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_306),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_89),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_299),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_280),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_90),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_132),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_421),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_8),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_0),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_403),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_333),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_259),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_230),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_162),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_275),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_27),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_165),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_76),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_239),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_203),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_372),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_341),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_139),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_194),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_435),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_204),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_392),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_276),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_330),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_262),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_419),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_128),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_226),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_153),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_117),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_342),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_246),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_15),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_395),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_200),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_430),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_282),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_219),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_163),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_434),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_168),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_387),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_356),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_60),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_59),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_166),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_102),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_210),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_22),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_254),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_292),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_432),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_398),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_220),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_232),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_9),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_48),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_38),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_123),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_270),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_255),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_29),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_411),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_169),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_307),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_391),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_385),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_72),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_198),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_369),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_189),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_423),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_39),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_312),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_218),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_352),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_416),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_436),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_344),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_67),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_310),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_370),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_57),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_228),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_297),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_5),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_73),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_271),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_187),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_402),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_371),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_377),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_125),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_79),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_414),
.Y(n_622)
);

BUFx8_ASAP7_75t_SL g623 ( 
.A(n_205),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_334),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_111),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_131),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_288),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_227),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_186),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_132),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_52),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_158),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_172),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_275),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_151),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_386),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_413),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_328),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_230),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_229),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_127),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_273),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_34),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_431),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_382),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_59),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_153),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_215),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_346),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_282),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_50),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_284),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_319),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_359),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_418),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_164),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_243),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_379),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_185),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_104),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_92),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_209),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_396),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_152),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_276),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_376),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_83),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_412),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_104),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_26),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_81),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_127),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_201),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_309),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_172),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_353),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_82),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_20),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_246),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_322),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_227),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_422),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_165),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_323),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_94),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_221),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_320),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_409),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_90),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_241),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_62),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_47),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_145),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_304),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_358),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_294),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_6),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_95),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_60),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_362),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_47),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_122),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_55),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_45),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_79),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_374),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_228),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_169),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_88),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_185),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_101),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_4),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_46),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_278),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_326),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_203),
.Y(n_716)
);

BUFx5_ASAP7_75t_L g717 ( 
.A(n_417),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_115),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_18),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_209),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_98),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_219),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_400),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_134),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_339),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_35),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_214),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_197),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_124),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_30),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_244),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_39),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_167),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_102),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_75),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_192),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_35),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_17),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_298),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_340),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_284),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_315),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_194),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_92),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_216),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_55),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_365),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_236),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_138),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_259),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_70),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_54),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_36),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_34),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_0),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_161),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_278),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_32),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_141),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_446),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_623),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_463),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_629),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_621),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_643),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_497),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_463),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_541),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_552),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_497),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_552),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_510),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_440),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_510),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_621),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_443),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_525),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_486),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_447),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_541),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_525),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_453),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_527),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_621),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_621),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_454),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_455),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_464),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_456),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_527),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_463),
.Y(n_792)
);

BUFx5_ASAP7_75t_L g793 ( 
.A(n_530),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_458),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_530),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_531),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_531),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_542),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_467),
.Y(n_799)
);

BUFx5_ASAP7_75t_L g800 ( 
.A(n_542),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_460),
.Y(n_801)
);

XNOR2xp5_ASAP7_75t_L g802 ( 
.A(n_738),
.B(n_1),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_551),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_462),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_487),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_551),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_556),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_556),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_486),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_465),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_569),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_457),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_468),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_469),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_569),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_470),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_570),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_472),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_511),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_518),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_561),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_463),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_474),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_475),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_478),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_481),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_570),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_578),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_480),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_578),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_463),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_490),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_492),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_446),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_493),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_580),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_494),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_446),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_580),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_593),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_593),
.Y(n_841)
);

CKINVDCx16_ASAP7_75t_R g842 ( 
.A(n_528),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_594),
.Y(n_843)
);

XNOR2xp5_ASAP7_75t_L g844 ( 
.A(n_479),
.B(n_1),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_495),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_541),
.Y(n_846)
);

INVxp33_ASAP7_75t_SL g847 ( 
.A(n_625),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_594),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_446),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_446),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_446),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_483),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_496),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_448),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_448),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_448),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_448),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_448),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_448),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_499),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_537),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_502),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_537),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_537),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_481),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_601),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_463),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_504),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_537),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_503),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_537),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_505),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_537),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_617),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_652),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_652),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_619),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_652),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_568),
.Y(n_879)
);

CKINVDCx16_ASAP7_75t_R g880 ( 
.A(n_644),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_506),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_603),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_609),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_603),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_604),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_604),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_652),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_618),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_618),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_622),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_507),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_508),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_633),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_663),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_622),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_627),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_648),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_627),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_723),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_636),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_509),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_512),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_636),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_645),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_514),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_609),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_441),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_645),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_653),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_720),
.B(n_2),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_517),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_522),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_653),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_654),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_442),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_654),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_524),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_655),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_526),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_655),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_658),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_609),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_532),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_658),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_534),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_535),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_666),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_642),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_666),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_674),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_673),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_538),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_539),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_540),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_674),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_682),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_449),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_742),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_543),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_544),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_546),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_550),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_682),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_452),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_684),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_684),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_553),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_473),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_554),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_555),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_501),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_695),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_695),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_652),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_739),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_739),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_740),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_557),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_740),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_747),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_562),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_564),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_652),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_747),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_742),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_677),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_481),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_742),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_584),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_677),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_584),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_690),
.Y(n_972)
);

BUFx10_ASAP7_75t_L g973 ( 
.A(n_677),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_584),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_567),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_677),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_631),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_677),
.Y(n_978)
);

CKINVDCx16_ASAP7_75t_R g979 ( 
.A(n_501),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_631),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_573),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_498),
.B(n_3),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_631),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_735),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_735),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_575),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_488),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_735),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_500),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_568),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_515),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_491),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_501),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_491),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_577),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_677),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_581),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_628),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_628),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_501),
.Y(n_1000)
);

INVxp33_ASAP7_75t_SL g1001 ( 
.A(n_583),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_491),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_568),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_585),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_588),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_589),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_547),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_606),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_591),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_519),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_595),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_596),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_628),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_606),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_563),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_630),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_630),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_606),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_598),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_521),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_700),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_630),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_700),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_602),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_700),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_444),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_529),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_607),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_444),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_545),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_450),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_612),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_613),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_450),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_547),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_614),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_451),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_451),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_620),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_549),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_626),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_634),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_461),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_461),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_635),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_559),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_639),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_702),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_566),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_568),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_641),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_471),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_471),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_624),
.B(n_4),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_579),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_476),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_498),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_476),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_477),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_477),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_650),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_489),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_590),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_651),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_650),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_650),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_568),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_681),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_656),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_657),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_489),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_681),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_659),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_610),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_610),
.B(n_6),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_513),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_568),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_660),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_662),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_664),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_513),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_516),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_516),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_523),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_667),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_523),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_533),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_592),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_533),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_624),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_669),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_670),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_672),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_536),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_536),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_548),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_548),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_681),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_711),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_678),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_711),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_711),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_736),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_597),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_736),
.Y(n_1105)
);

BUFx5_ASAP7_75t_L g1106 ( 
.A(n_558),
.Y(n_1106)
);

CKINVDCx16_ASAP7_75t_R g1107 ( 
.A(n_640),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_679),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_599),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_760),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_764),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_907),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_915),
.Y(n_1113)
);

INVxp33_ASAP7_75t_SL g1114 ( 
.A(n_802),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_789),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_764),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_937),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_944),
.Y(n_1118)
);

BUFx2_ASAP7_75t_SL g1119 ( 
.A(n_948),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_987),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_775),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_775),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_785),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_989),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_799),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_785),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_786),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_819),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_786),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_769),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_760),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_849),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_769),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_768),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_991),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_768),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_849),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_850),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1010),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1020),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_850),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_866),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1027),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_874),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_851),
.Y(n_1145)
);

INVxp67_ASAP7_75t_SL g1146 ( 
.A(n_780),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_851),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_762),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_877),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_854),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1030),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_854),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_834),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_855),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1040),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_855),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_856),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_856),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_857),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1046),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_857),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1049),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_821),
.B(n_687),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_858),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_899),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_938),
.B(n_1063),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1055),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_858),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1001),
.B(n_484),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_1088),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1104),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_859),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1109),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_880),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_859),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_780),
.B(n_736),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_894),
.Y(n_1177)
);

INVxp33_ASAP7_75t_L g1178 ( 
.A(n_763),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_861),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_846),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_778),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_809),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1063),
.B(n_605),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_812),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_861),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_761),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_761),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_863),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_846),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_863),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_773),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1015),
.B(n_649),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_864),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_773),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_771),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_864),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_776),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_834),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_869),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_869),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_852),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_868),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_776),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_893),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_897),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_931),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_779),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_972),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_871),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_871),
.Y(n_1210)
);

INVxp67_ASAP7_75t_SL g1211 ( 
.A(n_883),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_779),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_1048),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_771),
.Y(n_1214)
);

INVxp33_ASAP7_75t_SL g1215 ( 
.A(n_802),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_782),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_873),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_873),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_875),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_782),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_787),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_875),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_787),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_876),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_876),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_878),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_878),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_951),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_788),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_993),
.B(n_608),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_967),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_969),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_971),
.Y(n_1233)
);

NOR2xp67_ASAP7_75t_L g1234 ( 
.A(n_788),
.B(n_637),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_974),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_790),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_977),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_979),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_980),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_790),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_794),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_887),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_983),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_794),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_984),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_842),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_985),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_801),
.B(n_638),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_801),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_804),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_804),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_810),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_766),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_810),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_887),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_813),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_813),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_814),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_814),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_770),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_816),
.Y(n_1261)
);

INVxp33_ASAP7_75t_L g1262 ( 
.A(n_928),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_816),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_818),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_772),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_774),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_777),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_781),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_784),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_791),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_818),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_823),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_795),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_993),
.B(n_668),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_796),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_797),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_798),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_823),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_954),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1000),
.B(n_676),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_824),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_883),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_824),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_803),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_825),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_829),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_806),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_829),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_832),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_807),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_808),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_811),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_815),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_832),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_817),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_833),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_827),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_828),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_830),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_906),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_833),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_906),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_954),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_835),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_835),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_837),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_836),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_839),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_837),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_845),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_845),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_840),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_841),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_843),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_847),
.B(n_680),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_848),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_882),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_884),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_885),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_886),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_853),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_888),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1000),
.B(n_688),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_853),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_889),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_860),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_890),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_895),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_896),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_898),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_900),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_860),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_903),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_862),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_904),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_966),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_862),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_966),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_870),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_870),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_908),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_872),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_872),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_881),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_909),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_881),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_913),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_891),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_914),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_SL g1350 ( 
.A(n_1007),
.Y(n_1350)
);

BUFx2_ASAP7_75t_SL g1351 ( 
.A(n_1032),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_916),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_918),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_891),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_920),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1007),
.B(n_694),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_921),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_892),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_924),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_892),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_901),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_901),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_902),
.Y(n_1363)
);

NAND2xp33_ASAP7_75t_R g1364 ( 
.A(n_902),
.B(n_683),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_905),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_R g1366 ( 
.A(n_905),
.B(n_911),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_927),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_929),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1035),
.B(n_696),
.Y(n_1369)
);

CKINVDCx14_ASAP7_75t_R g1370 ( 
.A(n_783),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1032),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_911),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_912),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_930),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_935),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_936),
.Y(n_1376)
);

CKINVDCx16_ASAP7_75t_R g1377 ( 
.A(n_1057),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_912),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_943),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_917),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_917),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_919),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_945),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_919),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_946),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_952),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_923),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_953),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_955),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_956),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_970),
.Y(n_1391)
);

INVxp33_ASAP7_75t_SL g1392 ( 
.A(n_923),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_970),
.Y(n_1393)
);

INVxp33_ASAP7_75t_L g1394 ( 
.A(n_805),
.Y(n_1394)
);

CKINVDCx14_ASAP7_75t_R g1395 ( 
.A(n_783),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_925),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_976),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1035),
.B(n_706),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_976),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_925),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_978),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_978),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1131),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1169),
.A2(n_932),
.B1(n_933),
.B2(n_926),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1148),
.Y(n_1405)
);

XNOR2xp5_ASAP7_75t_L g1406 ( 
.A(n_1114),
.B(n_844),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1153),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1148),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1192),
.A2(n_1074),
.B1(n_1107),
.B2(n_1054),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1132),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1134),
.B(n_922),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1110),
.A2(n_1179),
.B(n_1175),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1153),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1231),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1146),
.B(n_1090),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1148),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1137),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1114),
.A2(n_844),
.B1(n_765),
.B2(n_466),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1198),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1198),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1138),
.Y(n_1421)
);

NOR2x1_ASAP7_75t_L g1422 ( 
.A(n_1351),
.B(n_965),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1134),
.B(n_965),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1141),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1145),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1176),
.B(n_1232),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1242),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1147),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1184),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1136),
.B(n_968),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1242),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1201),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1150),
.Y(n_1433)
);

OAI22x1_ASAP7_75t_SL g1434 ( 
.A1(n_1215),
.A2(n_686),
.B1(n_697),
.B2(n_685),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1152),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1279),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1189),
.B(n_1090),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1279),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1176),
.B(n_968),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1364),
.A2(n_932),
.B1(n_933),
.B2(n_926),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1136),
.B(n_998),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1180),
.B(n_998),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1211),
.B(n_1090),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1110),
.A2(n_1179),
.B(n_1175),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1176),
.B(n_826),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1185),
.A2(n_994),
.B(n_992),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1202),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1336),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1336),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1338),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1154),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1156),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1282),
.B(n_1090),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1180),
.B(n_1300),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1394),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1233),
.B(n_826),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1338),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1315),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1235),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1255),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1237),
.Y(n_1461)
);

INVx5_ASAP7_75t_L g1462 ( 
.A(n_1294),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1302),
.B(n_1090),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1157),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1158),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1255),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1166),
.B(n_934),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1159),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1161),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1164),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1215),
.A2(n_482),
.B1(n_485),
.B2(n_445),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1168),
.Y(n_1472)
);

INVx4_ASAP7_75t_L g1473 ( 
.A(n_1172),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1196),
.Y(n_1474)
);

AND2x2_ASAP7_75t_R g1475 ( 
.A(n_1370),
.B(n_558),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1303),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1303),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1199),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1185),
.A2(n_1008),
.B(n_1002),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1200),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1239),
.B(n_1243),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1209),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1188),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1163),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1351),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1323),
.B(n_793),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1245),
.B(n_865),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1188),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1234),
.A2(n_939),
.B1(n_941),
.B2(n_940),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1391),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1204),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1210),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1393),
.Y(n_1493)
);

BUFx8_ASAP7_75t_L g1494 ( 
.A(n_1350),
.Y(n_1494)
);

AOI22x1_ASAP7_75t_SL g1495 ( 
.A1(n_1271),
.A2(n_701),
.B1(n_703),
.B2(n_698),
.Y(n_1495)
);

CKINVDCx6p67_ASAP7_75t_R g1496 ( 
.A(n_1377),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1395),
.A2(n_910),
.B1(n_940),
.B2(n_939),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1190),
.A2(n_1018),
.B(n_1014),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1247),
.B(n_999),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1205),
.A2(n_520),
.B1(n_719),
.B2(n_615),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1183),
.B(n_941),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1217),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1218),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1219),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1369),
.B(n_793),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1190),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1248),
.A2(n_947),
.B1(n_949),
.B2(n_942),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1222),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1230),
.A2(n_996),
.B(n_1021),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1371),
.B(n_1253),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1224),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1274),
.A2(n_942),
.B1(n_949),
.B2(n_947),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1225),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1226),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1193),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1260),
.B(n_999),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1227),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1398),
.B(n_793),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1280),
.B(n_793),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1193),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1356),
.A2(n_950),
.B1(n_961),
.B2(n_958),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_R g1522 ( 
.A(n_1112),
.B(n_950),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1371),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_1025),
.B(n_1023),
.Y(n_1524)
);

INVx5_ASAP7_75t_L g1525 ( 
.A(n_1294),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1397),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1392),
.A2(n_958),
.B1(n_962),
.B2(n_961),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1265),
.B(n_1013),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1266),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1397),
.A2(n_996),
.B(n_959),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1399),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1267),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1268),
.B(n_793),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1399),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1269),
.B(n_865),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1401),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1270),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1401),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1402),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1130),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1273),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1402),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1206),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1275),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1276),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1111),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1277),
.B(n_988),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1208),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1116),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1284),
.B(n_793),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1287),
.Y(n_1551)
);

BUFx8_ASAP7_75t_L g1552 ( 
.A(n_1350),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1121),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1122),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1123),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1126),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1290),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1112),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1392),
.A2(n_975),
.B1(n_981),
.B2(n_962),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1291),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1213),
.A2(n_741),
.B1(n_707),
.B2(n_708),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1127),
.A2(n_960),
.B(n_957),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1129),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1292),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1293),
.A2(n_820),
.B1(n_981),
.B2(n_975),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1133),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1214),
.A2(n_710),
.B1(n_713),
.B2(n_704),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1295),
.B(n_988),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1297),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1298),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1299),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1113),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1307),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1308),
.B(n_1013),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1312),
.B(n_982),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1313),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1314),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1316),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1317),
.B(n_793),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1318),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1319),
.Y(n_1581)
);

INVxp33_ASAP7_75t_SL g1582 ( 
.A(n_1366),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1320),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1322),
.B(n_1325),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1327),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1328),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1329),
.B(n_800),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1330),
.B(n_1331),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1333),
.B(n_1016),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1335),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1341),
.B(n_1098),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1345),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1347),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1349),
.B(n_1352),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1113),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1353),
.B(n_800),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1355),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1130),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1357),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_L g1600 ( 
.A(n_1359),
.B(n_1367),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1368),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1374),
.B(n_1016),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1375),
.B(n_800),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1376),
.B(n_800),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1262),
.B(n_986),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1379),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1383),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1117),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1385),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1386),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1388),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1117),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1389),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1390),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1195),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1350),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_L g1617 ( 
.A(n_1254),
.B(n_717),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1257),
.B(n_800),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1263),
.B(n_800),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1178),
.B(n_995),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1289),
.A2(n_964),
.B(n_1017),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1340),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1400),
.A2(n_997),
.B1(n_1004),
.B2(n_995),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1346),
.Y(n_1624)
);

INVx5_ASAP7_75t_L g1625 ( 
.A(n_1246),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1191),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1354),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1360),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1194),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1197),
.B(n_1017),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1197),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1203),
.B(n_1098),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1203),
.B(n_800),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1207),
.A2(n_1061),
.B(n_1022),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1207),
.B(n_800),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1212),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1212),
.A2(n_1061),
.B(n_1022),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1216),
.A2(n_1004),
.B1(n_1005),
.B2(n_997),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1216),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1220),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1220),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1221),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1221),
.B(n_1065),
.Y(n_1643)
);

INVx5_ASAP7_75t_L g1644 ( 
.A(n_1223),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1223),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1229),
.A2(n_1066),
.B(n_1065),
.Y(n_1646)
);

AND2x6_ASAP7_75t_L g1647 ( 
.A(n_1182),
.B(n_746),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1229),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1236),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1236),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1240),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1181),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1240),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1241),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1241),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1244),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1244),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1249),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1250),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1250),
.A2(n_1068),
.B(n_1066),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1251),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1251),
.B(n_1005),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1252),
.B(n_1068),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1252),
.A2(n_1072),
.B(n_1099),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1256),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1256),
.B(n_1006),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1258),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1258),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1259),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1259),
.A2(n_1009),
.B1(n_1011),
.B2(n_1006),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1261),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1261),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1264),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1264),
.B(n_1072),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1272),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1272),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1278),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1278),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1281),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1283),
.A2(n_1012),
.B1(n_1019),
.B2(n_1011),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1283),
.Y(n_1681)
);

OAI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1458),
.A2(n_1019),
.B1(n_1024),
.B2(n_1012),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1467),
.A2(n_1288),
.B1(n_1311),
.B2(n_1305),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1530),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1455),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1418),
.A2(n_1125),
.B1(n_1128),
.B2(n_1115),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1406),
.A2(n_1144),
.B1(n_1149),
.B2(n_1142),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1407),
.Y(n_1688)
);

OAI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1618),
.A2(n_1619),
.B1(n_1409),
.B2(n_1633),
.Y(n_1689)
);

OAI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1635),
.A2(n_1305),
.B1(n_1311),
.B2(n_1288),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1632),
.B(n_1085),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1501),
.A2(n_1324),
.B1(n_1337),
.B2(n_1332),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1617),
.A2(n_1647),
.B1(n_1510),
.B2(n_1454),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1617),
.A2(n_1324),
.B1(n_1337),
.B2(n_1332),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1530),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1632),
.B(n_1108),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_R g1697 ( 
.A1(n_1605),
.A2(n_560),
.B1(n_571),
.B2(n_565),
.Y(n_1697)
);

OAI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1440),
.A2(n_1342),
.B1(n_1343),
.B2(n_1339),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1530),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1647),
.A2(n_1510),
.B1(n_1454),
.B2(n_1426),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1484),
.A2(n_1033),
.B1(n_1036),
.B2(n_1028),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1404),
.A2(n_1358),
.B1(n_1362),
.B2(n_1348),
.Y(n_1702)
);

AO22x2_ASAP7_75t_L g1703 ( 
.A1(n_1495),
.A2(n_756),
.B1(n_671),
.B2(n_560),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1429),
.B(n_1119),
.Y(n_1704)
);

AO22x2_ASAP7_75t_L g1705 ( 
.A1(n_1495),
.A2(n_565),
.B1(n_572),
.B2(n_571),
.Y(n_1705)
);

AO22x2_ASAP7_75t_L g1706 ( 
.A1(n_1623),
.A2(n_572),
.B1(n_576),
.B2(n_574),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1647),
.A2(n_1621),
.B1(n_1439),
.B2(n_1426),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1647),
.A2(n_1075),
.B1(n_1372),
.B2(n_1365),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1647),
.A2(n_1373),
.B1(n_1378),
.B2(n_1372),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1621),
.A2(n_1378),
.B1(n_1380),
.B2(n_1373),
.Y(n_1710)
);

AO22x2_ASAP7_75t_L g1711 ( 
.A1(n_1680),
.A2(n_1645),
.B1(n_1648),
.B2(n_1629),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1630),
.B(n_1108),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1620),
.B(n_1380),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1621),
.A2(n_1387),
.B1(n_1381),
.B2(n_1039),
.Y(n_1714)
);

AO22x2_ASAP7_75t_L g1715 ( 
.A1(n_1629),
.A2(n_574),
.B1(n_582),
.B2(n_576),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1532),
.A2(n_1387),
.B1(n_1381),
.B2(n_1039),
.Y(n_1716)
);

OAI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1532),
.A2(n_1041),
.B1(n_1042),
.B2(n_1036),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1407),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1578),
.B(n_1041),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1630),
.B(n_1119),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1413),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1429),
.B(n_1062),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1578),
.B(n_1042),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1441),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1406),
.A2(n_1165),
.B1(n_1173),
.B2(n_1170),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1630),
.B(n_1045),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1413),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1530),
.Y(n_1728)
);

AO22x2_ASAP7_75t_L g1729 ( 
.A1(n_1645),
.A2(n_582),
.B1(n_587),
.B2(n_586),
.Y(n_1729)
);

AND2x6_ASAP7_75t_L g1730 ( 
.A(n_1616),
.B(n_746),
.Y(n_1730)
);

AOI22x1_ASAP7_75t_SL g1731 ( 
.A1(n_1558),
.A2(n_1120),
.B1(n_1124),
.B2(n_1118),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1598),
.B(n_1047),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1441),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_R g1734 ( 
.A1(n_1627),
.A2(n_586),
.B1(n_600),
.B2(n_587),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1412),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1412),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1454),
.A2(n_1182),
.B1(n_1064),
.B2(n_1069),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1662),
.B(n_1051),
.Y(n_1738)
);

AND2x2_ASAP7_75t_SL g1739 ( 
.A(n_1626),
.B(n_746),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1666),
.B(n_1051),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1643),
.A2(n_1069),
.B1(n_1070),
.B2(n_1064),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1537),
.A2(n_1073),
.B1(n_1078),
.B2(n_1070),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1643),
.B(n_1073),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1643),
.B(n_1078),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1578),
.B(n_1079),
.Y(n_1745)
);

AO22x2_ASAP7_75t_L g1746 ( 
.A1(n_1648),
.A2(n_600),
.B1(n_616),
.B2(n_611),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1412),
.Y(n_1747)
);

AO22x2_ASAP7_75t_L g1748 ( 
.A1(n_1649),
.A2(n_611),
.B1(n_632),
.B2(n_616),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1419),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1663),
.B(n_1079),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1663),
.B(n_1080),
.Y(n_1751)
);

OAI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1537),
.A2(n_1091),
.B1(n_1092),
.B2(n_1080),
.Y(n_1752)
);

AO22x2_ASAP7_75t_L g1753 ( 
.A1(n_1649),
.A2(n_632),
.B1(n_647),
.B2(n_646),
.Y(n_1753)
);

BUFx10_ASAP7_75t_L g1754 ( 
.A(n_1663),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1541),
.A2(n_1100),
.B1(n_1093),
.B2(n_752),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1674),
.B(n_1445),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1544),
.A2(n_752),
.B1(n_749),
.B2(n_1174),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1621),
.A2(n_1396),
.B1(n_1286),
.B2(n_1296),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1419),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1420),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1674),
.A2(n_1301),
.B1(n_1304),
.B2(n_1285),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1674),
.B(n_1445),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1432),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1439),
.A2(n_1384),
.B1(n_1309),
.B2(n_1310),
.Y(n_1764)
);

OAI22xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1544),
.A2(n_646),
.B1(n_661),
.B2(n_647),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1412),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1590),
.A2(n_1321),
.B1(n_1326),
.B2(n_1306),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1597),
.B(n_1106),
.Y(n_1768)
);

AO22x2_ASAP7_75t_L g1769 ( 
.A1(n_1650),
.A2(n_661),
.B1(n_675),
.B2(n_665),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1590),
.A2(n_1344),
.B1(n_1361),
.B2(n_1334),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1535),
.B(n_1174),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1545),
.A2(n_665),
.B1(n_689),
.B2(n_675),
.Y(n_1772)
);

AO22x2_ASAP7_75t_L g1773 ( 
.A1(n_1650),
.A2(n_689),
.B1(n_692),
.B2(n_691),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1471),
.A2(n_1500),
.B1(n_1561),
.B2(n_1382),
.Y(n_1774)
);

OR2x6_ASAP7_75t_L g1775 ( 
.A(n_1432),
.B(n_691),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1535),
.B(n_1177),
.Y(n_1776)
);

OR2x6_ASAP7_75t_L g1777 ( 
.A(n_1447),
.B(n_692),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1441),
.Y(n_1778)
);

AO22x2_ASAP7_75t_L g1779 ( 
.A1(n_1661),
.A2(n_693),
.B1(n_705),
.B2(n_699),
.Y(n_1779)
);

AO22x2_ASAP7_75t_L g1780 ( 
.A1(n_1661),
.A2(n_693),
.B1(n_705),
.B2(n_699),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1590),
.A2(n_1363),
.B1(n_715),
.B2(n_725),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1593),
.A2(n_1187),
.B1(n_1186),
.B2(n_1228),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1551),
.A2(n_709),
.B1(n_714),
.B2(n_712),
.Y(n_1783)
);

OAI22xp33_ASAP7_75t_SL g1784 ( 
.A1(n_1551),
.A2(n_709),
.B1(n_714),
.B2(n_712),
.Y(n_1784)
);

OAI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1560),
.A2(n_1577),
.B1(n_1583),
.B2(n_1571),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1411),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1444),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1593),
.A2(n_1187),
.B1(n_1186),
.B2(n_1238),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1447),
.B(n_1118),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1597),
.B(n_1106),
.Y(n_1790)
);

AO22x2_ASAP7_75t_L g1791 ( 
.A1(n_1669),
.A2(n_724),
.B1(n_726),
.B2(n_718),
.Y(n_1791)
);

AO22x2_ASAP7_75t_L g1792 ( 
.A1(n_1669),
.A2(n_1672),
.B1(n_1681),
.B2(n_1677),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1560),
.A2(n_716),
.B1(n_459),
.B2(n_718),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1547),
.B(n_1124),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1420),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1547),
.B(n_1135),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1427),
.Y(n_1797)
);

NAND3x1_ASAP7_75t_L g1798 ( 
.A(n_1638),
.B(n_726),
.C(n_724),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1571),
.A2(n_459),
.B1(n_728),
.B2(n_727),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1436),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1577),
.A2(n_728),
.B1(n_729),
.B2(n_727),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1491),
.B(n_1543),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1436),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1599),
.A2(n_1140),
.B1(n_1143),
.B2(n_1139),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1450),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1567),
.A2(n_1155),
.B1(n_1160),
.B2(n_1151),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1444),
.Y(n_1807)
);

AO22x2_ASAP7_75t_L g1808 ( 
.A1(n_1672),
.A2(n_732),
.B1(n_733),
.B2(n_729),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1450),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1457),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1543),
.B(n_1151),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1411),
.B(n_1026),
.Y(n_1812)
);

AO22x2_ASAP7_75t_L g1813 ( 
.A1(n_1677),
.A2(n_733),
.B1(n_745),
.B2(n_732),
.Y(n_1813)
);

INVx8_ASAP7_75t_L g1814 ( 
.A(n_1625),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1485),
.B(n_1160),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1444),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1558),
.A2(n_1167),
.B1(n_1171),
.B2(n_1162),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1599),
.A2(n_1167),
.B1(n_1171),
.B2(n_1162),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1599),
.A2(n_1106),
.B1(n_717),
.B2(n_1031),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1457),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1444),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1536),
.Y(n_1822)
);

BUFx10_ASAP7_75t_L g1823 ( 
.A(n_1572),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1520),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1583),
.A2(n_748),
.B1(n_750),
.B2(n_745),
.Y(n_1825)
);

AO22x2_ASAP7_75t_L g1826 ( 
.A1(n_1681),
.A2(n_750),
.B1(n_751),
.B2(n_748),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1536),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1485),
.B(n_1032),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1568),
.B(n_1029),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1456),
.B(n_1034),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1670),
.B(n_721),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1548),
.B(n_751),
.Y(n_1832)
);

OAI22xp33_ASAP7_75t_SL g1833 ( 
.A1(n_1585),
.A2(n_754),
.B1(n_757),
.B2(n_753),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1582),
.B(n_722),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1536),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1512),
.A2(n_1106),
.B1(n_717),
.B2(n_1038),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1456),
.B(n_1037),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1597),
.B(n_1106),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1536),
.Y(n_1839)
);

AO22x2_ASAP7_75t_L g1840 ( 
.A1(n_1497),
.A2(n_754),
.B1(n_757),
.B2(n_753),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1548),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1536),
.Y(n_1842)
);

OA22x2_ASAP7_75t_L g1843 ( 
.A1(n_1559),
.A2(n_731),
.B1(n_734),
.B2(n_730),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1521),
.A2(n_1106),
.B1(n_717),
.B2(n_1044),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1487),
.B(n_1043),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1487),
.B(n_1052),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1442),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_SL g1848 ( 
.A1(n_1585),
.A2(n_743),
.B1(n_744),
.B2(n_737),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1588),
.A2(n_1594),
.B1(n_1423),
.B2(n_1430),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1460),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1566),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1595),
.A2(n_758),
.B1(n_759),
.B2(n_755),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1520),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1627),
.B(n_1053),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1523),
.A2(n_1101),
.B1(n_1102),
.B2(n_1099),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1527),
.B(n_1056),
.Y(n_1856)
);

INVxp67_ASAP7_75t_SL g1857 ( 
.A(n_1431),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_SL g1858 ( 
.A1(n_1595),
.A2(n_1059),
.B1(n_1060),
.B2(n_1058),
.Y(n_1858)
);

OA22x2_ASAP7_75t_L g1859 ( 
.A1(n_1628),
.A2(n_1076),
.B1(n_1081),
.B2(n_1071),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1483),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1588),
.A2(n_1106),
.B1(n_717),
.B2(n_1083),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1609),
.A2(n_1613),
.B1(n_1489),
.B2(n_1507),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1462),
.B(n_1082),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1608),
.A2(n_1086),
.B1(n_1087),
.B2(n_1084),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1592),
.A2(n_1106),
.B1(n_1089),
.B2(n_1095),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1592),
.A2(n_1094),
.B1(n_1097),
.B2(n_1096),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1610),
.A2(n_1102),
.B1(n_1103),
.B2(n_1101),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1610),
.A2(n_1103),
.B1(n_1105),
.B2(n_717),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1611),
.A2(n_1105),
.B1(n_717),
.B2(n_963),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1611),
.A2(n_767),
.B1(n_792),
.B2(n_762),
.Y(n_1870)
);

AND2x2_ASAP7_75t_SL g1871 ( 
.A(n_1626),
.B(n_762),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1540),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1614),
.A2(n_767),
.B1(n_792),
.B2(n_762),
.Y(n_1873)
);

OAI22xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1614),
.A2(n_11),
.B1(n_7),
.B2(n_10),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_SL g1875 ( 
.A1(n_1608),
.A2(n_12),
.B1(n_7),
.B2(n_11),
.Y(n_1875)
);

NAND3x1_ASAP7_75t_L g1876 ( 
.A(n_1653),
.B(n_12),
.C(n_13),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1462),
.A2(n_767),
.B1(n_792),
.B2(n_762),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1462),
.A2(n_1077),
.B1(n_792),
.B2(n_822),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1462),
.B(n_838),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1466),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1584),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1476),
.Y(n_1882)
);

OAI22xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1631),
.A2(n_1639),
.B1(n_1656),
.B2(n_1642),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1516),
.A2(n_717),
.B1(n_963),
.B2(n_838),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1476),
.Y(n_1885)
);

OAI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1462),
.A2(n_1077),
.B1(n_792),
.B2(n_822),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1525),
.B(n_838),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1477),
.Y(n_1888)
);

AO22x2_ASAP7_75t_L g1889 ( 
.A1(n_1631),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1483),
.Y(n_1890)
);

OR2x6_ASAP7_75t_L g1891 ( 
.A(n_1626),
.B(n_767),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1516),
.A2(n_1528),
.B1(n_1589),
.B2(n_1574),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1628),
.B(n_19),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1477),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1490),
.Y(n_1895)
);

OAI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1525),
.A2(n_822),
.B1(n_831),
.B2(n_767),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1525),
.B(n_963),
.Y(n_1897)
);

OAI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1525),
.A2(n_831),
.B1(n_867),
.B2(n_822),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1516),
.A2(n_717),
.B1(n_973),
.B2(n_831),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1483),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1588),
.A2(n_973),
.B1(n_831),
.B2(n_867),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1582),
.B(n_19),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1525),
.B(n_973),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1490),
.Y(n_1904)
);

OAI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1609),
.A2(n_1077),
.B1(n_831),
.B2(n_867),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1488),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1411),
.B(n_287),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1639),
.B(n_1077),
.Y(n_1908)
);

AND2x2_ASAP7_75t_SL g1909 ( 
.A(n_1626),
.B(n_822),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1488),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1423),
.B(n_289),
.Y(n_1911)
);

OAI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1613),
.A2(n_1580),
.B1(n_1586),
.B2(n_1573),
.Y(n_1912)
);

OAI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1573),
.A2(n_1077),
.B1(n_879),
.B2(n_990),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1488),
.Y(n_1914)
);

OAI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1580),
.A2(n_879),
.B1(n_990),
.B2(n_867),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1493),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1493),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1642),
.A2(n_1665),
.B1(n_1667),
.B2(n_1656),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1526),
.Y(n_1919)
);

OAI22xp33_ASAP7_75t_SL g1920 ( 
.A1(n_1665),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1506),
.Y(n_1921)
);

OA22x2_ASAP7_75t_L g1922 ( 
.A1(n_1622),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1667),
.B(n_1067),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1671),
.B(n_1067),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1423),
.B(n_290),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1430),
.B(n_291),
.Y(n_1926)
);

AO22x2_ASAP7_75t_L g1927 ( 
.A1(n_1671),
.A2(n_28),
.B1(n_24),
.B2(n_25),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1430),
.Y(n_1928)
);

AO22x2_ASAP7_75t_L g1929 ( 
.A1(n_1678),
.A2(n_31),
.B1(n_25),
.B2(n_28),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1678),
.B(n_1067),
.Y(n_1930)
);

OAI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1679),
.A2(n_1459),
.B1(n_1461),
.B2(n_1414),
.Y(n_1931)
);

AO22x2_ASAP7_75t_L g1932 ( 
.A1(n_1679),
.A2(n_36),
.B1(n_32),
.B2(n_33),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1526),
.Y(n_1933)
);

OA22x2_ASAP7_75t_L g1934 ( 
.A1(n_1624),
.A2(n_38),
.B1(n_33),
.B2(n_37),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1594),
.A2(n_879),
.B1(n_990),
.B2(n_867),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1442),
.B(n_293),
.Y(n_1936)
);

OAI22xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1653),
.A2(n_42),
.B1(n_37),
.B2(n_40),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1506),
.Y(n_1938)
);

AO22x2_ASAP7_75t_L g1939 ( 
.A1(n_1673),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1506),
.Y(n_1940)
);

OAI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1586),
.A2(n_990),
.B1(n_1003),
.B2(n_879),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1529),
.B(n_43),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1616),
.A2(n_990),
.B1(n_1003),
.B2(n_879),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1673),
.B(n_1067),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1442),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1531),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1594),
.A2(n_1050),
.B1(n_1067),
.B2(n_1003),
.Y(n_1947)
);

AO22x2_ASAP7_75t_L g1948 ( 
.A1(n_1655),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1515),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1515),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1529),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1515),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1531),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1953),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1824),
.B(n_1415),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1824),
.B(n_1437),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1831),
.B(n_1615),
.C(n_1626),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1860),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1853),
.B(n_1443),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1763),
.Y(n_1960)
);

OR2x6_ASAP7_75t_L g1961 ( 
.A(n_1814),
.B(n_1676),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1853),
.B(n_1453),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1860),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1814),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1756),
.A2(n_1664),
.B1(n_1473),
.B2(n_1569),
.Y(n_1965)
);

AND2x6_ASAP7_75t_L g1966 ( 
.A(n_1735),
.B(n_1636),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1890),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1953),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1890),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1739),
.B(n_1644),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1928),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1762),
.A2(n_1664),
.B1(n_1473),
.B2(n_1569),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1900),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1900),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1906),
.Y(n_1975)
);

INVx4_ASAP7_75t_SL g1976 ( 
.A(n_1735),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1906),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1910),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1693),
.B(n_1863),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1738),
.B(n_1463),
.Y(n_1980)
);

AND3x1_ASAP7_75t_L g1981 ( 
.A(n_1758),
.B(n_1600),
.C(n_1575),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1720),
.B(n_1644),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1740),
.B(n_1403),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1700),
.A2(n_1644),
.B1(n_1676),
.B2(n_1636),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1691),
.A2(n_1655),
.B(n_1581),
.Y(n_1985)
);

AND2x6_ASAP7_75t_L g1986 ( 
.A(n_1736),
.B(n_1636),
.Y(n_1986)
);

INVx6_ASAP7_75t_L g1987 ( 
.A(n_1928),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1914),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1921),
.Y(n_1989)
);

NAND2xp33_ASAP7_75t_SL g1990 ( 
.A(n_1862),
.B(n_1636),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1921),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1829),
.B(n_1664),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1938),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1908),
.B(n_1403),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1923),
.B(n_1410),
.Y(n_1995)
);

INVxp67_ASAP7_75t_SL g1996 ( 
.A(n_1928),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1924),
.B(n_1410),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1938),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1936),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1952),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1952),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1940),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1940),
.Y(n_2003)
);

BUFx10_ASAP7_75t_L g2004 ( 
.A(n_1713),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1754),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1949),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1949),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1830),
.B(n_1664),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1802),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1930),
.B(n_1417),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1754),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1724),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1950),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1950),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1785),
.B(n_1417),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1688),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_L g2017 ( 
.A(n_1736),
.B(n_1640),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1837),
.B(n_1640),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1709),
.B(n_1640),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1718),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1936),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1710),
.B(n_1640),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1854),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1684),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_1685),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1721),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1684),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1822),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1683),
.B(n_1641),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_L g2030 ( 
.A(n_1741),
.B(n_1651),
.C(n_1641),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1944),
.B(n_1724),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1695),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1695),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1710),
.B(n_1641),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1733),
.B(n_1421),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1871),
.B(n_1641),
.Y(n_2036)
);

INVx2_ASAP7_75t_SL g2037 ( 
.A(n_1733),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1778),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1851),
.B(n_1641),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1699),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1778),
.A2(n_1473),
.B1(n_1569),
.B2(n_1557),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1847),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1907),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1845),
.B(n_1651),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1847),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1699),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1719),
.B(n_1421),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1723),
.B(n_1745),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1850),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1728),
.Y(n_2050)
);

AO21x2_ASAP7_75t_L g2051 ( 
.A1(n_1707),
.A2(n_1634),
.B(n_1509),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1880),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1728),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1690),
.B(n_1651),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1882),
.Y(n_2055)
);

BUFx10_ASAP7_75t_L g2056 ( 
.A(n_1902),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1885),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1888),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1894),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1895),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1909),
.B(n_1424),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1708),
.B(n_1651),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1692),
.B(n_1651),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1904),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_1722),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1846),
.B(n_1654),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1732),
.B(n_1654),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1872),
.B(n_1654),
.Y(n_2068)
);

INVx1_ASAP7_75t_SL g2069 ( 
.A(n_1841),
.Y(n_2069)
);

AND2x6_ASAP7_75t_L g2070 ( 
.A(n_1747),
.B(n_1654),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1907),
.A2(n_1911),
.B1(n_1926),
.B2(n_1925),
.Y(n_2071)
);

NAND3xp33_ASAP7_75t_L g2072 ( 
.A(n_1714),
.B(n_1658),
.C(n_1657),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1945),
.B(n_1424),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_L g2074 ( 
.A(n_1747),
.B(n_1657),
.Y(n_2074)
);

INVx8_ASAP7_75t_L g2075 ( 
.A(n_1891),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1916),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1827),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1834),
.B(n_1657),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1917),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1716),
.B(n_1657),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1919),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1911),
.A2(n_1569),
.B1(n_1570),
.B2(n_1557),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1933),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_1925),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1696),
.B(n_1425),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1926),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1946),
.Y(n_2087)
);

NAND3xp33_ASAP7_75t_L g2088 ( 
.A(n_1714),
.B(n_1659),
.C(n_1658),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1823),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1789),
.B(n_1652),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1892),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1750),
.B(n_1658),
.Y(n_2092)
);

CKINVDCx20_ASAP7_75t_R g2093 ( 
.A(n_1687),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1794),
.B(n_1658),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1689),
.A2(n_1570),
.B1(n_1576),
.B2(n_1557),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1951),
.B(n_1425),
.Y(n_2096)
);

INVx6_ASAP7_75t_L g2097 ( 
.A(n_1891),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1892),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1727),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1749),
.Y(n_2100)
);

BUFx10_ASAP7_75t_L g2101 ( 
.A(n_1856),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1759),
.Y(n_2102)
);

BUFx10_ASAP7_75t_L g2103 ( 
.A(n_1942),
.Y(n_2103)
);

BUFx10_ASAP7_75t_L g2104 ( 
.A(n_1812),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1760),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1766),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1795),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_1722),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1797),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1800),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1803),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_1796),
.Y(n_2112)
);

AND2x6_ASAP7_75t_L g2113 ( 
.A(n_1766),
.B(n_1659),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1805),
.Y(n_2114)
);

OR2x2_ASAP7_75t_SL g2115 ( 
.A(n_1811),
.B(n_1659),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1694),
.B(n_1659),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1809),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1810),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1820),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1787),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_1812),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1883),
.B(n_1428),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1786),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1918),
.B(n_1668),
.Y(n_2124)
);

BUFx2_ASAP7_75t_L g2125 ( 
.A(n_1775),
.Y(n_2125)
);

NAND3xp33_ASAP7_75t_L g2126 ( 
.A(n_1737),
.B(n_1675),
.C(n_1668),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_1775),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_1835),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1859),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_L g2130 ( 
.A(n_1787),
.B(n_1668),
.Y(n_2130)
);

OAI22xp33_ASAP7_75t_SL g2131 ( 
.A1(n_1893),
.A2(n_1612),
.B1(n_1422),
.B2(n_1581),
.Y(n_2131)
);

CKINVDCx20_ASAP7_75t_R g2132 ( 
.A(n_1725),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_1771),
.B(n_1652),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1807),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_SL g2135 ( 
.A(n_1817),
.B(n_1612),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1807),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1816),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1816),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1821),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1821),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1839),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1842),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1712),
.B(n_1428),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1912),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1879),
.B(n_1433),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1887),
.B(n_1433),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1768),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1849),
.B(n_1668),
.Y(n_2148)
);

INVx1_ASAP7_75t_SL g2149 ( 
.A(n_1776),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1730),
.Y(n_2150)
);

INVx5_ASAP7_75t_L g2151 ( 
.A(n_1730),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_1702),
.B(n_1668),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_1764),
.B(n_1496),
.Y(n_2153)
);

NAND3xp33_ASAP7_75t_L g2154 ( 
.A(n_1726),
.B(n_1676),
.C(n_1675),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1707),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1865),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1790),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1743),
.B(n_1675),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1865),
.Y(n_2159)
);

AO22x2_ASAP7_75t_L g2160 ( 
.A1(n_1939),
.A2(n_1435),
.B1(n_1452),
.B2(n_1451),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1823),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1744),
.A2(n_1570),
.B1(n_1606),
.B2(n_1576),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1838),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1730),
.Y(n_2164)
);

BUFx10_ASAP7_75t_L g2165 ( 
.A(n_1704),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1868),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_1730),
.Y(n_2167)
);

OR2x6_ASAP7_75t_L g2168 ( 
.A(n_1704),
.B(n_1675),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_1897),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1751),
.B(n_1675),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1903),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1868),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1939),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1857),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1931),
.B(n_1676),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1836),
.Y(n_2176)
);

NAND3xp33_ASAP7_75t_L g2177 ( 
.A(n_1781),
.B(n_1676),
.C(n_1625),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_1758),
.B(n_1564),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1844),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1819),
.Y(n_2180)
);

AND2x2_ASAP7_75t_SL g2181 ( 
.A(n_1884),
.B(n_1637),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1777),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1855),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1792),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1717),
.B(n_1625),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_1861),
.B(n_1564),
.Y(n_2186)
);

AND3x2_ASAP7_75t_L g2187 ( 
.A(n_1948),
.B(n_1552),
.C(n_1494),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1742),
.B(n_1625),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_1876),
.Y(n_2189)
);

INVxp33_ASAP7_75t_L g2190 ( 
.A(n_1686),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1752),
.B(n_1625),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1698),
.B(n_1565),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1815),
.B(n_1576),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1889),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1889),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1927),
.Y(n_2196)
);

AND2x6_ASAP7_75t_L g2197 ( 
.A(n_1884),
.B(n_1519),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_1804),
.B(n_1481),
.C(n_1601),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1757),
.B(n_1451),
.Y(n_2199)
);

INVx4_ASAP7_75t_L g2200 ( 
.A(n_1927),
.Y(n_2200)
);

AOI22xp33_ASAP7_75t_L g2201 ( 
.A1(n_1843),
.A2(n_1606),
.B1(n_1465),
.B2(n_1468),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1755),
.B(n_1452),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1929),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1866),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1777),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1929),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1932),
.Y(n_2207)
);

AND2x6_ASAP7_75t_L g2208 ( 
.A(n_1869),
.B(n_1899),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_1711),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_1832),
.Y(n_2210)
);

INVxp33_ASAP7_75t_L g2211 ( 
.A(n_1761),
.Y(n_2211)
);

NOR2x1p5_ASAP7_75t_L g2212 ( 
.A(n_1697),
.B(n_1494),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1867),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1932),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1711),
.B(n_1465),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_1782),
.B(n_1606),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_1788),
.B(n_1522),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1899),
.Y(n_2218)
);

INVx5_ASAP7_75t_L g2219 ( 
.A(n_1937),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1840),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_1798),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_1818),
.B(n_1601),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1974),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_2106),
.Y(n_2224)
);

INVxp67_ASAP7_75t_L g2225 ( 
.A(n_2009),
.Y(n_2225)
);

BUFx4_ASAP7_75t_L g2226 ( 
.A(n_2220),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_1960),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2043),
.B(n_1481),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1974),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2089),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_1999),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1978),
.Y(n_2232)
);

AND2x6_ASAP7_75t_L g2233 ( 
.A(n_1999),
.B(n_1869),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1978),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1999),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1989),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1989),
.Y(n_2237)
);

OAI22xp33_ASAP7_75t_SL g2238 ( 
.A1(n_2189),
.A2(n_1828),
.B1(n_1767),
.B2(n_1770),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1993),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1993),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2149),
.B(n_1806),
.Y(n_2241)
);

AND2x4_ASAP7_75t_L g2242 ( 
.A(n_2043),
.B(n_1607),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1998),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1998),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2155),
.B(n_1637),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2048),
.B(n_1701),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_2009),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2002),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2002),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_2106),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2003),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2003),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_2089),
.Y(n_2253)
);

INVx4_ASAP7_75t_L g2254 ( 
.A(n_1999),
.Y(n_2254)
);

INVx4_ASAP7_75t_L g2255 ( 
.A(n_1999),
.Y(n_2255)
);

INVx4_ASAP7_75t_L g2256 ( 
.A(n_2021),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2006),
.Y(n_2257)
);

BUFx3_ASAP7_75t_L g2258 ( 
.A(n_1960),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_2086),
.B(n_1607),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2006),
.Y(n_2260)
);

INVx2_ASAP7_75t_SL g2261 ( 
.A(n_2025),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1968),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2106),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2071),
.B(n_1486),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2086),
.B(n_1591),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_2158),
.B(n_1591),
.Y(n_2266)
);

AOI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2155),
.A2(n_1990),
.B1(n_2173),
.B2(n_2098),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2021),
.B(n_1505),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2000),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_2106),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2001),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2007),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2021),
.B(n_1518),
.Y(n_2273)
);

AO22x2_ASAP7_75t_L g2274 ( 
.A1(n_2200),
.A2(n_1948),
.B1(n_1875),
.B2(n_1731),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_2106),
.Y(n_2275)
);

BUFx8_ASAP7_75t_L g2276 ( 
.A(n_2065),
.Y(n_2276)
);

NOR2x1p5_ASAP7_75t_L g2277 ( 
.A(n_2011),
.B(n_1494),
.Y(n_2277)
);

BUFx3_ASAP7_75t_L g2278 ( 
.A(n_2011),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_L g2279 ( 
.A(n_2112),
.B(n_1682),
.Y(n_2279)
);

NAND2xp33_ASAP7_75t_L g2280 ( 
.A(n_2021),
.B(n_1774),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1968),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1992),
.B(n_1637),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1954),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_L g2284 ( 
.A(n_2021),
.B(n_1901),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2007),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1954),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2013),
.Y(n_2287)
);

BUFx2_ASAP7_75t_L g2288 ( 
.A(n_2069),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2133),
.Y(n_2289)
);

AO22x2_ASAP7_75t_L g2290 ( 
.A1(n_2200),
.A2(n_2195),
.B1(n_2196),
.B2(n_2194),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_2140),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_1990),
.A2(n_2173),
.B1(n_2091),
.B2(n_2208),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2013),
.Y(n_2293)
);

INVx4_ASAP7_75t_L g2294 ( 
.A(n_1987),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2140),
.Y(n_2295)
);

NAND2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2084),
.B(n_1637),
.Y(n_2296)
);

AND2x6_ASAP7_75t_L g2297 ( 
.A(n_2140),
.B(n_1935),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2018),
.B(n_2044),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2014),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2044),
.B(n_1848),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2014),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2140),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2066),
.B(n_1715),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1958),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1963),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_2084),
.Y(n_2306)
);

OAI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2084),
.A2(n_1840),
.B1(n_1947),
.B2(n_1660),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_2170),
.B(n_1469),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_SL g2309 ( 
.A(n_2165),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2066),
.B(n_1469),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2099),
.Y(n_2311)
);

BUFx6f_ASAP7_75t_L g2312 ( 
.A(n_2084),
.Y(n_2312)
);

AND2x6_ASAP7_75t_L g2313 ( 
.A(n_2084),
.B(n_1472),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1992),
.B(n_1646),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1967),
.Y(n_2315)
);

OAI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2082),
.A2(n_1660),
.B1(n_1646),
.B2(n_1480),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1973),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1975),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_1983),
.B(n_1472),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1977),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2101),
.B(n_1852),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2099),
.Y(n_2322)
);

AOI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2094),
.A2(n_1480),
.B1(n_1492),
.B2(n_1482),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2008),
.B(n_1646),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2100),
.Y(n_2325)
);

NAND3x1_ASAP7_75t_L g2326 ( 
.A(n_2192),
.B(n_1434),
.C(n_1475),
.Y(n_2326)
);

INVx4_ASAP7_75t_L g2327 ( 
.A(n_1987),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2008),
.B(n_1646),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2121),
.B(n_1482),
.Y(n_2329)
);

BUFx3_ASAP7_75t_L g2330 ( 
.A(n_1964),
.Y(n_2330)
);

NAND2x1p5_ASAP7_75t_L g2331 ( 
.A(n_1971),
.B(n_1660),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1980),
.B(n_1660),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1991),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2101),
.B(n_1492),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2023),
.B(n_1715),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2134),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_2121),
.B(n_1503),
.Y(n_2337)
);

INVx6_ASAP7_75t_L g2338 ( 
.A(n_2104),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2023),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2133),
.Y(n_2340)
);

AND2x6_ASAP7_75t_L g2341 ( 
.A(n_2173),
.B(n_1503),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1955),
.B(n_1508),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_SL g2343 ( 
.A(n_2161),
.B(n_1552),
.Y(n_2343)
);

INVx4_ASAP7_75t_L g2344 ( 
.A(n_1987),
.Y(n_2344)
);

AO22x2_ASAP7_75t_L g2345 ( 
.A1(n_2200),
.A2(n_1734),
.B1(n_1934),
.B2(n_1922),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_SL g2346 ( 
.A1(n_2093),
.A2(n_1864),
.B1(n_1858),
.B2(n_1703),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2100),
.Y(n_2347)
);

INVxp33_ASAP7_75t_L g2348 ( 
.A(n_2068),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2005),
.B(n_1508),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2134),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2107),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2107),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1956),
.B(n_1511),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1959),
.B(n_1511),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2075),
.Y(n_2355)
);

INVx1_ASAP7_75t_SL g2356 ( 
.A(n_2090),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2067),
.B(n_1729),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_1987),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2136),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2138),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2138),
.Y(n_2361)
);

BUFx2_ASAP7_75t_L g2362 ( 
.A(n_2108),
.Y(n_2362)
);

AO22x2_ASAP7_75t_L g2363 ( 
.A1(n_2194),
.A2(n_1706),
.B1(n_1746),
.B2(n_1729),
.Y(n_2363)
);

CKINVDCx14_ASAP7_75t_R g2364 ( 
.A(n_2108),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2139),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2111),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2139),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2120),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_2075),
.Y(n_2369)
);

A2O1A1Ixp33_ASAP7_75t_L g2370 ( 
.A1(n_2152),
.A2(n_1634),
.B(n_1509),
.C(n_1517),
.Y(n_2370)
);

INVx4_ASAP7_75t_L g2371 ( 
.A(n_1961),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2005),
.B(n_1514),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2101),
.B(n_1514),
.Y(n_2373)
);

INVx8_ASAP7_75t_L g2374 ( 
.A(n_2075),
.Y(n_2374)
);

INVx3_ASAP7_75t_L g2375 ( 
.A(n_1971),
.Y(n_2375)
);

INVx8_ASAP7_75t_L g2376 ( 
.A(n_2075),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1962),
.B(n_1517),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2085),
.B(n_1748),
.Y(n_2378)
);

INVx4_ASAP7_75t_L g2379 ( 
.A(n_1961),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2029),
.B(n_1553),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2120),
.Y(n_2381)
);

NAND2xp33_ASAP7_75t_L g2382 ( 
.A(n_1966),
.B(n_1706),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2063),
.B(n_1553),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2137),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2211),
.B(n_1765),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2111),
.Y(n_2386)
);

NAND2x1p5_ASAP7_75t_L g2387 ( 
.A(n_2151),
.B(n_1553),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2137),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2016),
.Y(n_2389)
);

BUFx2_ASAP7_75t_L g2390 ( 
.A(n_2090),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2092),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2119),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2016),
.Y(n_2393)
);

INVxp67_ASAP7_75t_SL g2394 ( 
.A(n_2024),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2047),
.B(n_1555),
.Y(n_2395)
);

AOI22x1_ASAP7_75t_L g2396 ( 
.A1(n_2176),
.A2(n_1748),
.B1(n_1769),
.B2(n_1753),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2024),
.B(n_1555),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2211),
.B(n_1772),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2020),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2020),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2129),
.B(n_1964),
.Y(n_2401)
);

AND2x6_ASAP7_75t_L g2402 ( 
.A(n_2189),
.B(n_1533),
.Y(n_2402)
);

INVx1_ASAP7_75t_SL g2403 ( 
.A(n_2125),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2119),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2055),
.Y(n_2405)
);

INVx3_ASAP7_75t_L g2406 ( 
.A(n_1969),
.Y(n_2406)
);

NOR2x1p5_ASAP7_75t_L g2407 ( 
.A(n_2153),
.B(n_1552),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2026),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2057),
.Y(n_2409)
);

BUFx3_ASAP7_75t_L g2410 ( 
.A(n_2165),
.Y(n_2410)
);

INVxp67_ASAP7_75t_SL g2411 ( 
.A(n_2027),
.Y(n_2411)
);

AOI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2054),
.A2(n_1703),
.B1(n_1579),
.B2(n_1587),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2026),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2058),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2027),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2080),
.A2(n_1596),
.B1(n_1603),
.B2(n_1550),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2178),
.B(n_1783),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2032),
.B(n_2033),
.Y(n_2418)
);

OAI22xp5_ASAP7_75t_L g2419 ( 
.A1(n_1965),
.A2(n_1769),
.B1(n_1773),
.B2(n_1753),
.Y(n_2419)
);

INVx3_ASAP7_75t_L g2420 ( 
.A(n_1969),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2097),
.Y(n_2421)
);

CKINVDCx20_ASAP7_75t_R g2422 ( 
.A(n_2132),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2040),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2178),
.B(n_1784),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2059),
.Y(n_2425)
);

NAND2x1_ASAP7_75t_L g2426 ( 
.A(n_1966),
.B(n_1408),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2040),
.B(n_1555),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2046),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_1969),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2046),
.B(n_1604),
.Y(n_2430)
);

AOI22x1_ASAP7_75t_L g2431 ( 
.A1(n_2176),
.A2(n_2179),
.B1(n_2144),
.B2(n_2180),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2050),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2059),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2097),
.Y(n_2434)
);

AND2x4_ASAP7_75t_L g2435 ( 
.A(n_2123),
.B(n_1528),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2050),
.Y(n_2436)
);

AND2x4_ASAP7_75t_L g2437 ( 
.A(n_2184),
.B(n_1528),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_L g2438 ( 
.A1(n_1972),
.A2(n_1779),
.B1(n_1780),
.B2(n_1773),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2060),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2078),
.A2(n_1589),
.B1(n_1602),
.B2(n_1574),
.Y(n_2440)
);

O2A1O1Ixp33_ASAP7_75t_L g2441 ( 
.A1(n_2246),
.A2(n_2217),
.B(n_2131),
.C(n_2034),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2298),
.B(n_2143),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2336),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2258),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2350),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2394),
.B(n_2209),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2394),
.B(n_2209),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2411),
.B(n_2015),
.Y(n_2448)
);

A2O1A1Ixp33_ASAP7_75t_L g2449 ( 
.A1(n_2246),
.A2(n_2222),
.B(n_2088),
.C(n_2072),
.Y(n_2449)
);

OR2x6_ASAP7_75t_L g2450 ( 
.A(n_2374),
.B(n_2376),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2289),
.B(n_2004),
.Y(n_2451)
);

NAND2x1p5_ASAP7_75t_L g2452 ( 
.A(n_2371),
.B(n_2151),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2411),
.B(n_2145),
.Y(n_2453)
);

INVx4_ASAP7_75t_L g2454 ( 
.A(n_2374),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2348),
.B(n_2004),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2359),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2241),
.A2(n_2039),
.B1(n_1957),
.B2(n_2135),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2342),
.B(n_2146),
.Y(n_2458)
);

NOR2xp67_ASAP7_75t_L g2459 ( 
.A(n_2230),
.B(n_2161),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2348),
.B(n_2004),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2342),
.B(n_2156),
.Y(n_2461)
);

AOI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_2241),
.A2(n_2132),
.B1(n_1981),
.B2(n_1985),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2360),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_2421),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2340),
.B(n_2182),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2361),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2353),
.B(n_2204),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2356),
.B(n_2261),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2229),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2264),
.A2(n_2074),
.B(n_2017),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2365),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_SL g2472 ( 
.A(n_2253),
.B(n_2190),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2238),
.B(n_2390),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2421),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2385),
.A2(n_2188),
.B1(n_2126),
.B2(n_2116),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_2385),
.A2(n_2189),
.B1(n_2221),
.B2(n_2219),
.Y(n_2476)
);

INVx4_ASAP7_75t_L g2477 ( 
.A(n_2374),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2354),
.B(n_2096),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2378),
.B(n_2056),
.Y(n_2479)
);

INVx5_ASAP7_75t_L g2480 ( 
.A(n_2224),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2232),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2398),
.B(n_2056),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2367),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2398),
.B(n_2056),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2377),
.B(n_2202),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2290),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2239),
.Y(n_2487)
);

NOR2x1p5_ASAP7_75t_L g2488 ( 
.A(n_2227),
.B(n_2153),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2258),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2279),
.B(n_2300),
.C(n_2280),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2290),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2290),
.Y(n_2492)
);

NAND2x1p5_ASAP7_75t_L g2493 ( 
.A(n_2371),
.B(n_2151),
.Y(n_2493)
);

AOI22xp33_ASAP7_75t_L g2494 ( 
.A1(n_2417),
.A2(n_2221),
.B1(n_2219),
.B2(n_2022),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2266),
.B(n_2183),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2266),
.B(n_2199),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2269),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2391),
.B(n_2073),
.Y(n_2498)
);

NAND3xp33_ASAP7_75t_L g2499 ( 
.A(n_2279),
.B(n_2198),
.C(n_2030),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2391),
.B(n_2195),
.Y(n_2500)
);

AOI22xp5_ASAP7_75t_L g2501 ( 
.A1(n_2417),
.A2(n_2154),
.B1(n_2212),
.B2(n_2148),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2424),
.A2(n_2219),
.B1(n_2186),
.B2(n_2019),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2288),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2228),
.B(n_2182),
.Y(n_2504)
);

AOI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_2303),
.A2(n_2219),
.B1(n_2186),
.B2(n_2175),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_L g2506 ( 
.A(n_2225),
.B(n_2103),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2321),
.A2(n_2219),
.B1(n_2186),
.B2(n_2208),
.Y(n_2507)
);

NOR2xp67_ASAP7_75t_L g2508 ( 
.A(n_2339),
.B(n_2177),
.Y(n_2508)
);

NOR2x2_ASAP7_75t_L g2509 ( 
.A(n_2274),
.B(n_2203),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2308),
.B(n_2203),
.Y(n_2510)
);

INVx6_ASAP7_75t_L g2511 ( 
.A(n_2376),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2271),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2243),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2308),
.B(n_2206),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2224),
.Y(n_2515)
);

AOI22xp5_ASAP7_75t_L g2516 ( 
.A1(n_2280),
.A2(n_2193),
.B1(n_2191),
.B2(n_2185),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2225),
.B(n_2103),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2272),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2267),
.B(n_2156),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2321),
.A2(n_2326),
.B1(n_2346),
.B2(n_2228),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2247),
.B(n_2103),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2373),
.B(n_2115),
.Y(n_2522)
);

AND2x4_ASAP7_75t_L g2523 ( 
.A(n_2401),
.B(n_1996),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2267),
.B(n_2159),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2357),
.B(n_1705),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2251),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2262),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2373),
.B(n_2127),
.Y(n_2528)
);

AOI22xp5_ASAP7_75t_L g2529 ( 
.A1(n_2265),
.A2(n_2036),
.B1(n_1984),
.B2(n_2062),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2339),
.B(n_2182),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2335),
.B(n_1705),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2281),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2278),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2292),
.B(n_2250),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2285),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_SL g2536 ( 
.A(n_2343),
.B(n_2168),
.Y(n_2536)
);

OAI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2292),
.A2(n_2218),
.B1(n_2438),
.B2(n_2419),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2250),
.B(n_2159),
.Y(n_2538)
);

BUFx3_ASAP7_75t_L g2539 ( 
.A(n_2330),
.Y(n_2539)
);

AOI22xp33_ASAP7_75t_L g2540 ( 
.A1(n_2274),
.A2(n_2208),
.B1(n_2214),
.B2(n_2207),
.Y(n_2540)
);

BUFx8_ASAP7_75t_L g2541 ( 
.A(n_2309),
.Y(n_2541)
);

OR2x2_ASAP7_75t_L g2542 ( 
.A(n_2403),
.B(n_2215),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2270),
.B(n_2144),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2287),
.Y(n_2544)
);

AOI22xp5_ASAP7_75t_SL g2545 ( 
.A1(n_2422),
.A2(n_1881),
.B1(n_1920),
.B2(n_1874),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2270),
.B(n_2053),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2275),
.B(n_2053),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2275),
.B(n_1994),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_2421),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2283),
.Y(n_2550)
);

NAND2x1p5_ASAP7_75t_L g2551 ( 
.A(n_2379),
.B(n_2151),
.Y(n_2551)
);

INVx8_ASAP7_75t_L g2552 ( 
.A(n_2376),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2293),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2319),
.B(n_1995),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2345),
.B(n_1997),
.Y(n_2555)
);

INVx4_ASAP7_75t_L g2556 ( 
.A(n_2421),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2265),
.B(n_2205),
.Y(n_2557)
);

NAND2xp33_ASAP7_75t_L g2558 ( 
.A(n_2313),
.B(n_1966),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2286),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2299),
.A2(n_2218),
.B1(n_2160),
.B2(n_2095),
.Y(n_2560)
);

AND2x6_ASAP7_75t_SL g2561 ( 
.A(n_2401),
.B(n_2168),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2223),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2301),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2437),
.B(n_2345),
.Y(n_2564)
);

O2A1O1Ixp33_ASAP7_75t_L g2565 ( 
.A1(n_2334),
.A2(n_2124),
.B(n_2216),
.C(n_1833),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2345),
.B(n_2010),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2395),
.B(n_2163),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2434),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2434),
.B(n_2205),
.Y(n_2569)
);

O2A1O1Ixp5_ASAP7_75t_L g2570 ( 
.A1(n_2380),
.A2(n_1970),
.B(n_1982),
.C(n_2179),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2234),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2395),
.B(n_2163),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2242),
.A2(n_2259),
.B1(n_2274),
.B2(n_2435),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2329),
.B(n_2061),
.Y(n_2574)
);

INVx2_ASAP7_75t_SL g2575 ( 
.A(n_2278),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2337),
.B(n_2147),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2434),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2363),
.B(n_2147),
.Y(n_2578)
);

A2O1A1Ixp33_ASAP7_75t_L g2579 ( 
.A1(n_2412),
.A2(n_2122),
.B(n_2201),
.C(n_1979),
.Y(n_2579)
);

OAI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2363),
.A2(n_2160),
.B1(n_2396),
.B2(n_2418),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2349),
.B(n_2157),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2434),
.B(n_2205),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2304),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2349),
.B(n_2157),
.Y(n_2584)
);

A2O1A1Ixp33_ASAP7_75t_SL g2585 ( 
.A1(n_2364),
.A2(n_2167),
.B(n_2150),
.C(n_2169),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2362),
.B(n_2210),
.Y(n_2586)
);

INVx2_ASAP7_75t_SL g2587 ( 
.A(n_2330),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_2355),
.B(n_2168),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2364),
.Y(n_2589)
);

AND2x6_ASAP7_75t_SL g2590 ( 
.A(n_2422),
.B(n_1961),
.Y(n_2590)
);

BUFx2_ASAP7_75t_L g2591 ( 
.A(n_2276),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2418),
.B(n_2166),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2431),
.B(n_2166),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2368),
.B(n_2208),
.Y(n_2594)
);

O2A1O1Ixp33_ASAP7_75t_L g2595 ( 
.A1(n_2382),
.A2(n_1801),
.B(n_1825),
.C(n_1793),
.Y(n_2595)
);

BUFx2_ASAP7_75t_L g2596 ( 
.A(n_2276),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2381),
.B(n_2208),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2372),
.B(n_2210),
.Y(n_2598)
);

NOR3xp33_ASAP7_75t_L g2599 ( 
.A(n_2264),
.B(n_1799),
.C(n_2035),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2389),
.B(n_2049),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2384),
.B(n_1988),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2242),
.A2(n_2210),
.B1(n_2097),
.B2(n_2104),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2388),
.B(n_1988),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2305),
.Y(n_2604)
);

INVxp67_ASAP7_75t_L g2605 ( 
.A(n_2410),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2415),
.B(n_1988),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2315),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2236),
.Y(n_2608)
);

OR2x6_ASAP7_75t_L g2609 ( 
.A(n_2450),
.B(n_2379),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2562),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2583),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2571),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2457),
.B(n_2323),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_2503),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2541),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2539),
.Y(n_2616)
);

INVxp67_ASAP7_75t_L g2617 ( 
.A(n_2468),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_2541),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2480),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2480),
.Y(n_2620)
);

INVx3_ASAP7_75t_L g2621 ( 
.A(n_2480),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2608),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2550),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2604),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2442),
.B(n_2259),
.Y(n_2625)
);

NAND2x1p5_ASAP7_75t_L g2626 ( 
.A(n_2480),
.B(n_2224),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2607),
.Y(n_2627)
);

INVx3_ASAP7_75t_L g2628 ( 
.A(n_2452),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2444),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2552),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2559),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2490),
.A2(n_1808),
.B1(n_1813),
.B2(n_1791),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2489),
.Y(n_2633)
);

OAI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2462),
.A2(n_1961),
.B1(n_2440),
.B2(n_2162),
.Y(n_2634)
);

BUFx2_ASAP7_75t_L g2635 ( 
.A(n_2589),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2482),
.A2(n_2407),
.B1(n_2402),
.B2(n_2277),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2467),
.B(n_2317),
.Y(n_2637)
);

INVx5_ASAP7_75t_L g2638 ( 
.A(n_2450),
.Y(n_2638)
);

INVx5_ASAP7_75t_L g2639 ( 
.A(n_2450),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2542),
.B(n_2393),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2443),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2445),
.Y(n_2642)
);

INVx4_ASAP7_75t_L g2643 ( 
.A(n_2552),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2452),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2588),
.B(n_2231),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_2552),
.Y(n_2646)
);

BUFx4f_ASAP7_75t_L g2647 ( 
.A(n_2511),
.Y(n_2647)
);

BUFx3_ASAP7_75t_L g2648 ( 
.A(n_2511),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2493),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2478),
.B(n_2318),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2456),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2458),
.B(n_2383),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_2533),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2458),
.B(n_2383),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2463),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2466),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_2464),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2476),
.A2(n_2097),
.B1(n_2041),
.B2(n_2338),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2485),
.B(n_2320),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2464),
.Y(n_2660)
);

AOI22xp33_ASAP7_75t_L g2661 ( 
.A1(n_2537),
.A2(n_1813),
.B1(n_1826),
.B2(n_1808),
.Y(n_2661)
);

CKINVDCx16_ASAP7_75t_R g2662 ( 
.A(n_2472),
.Y(n_2662)
);

BUFx3_ASAP7_75t_L g2663 ( 
.A(n_2511),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2484),
.A2(n_2402),
.B1(n_2309),
.B2(n_2310),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2471),
.Y(n_2665)
);

INVx1_ASAP7_75t_SL g2666 ( 
.A(n_2479),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2483),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2497),
.Y(n_2668)
);

AND2x4_ASAP7_75t_L g2669 ( 
.A(n_2588),
.B(n_2231),
.Y(n_2669)
);

NOR3xp33_ASAP7_75t_SL g2670 ( 
.A(n_2455),
.B(n_2460),
.C(n_2451),
.Y(n_2670)
);

AND2x4_ASAP7_75t_L g2671 ( 
.A(n_2454),
.B(n_2235),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_R g2672 ( 
.A(n_2536),
.B(n_2355),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2512),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2498),
.B(n_2333),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2501),
.B(n_2224),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_2464),
.Y(n_2676)
);

INVx5_ASAP7_75t_L g2677 ( 
.A(n_2561),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2518),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2454),
.B(n_2235),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2522),
.B(n_2496),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2535),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2461),
.B(n_2399),
.Y(n_2682)
);

NAND2x1p5_ASAP7_75t_L g2683 ( 
.A(n_2477),
.B(n_2263),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2544),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2553),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2563),
.Y(n_2686)
);

BUFx6f_ASAP7_75t_L g2687 ( 
.A(n_2474),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2600),
.Y(n_2688)
);

INVxp33_ASAP7_75t_L g2689 ( 
.A(n_2528),
.Y(n_2689)
);

CKINVDCx20_ASAP7_75t_R g2690 ( 
.A(n_2591),
.Y(n_2690)
);

INVx2_ASAP7_75t_SL g2691 ( 
.A(n_2575),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2441),
.B(n_2263),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2477),
.B(n_2355),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2469),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2481),
.Y(n_2695)
);

BUFx6f_ASAP7_75t_L g2696 ( 
.A(n_2474),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2461),
.B(n_2400),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_2474),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2473),
.A2(n_2402),
.B1(n_2104),
.B2(n_2382),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2487),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2537),
.A2(n_1826),
.B1(n_2187),
.B2(n_2160),
.Y(n_2701)
);

INVx4_ASAP7_75t_L g2702 ( 
.A(n_2549),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2525),
.B(n_2564),
.Y(n_2703)
);

INVx3_ASAP7_75t_L g2704 ( 
.A(n_2549),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2513),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2499),
.A2(n_2160),
.B1(n_2413),
.B2(n_2408),
.Y(n_2706)
);

INVx4_ASAP7_75t_L g2707 ( 
.A(n_2549),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2523),
.B(n_2355),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2526),
.Y(n_2709)
);

A2O1A1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2475),
.A2(n_2449),
.B(n_2516),
.C(n_2595),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2527),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2532),
.Y(n_2712)
);

BUFx3_ASAP7_75t_L g2713 ( 
.A(n_2587),
.Y(n_2713)
);

BUFx4f_ASAP7_75t_L g2714 ( 
.A(n_2523),
.Y(n_2714)
);

INVx5_ASAP7_75t_L g2715 ( 
.A(n_2568),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2508),
.B(n_2263),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2493),
.Y(n_2717)
);

INVx3_ASAP7_75t_L g2718 ( 
.A(n_2551),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2495),
.B(n_2375),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2494),
.B(n_2263),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2581),
.B(n_2375),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2568),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2568),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2601),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2448),
.B(n_2291),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2601),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2500),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_2596),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2584),
.B(n_2311),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2574),
.B(n_2322),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2603),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2576),
.B(n_2325),
.Y(n_2732)
);

BUFx3_ASAP7_75t_L g2733 ( 
.A(n_2577),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2557),
.B(n_2369),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_R g2735 ( 
.A(n_2590),
.B(n_2369),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2577),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2504),
.B(n_2369),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2551),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2603),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2606),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2586),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2606),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2486),
.Y(n_2743)
);

BUFx4f_ASAP7_75t_L g2744 ( 
.A(n_2577),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2546),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2546),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2547),
.Y(n_2747)
);

BUFx3_ASAP7_75t_L g2748 ( 
.A(n_2530),
.Y(n_2748)
);

OR2x6_ASAP7_75t_SL g2749 ( 
.A(n_2555),
.B(n_2226),
.Y(n_2749)
);

INVxp67_ASAP7_75t_SL g2750 ( 
.A(n_2453),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2594),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2515),
.Y(n_2752)
);

BUFx3_ASAP7_75t_L g2753 ( 
.A(n_2515),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2538),
.B(n_2347),
.Y(n_2754)
);

AOI22xp33_ASAP7_75t_L g2755 ( 
.A1(n_2599),
.A2(n_2507),
.B1(n_2502),
.B2(n_2566),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2556),
.Y(n_2756)
);

BUFx2_ASAP7_75t_L g2757 ( 
.A(n_2488),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2510),
.B(n_2351),
.Y(n_2758)
);

INVx5_ASAP7_75t_L g2759 ( 
.A(n_2556),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2448),
.B(n_2453),
.Y(n_2760)
);

AND2x4_ASAP7_75t_L g2761 ( 
.A(n_2514),
.B(n_2369),
.Y(n_2761)
);

AND2x4_ASAP7_75t_L g2762 ( 
.A(n_2598),
.B(n_2254),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2491),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2529),
.B(n_2291),
.Y(n_2764)
);

BUFx2_ASAP7_75t_L g2765 ( 
.A(n_2605),
.Y(n_2765)
);

OAI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2540),
.A2(n_2338),
.B1(n_2012),
.B2(n_2213),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2492),
.Y(n_2767)
);

INVx3_ASAP7_75t_L g2768 ( 
.A(n_2446),
.Y(n_2768)
);

OAI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2520),
.A2(n_2338),
.B1(n_2169),
.B2(n_2171),
.Y(n_2769)
);

BUFx3_ASAP7_75t_L g2770 ( 
.A(n_2602),
.Y(n_2770)
);

BUFx6f_ASAP7_75t_L g2771 ( 
.A(n_2594),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2597),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2548),
.B(n_2352),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2569),
.B(n_2254),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2543),
.B(n_2366),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_L g2776 ( 
.A(n_2519),
.B(n_2302),
.Y(n_2776)
);

AND3x2_ASAP7_75t_SL g2777 ( 
.A(n_2509),
.B(n_2295),
.C(n_2386),
.Y(n_2777)
);

BUFx5_ASAP7_75t_L g2778 ( 
.A(n_2558),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2642),
.Y(n_2779)
);

INVx4_ASAP7_75t_L g2780 ( 
.A(n_2620),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2703),
.B(n_2531),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2614),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2680),
.B(n_2506),
.Y(n_2783)
);

AOI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2710),
.A2(n_2130),
.B(n_2470),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2642),
.Y(n_2785)
);

OAI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2613),
.A2(n_2579),
.B(n_2570),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2651),
.Y(n_2787)
);

NAND2xp33_ASAP7_75t_SL g2788 ( 
.A(n_2672),
.B(n_2519),
.Y(n_2788)
);

BUFx8_ASAP7_75t_SL g2789 ( 
.A(n_2615),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2651),
.Y(n_2790)
);

INVx6_ASAP7_75t_L g2791 ( 
.A(n_2662),
.Y(n_2791)
);

OAI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2689),
.A2(n_2573),
.B1(n_2505),
.B2(n_2521),
.Y(n_2792)
);

AO21x1_ASAP7_75t_L g2793 ( 
.A1(n_2692),
.A2(n_2580),
.B(n_2565),
.Y(n_2793)
);

AOI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2770),
.A2(n_2402),
.B1(n_2465),
.B2(n_2233),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_L g2795 ( 
.A(n_2689),
.B(n_2517),
.Y(n_2795)
);

OAI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2661),
.A2(n_2524),
.B1(n_2545),
.B2(n_2578),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2670),
.B(n_2554),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2750),
.B(n_2543),
.Y(n_2798)
);

INVx2_ASAP7_75t_SL g2799 ( 
.A(n_2616),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2656),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2614),
.B(n_2459),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2760),
.A2(n_2130),
.B(n_2567),
.Y(n_2802)
);

OR2x6_ASAP7_75t_SL g2803 ( 
.A(n_2615),
.B(n_2580),
.Y(n_2803)
);

OAI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_2661),
.A2(n_2524),
.B1(n_2447),
.B2(n_2534),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2632),
.A2(n_2447),
.B1(n_2534),
.B2(n_2560),
.Y(n_2805)
);

AOI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2636),
.A2(n_2582),
.B1(n_2313),
.B2(n_2284),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2727),
.B(n_2592),
.Y(n_2807)
);

AOI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2760),
.A2(n_2692),
.B(n_2572),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2664),
.A2(n_2313),
.B1(n_2284),
.B2(n_2341),
.Y(n_2809)
);

BUFx8_ASAP7_75t_L g2810 ( 
.A(n_2633),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2666),
.B(n_2358),
.Y(n_2811)
);

NOR2xp67_ASAP7_75t_SL g2812 ( 
.A(n_2638),
.B(n_2151),
.Y(n_2812)
);

CKINVDCx8_ASAP7_75t_R g2813 ( 
.A(n_2618),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2764),
.A2(n_2650),
.B(n_2659),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2656),
.Y(n_2815)
);

AND2x4_ASAP7_75t_L g2816 ( 
.A(n_2748),
.B(n_2597),
.Y(n_2816)
);

O2A1O1Ixp33_ASAP7_75t_L g2817 ( 
.A1(n_2634),
.A2(n_2585),
.B(n_2560),
.C(n_2593),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2665),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2741),
.B(n_2255),
.Y(n_2819)
);

OR2x6_ASAP7_75t_SL g2820 ( 
.A(n_2618),
.B(n_2307),
.Y(n_2820)
);

OAI21x1_ASAP7_75t_L g2821 ( 
.A1(n_2675),
.A2(n_2273),
.B(n_2268),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2625),
.B(n_2237),
.Y(n_2822)
);

AOI21x1_ASAP7_75t_L g2823 ( 
.A1(n_2716),
.A2(n_2332),
.B(n_2316),
.Y(n_2823)
);

OAI22x1_ASAP7_75t_L g2824 ( 
.A1(n_2677),
.A2(n_2244),
.B1(n_2248),
.B2(n_2240),
.Y(n_2824)
);

NAND2xp33_ASAP7_75t_L g2825 ( 
.A(n_2672),
.B(n_2313),
.Y(n_2825)
);

NOR2xp67_ASAP7_75t_L g2826 ( 
.A(n_2617),
.B(n_2256),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2665),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2667),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2637),
.B(n_2249),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2748),
.Y(n_2830)
);

AND2x4_ASAP7_75t_L g2831 ( 
.A(n_2645),
.B(n_2306),
.Y(n_2831)
);

BUFx8_ASAP7_75t_SL g2832 ( 
.A(n_2690),
.Y(n_2832)
);

INVx1_ASAP7_75t_SL g2833 ( 
.A(n_2640),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2667),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2668),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2688),
.B(n_2392),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2652),
.A2(n_2332),
.B(n_2181),
.Y(n_2837)
);

O2A1O1Ixp5_ASAP7_75t_SL g2838 ( 
.A1(n_2716),
.A2(n_2257),
.B(n_2260),
.C(n_2252),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2668),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2652),
.A2(n_2181),
.B(n_2282),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2769),
.A2(n_2341),
.B1(n_2233),
.B2(n_1574),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2647),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2761),
.B(n_2404),
.Y(n_2843)
);

INVx5_ASAP7_75t_L g2844 ( 
.A(n_2609),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2728),
.Y(n_2845)
);

OAI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2654),
.A2(n_2416),
.B(n_2370),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_SL g2847 ( 
.A(n_2677),
.B(n_2291),
.Y(n_2847)
);

AOI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2654),
.A2(n_2314),
.B(n_2282),
.Y(n_2848)
);

AOI22x1_ASAP7_75t_L g2849 ( 
.A1(n_2757),
.A2(n_2327),
.B1(n_2344),
.B2(n_2294),
.Y(n_2849)
);

NOR2xp33_ASAP7_75t_L g2850 ( 
.A(n_2635),
.B(n_2327),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2632),
.A2(n_2291),
.B1(n_2428),
.B2(n_2423),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2761),
.B(n_2405),
.Y(n_2852)
);

INVx3_ASAP7_75t_L g2853 ( 
.A(n_2702),
.Y(n_2853)
);

AOI211xp5_ASAP7_75t_SL g2854 ( 
.A1(n_2658),
.A2(n_1878),
.B(n_1886),
.C(n_1877),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2674),
.B(n_2432),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2701),
.A2(n_2436),
.B1(n_2172),
.B2(n_2427),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2755),
.A2(n_2341),
.B1(n_2233),
.B2(n_1589),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2682),
.A2(n_2324),
.B(n_2314),
.Y(n_2858)
);

HB1xp67_ASAP7_75t_L g2859 ( 
.A(n_2771),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2770),
.A2(n_2233),
.B1(n_2341),
.B2(n_2197),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2697),
.A2(n_2328),
.B(n_2324),
.Y(n_2861)
);

A2O1A1Ixp33_ASAP7_75t_L g2862 ( 
.A1(n_2755),
.A2(n_2164),
.B(n_2171),
.C(n_2169),
.Y(n_2862)
);

OAI22xp5_ASAP7_75t_SL g2863 ( 
.A1(n_2690),
.A2(n_2306),
.B1(n_2312),
.B2(n_2344),
.Y(n_2863)
);

O2A1O1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2720),
.A2(n_2370),
.B(n_2042),
.C(n_2167),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2765),
.B(n_2306),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2725),
.A2(n_2031),
.B(n_2426),
.Y(n_2866)
);

AOI22xp5_ASAP7_75t_L g2867 ( 
.A1(n_2677),
.A2(n_2699),
.B1(n_2728),
.B2(n_2714),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2720),
.A2(n_2197),
.B(n_2245),
.Y(n_2868)
);

BUFx8_ASAP7_75t_SL g2869 ( 
.A(n_2629),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2771),
.Y(n_2870)
);

O2A1O1Ixp33_ASAP7_75t_L g2871 ( 
.A1(n_2766),
.A2(n_2167),
.B(n_2150),
.C(n_2164),
.Y(n_2871)
);

INVx5_ASAP7_75t_L g2872 ( 
.A(n_2609),
.Y(n_2872)
);

INVx3_ASAP7_75t_L g2873 ( 
.A(n_2702),
.Y(n_2873)
);

OAI21xp33_ASAP7_75t_SL g2874 ( 
.A1(n_2706),
.A2(n_2245),
.B(n_2397),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2730),
.B(n_2768),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2768),
.B(n_2719),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2706),
.A2(n_2172),
.B1(n_2427),
.B2(n_2397),
.Y(n_2877)
);

AOI21x1_ASAP7_75t_L g2878 ( 
.A1(n_2775),
.A2(n_1943),
.B(n_2052),
.Y(n_2878)
);

OAI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2749),
.A2(n_2406),
.B1(n_2429),
.B2(n_2420),
.Y(n_2879)
);

O2A1O1Ixp33_ASAP7_75t_SL g2880 ( 
.A1(n_2754),
.A2(n_2691),
.B(n_2653),
.C(n_2773),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2745),
.B(n_2746),
.Y(n_2881)
);

AOI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2714),
.A2(n_2174),
.B(n_2430),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2645),
.B(n_2409),
.Y(n_2883)
);

INVxp67_ASAP7_75t_L g2884 ( 
.A(n_2713),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_SL g2885 ( 
.A(n_2647),
.B(n_2638),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2708),
.A2(n_2233),
.B1(n_1602),
.B2(n_1499),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2645),
.B(n_2414),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2746),
.A2(n_2174),
.B(n_2430),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2669),
.B(n_2623),
.Y(n_2889)
);

AND2x4_ASAP7_75t_L g2890 ( 
.A(n_2669),
.B(n_2312),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2669),
.B(n_2425),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2616),
.B(n_2312),
.Y(n_2892)
);

NOR2xp67_ASAP7_75t_L g2893 ( 
.A(n_2694),
.B(n_2695),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2681),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2685),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2747),
.B(n_2433),
.Y(n_2896)
);

OA22x2_ASAP7_75t_L g2897 ( 
.A1(n_2734),
.A2(n_2439),
.B1(n_2079),
.B2(n_2081),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2735),
.B(n_2312),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2735),
.B(n_2076),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2713),
.B(n_2083),
.Y(n_2900)
);

AOI21xp33_ASAP7_75t_L g2901 ( 
.A1(n_2776),
.A2(n_2051),
.B(n_2102),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2611),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2638),
.A2(n_2051),
.B(n_2296),
.Y(n_2903)
);

BUFx2_ASAP7_75t_L g2904 ( 
.A(n_2722),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2729),
.B(n_1546),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2732),
.B(n_1546),
.Y(n_2906)
);

O2A1O1Ixp33_ASAP7_75t_L g2907 ( 
.A1(n_2624),
.A2(n_2038),
.B(n_2045),
.C(n_2037),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2722),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2708),
.B(n_1499),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2758),
.B(n_1549),
.Y(n_2910)
);

O2A1O1Ixp33_ASAP7_75t_L g2911 ( 
.A1(n_2627),
.A2(n_2038),
.B(n_2045),
.C(n_2037),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2685),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2708),
.B(n_1499),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_R g2914 ( 
.A(n_2630),
.B(n_1966),
.Y(n_2914)
);

INVx3_ASAP7_75t_SL g2915 ( 
.A(n_2693),
.Y(n_2915)
);

NAND3xp33_ASAP7_75t_L g2916 ( 
.A(n_2721),
.B(n_2109),
.C(n_2105),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2751),
.B(n_2772),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_L g2918 ( 
.A(n_2771),
.B(n_1554),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2609),
.B(n_2406),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2743),
.Y(n_2920)
);

OAI21xp33_ASAP7_75t_SL g2921 ( 
.A1(n_2763),
.A2(n_2429),
.B(n_2420),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2638),
.A2(n_2051),
.B(n_2296),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2767),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2772),
.B(n_1554),
.Y(n_2924)
);

NOR2xp33_ASAP7_75t_L g2925 ( 
.A(n_2771),
.B(n_1556),
.Y(n_2925)
);

O2A1O1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2641),
.A2(n_2114),
.B(n_2117),
.C(n_2110),
.Y(n_2926)
);

A2O1A1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_2762),
.A2(n_2118),
.B(n_2064),
.C(n_2087),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2639),
.A2(n_2331),
.B(n_2387),
.Y(n_2928)
);

O2A1O1Ixp5_ASAP7_75t_L g2929 ( 
.A1(n_2734),
.A2(n_1898),
.B(n_1896),
.C(n_2142),
.Y(n_2929)
);

NOR2xp67_ASAP7_75t_SL g2930 ( 
.A(n_2639),
.B(n_2060),
.Y(n_2930)
);

OAI21xp33_ASAP7_75t_SL g2931 ( 
.A1(n_2655),
.A2(n_2142),
.B(n_2087),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2639),
.A2(n_2387),
.B(n_1986),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2673),
.A2(n_2064),
.B1(n_2077),
.B2(n_2028),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2678),
.Y(n_2934)
);

O2A1O1Ixp33_ASAP7_75t_L g2935 ( 
.A1(n_2684),
.A2(n_1563),
.B(n_1556),
.C(n_1870),
.Y(n_2935)
);

OAI22xp33_ASAP7_75t_SL g2936 ( 
.A1(n_2686),
.A2(n_2028),
.B1(n_2128),
.B2(n_2077),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2737),
.B(n_1563),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2724),
.A2(n_1986),
.B(n_1966),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2724),
.A2(n_2028),
.B1(n_2128),
.B2(n_2077),
.Y(n_2939)
);

NOR2x1_ASAP7_75t_SL g2940 ( 
.A(n_2620),
.B(n_1966),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_2705),
.B(n_295),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2726),
.A2(n_2739),
.B1(n_2740),
.B2(n_2731),
.Y(n_2942)
);

BUFx6f_ASAP7_75t_L g2943 ( 
.A(n_2648),
.Y(n_2943)
);

OA22x2_ASAP7_75t_L g2944 ( 
.A1(n_2737),
.A2(n_2141),
.B1(n_2128),
.B2(n_50),
.Y(n_2944)
);

OR2x6_ASAP7_75t_L g2945 ( 
.A(n_2643),
.B(n_2726),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2798),
.B(n_2731),
.Y(n_2946)
);

OAI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2786),
.A2(n_2762),
.B(n_2740),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2779),
.Y(n_2948)
);

NAND3xp33_ASAP7_75t_L g2949 ( 
.A(n_2786),
.B(n_2712),
.C(n_2709),
.Y(n_2949)
);

AO31x2_ASAP7_75t_L g2950 ( 
.A1(n_2793),
.A2(n_2742),
.A3(n_2612),
.B(n_2622),
.Y(n_2950)
);

OAI21x1_ASAP7_75t_SL g2951 ( 
.A1(n_2814),
.A2(n_2643),
.B(n_2622),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2784),
.A2(n_2759),
.B(n_2620),
.Y(n_2952)
);

OAI21x1_ASAP7_75t_L g2953 ( 
.A1(n_2838),
.A2(n_2932),
.B(n_2878),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2920),
.Y(n_2954)
);

NOR2xp67_ASAP7_75t_SL g2955 ( 
.A(n_2813),
.B(n_2844),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2833),
.B(n_2610),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2833),
.B(n_2631),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2943),
.Y(n_2958)
);

OAI21x1_ASAP7_75t_SL g2959 ( 
.A1(n_2808),
.A2(n_2643),
.B(n_2631),
.Y(n_2959)
);

AO31x2_ASAP7_75t_L g2960 ( 
.A1(n_2824),
.A2(n_2711),
.A3(n_2700),
.B(n_2707),
.Y(n_2960)
);

NAND3xp33_ASAP7_75t_L g2961 ( 
.A(n_2797),
.B(n_2711),
.C(n_2700),
.Y(n_2961)
);

AO21x1_ASAP7_75t_L g2962 ( 
.A1(n_2788),
.A2(n_2777),
.B(n_2774),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2876),
.B(n_2774),
.Y(n_2963)
);

OAI21x1_ASAP7_75t_L g2964 ( 
.A1(n_2938),
.A2(n_2644),
.B(n_2628),
.Y(n_2964)
);

AO21x2_ASAP7_75t_L g2965 ( 
.A1(n_2901),
.A2(n_1873),
.B(n_1913),
.Y(n_2965)
);

AOI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2930),
.A2(n_2693),
.B(n_2679),
.Y(n_2966)
);

A2O1A1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2817),
.A2(n_2744),
.B(n_2663),
.C(n_2648),
.Y(n_2967)
);

INVx3_ASAP7_75t_L g2968 ( 
.A(n_2943),
.Y(n_2968)
);

BUFx2_ASAP7_75t_L g2969 ( 
.A(n_2830),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2783),
.B(n_2671),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2807),
.B(n_2778),
.Y(n_2971)
);

INVx4_ASAP7_75t_L g2972 ( 
.A(n_2943),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2923),
.Y(n_2973)
);

OAI21x1_ASAP7_75t_L g2974 ( 
.A1(n_2823),
.A2(n_2644),
.B(n_2628),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2796),
.A2(n_2620),
.B1(n_2663),
.B2(n_2626),
.Y(n_2975)
);

AND2x2_ASAP7_75t_SL g2976 ( 
.A(n_2825),
.B(n_2630),
.Y(n_2976)
);

OAI21x1_ASAP7_75t_L g2977 ( 
.A1(n_2903),
.A2(n_2717),
.B(n_2649),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2781),
.B(n_2657),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2875),
.B(n_2752),
.Y(n_2979)
);

INVx3_ASAP7_75t_L g2980 ( 
.A(n_2780),
.Y(n_2980)
);

OAI21x1_ASAP7_75t_L g2981 ( 
.A1(n_2922),
.A2(n_2717),
.B(n_2649),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2795),
.B(n_2657),
.Y(n_2982)
);

OAI21x1_ASAP7_75t_L g2983 ( 
.A1(n_2821),
.A2(n_2928),
.B(n_2866),
.Y(n_2983)
);

OAI21xp5_ASAP7_75t_SL g2984 ( 
.A1(n_2857),
.A2(n_2693),
.B(n_2683),
.Y(n_2984)
);

NAND3xp33_ASAP7_75t_SL g2985 ( 
.A(n_2899),
.B(n_2683),
.C(n_2702),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2796),
.A2(n_2621),
.B1(n_2619),
.B2(n_2715),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2934),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2785),
.Y(n_2988)
);

O2A1O1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2792),
.A2(n_2738),
.B(n_2718),
.C(n_2619),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2881),
.B(n_2660),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2816),
.B(n_2660),
.Y(n_2991)
);

AND2x2_ASAP7_75t_SL g2992 ( 
.A(n_2885),
.B(n_2630),
.Y(n_2992)
);

OAI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2803),
.A2(n_2621),
.B1(n_2619),
.B2(n_2715),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2942),
.B(n_2778),
.Y(n_2994)
);

OAI21x1_ASAP7_75t_SL g2995 ( 
.A1(n_2907),
.A2(n_2707),
.B(n_2778),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2787),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2800),
.Y(n_2997)
);

INVx1_ASAP7_75t_SL g2998 ( 
.A(n_2859),
.Y(n_2998)
);

OA21x2_ASAP7_75t_L g2999 ( 
.A1(n_2846),
.A2(n_2868),
.B(n_2802),
.Y(n_2999)
);

AO21x1_ASAP7_75t_L g3000 ( 
.A1(n_2879),
.A2(n_2819),
.B(n_2851),
.Y(n_3000)
);

AO21x1_ASAP7_75t_L g3001 ( 
.A1(n_2879),
.A2(n_2707),
.B(n_2679),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2827),
.Y(n_3002)
);

AO21x1_ASAP7_75t_L g3003 ( 
.A1(n_2851),
.A2(n_2679),
.B(n_2671),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2816),
.B(n_2698),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2889),
.B(n_2698),
.Y(n_3005)
);

OAI21x1_ASAP7_75t_L g3006 ( 
.A1(n_2864),
.A2(n_2756),
.B(n_2141),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2902),
.B(n_2704),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2791),
.B(n_2832),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2791),
.B(n_2704),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2870),
.B(n_2733),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2888),
.A2(n_2756),
.B(n_2141),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_2882),
.A2(n_2759),
.B(n_2715),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2917),
.B(n_2753),
.Y(n_3013)
);

OAI21x1_ASAP7_75t_L g3014 ( 
.A1(n_2897),
.A2(n_2756),
.B(n_1538),
.Y(n_3014)
);

OAI21x1_ASAP7_75t_L g3015 ( 
.A1(n_2897),
.A2(n_1538),
.B(n_1534),
.Y(n_3015)
);

A2O1A1Ixp33_ASAP7_75t_L g3016 ( 
.A1(n_2874),
.A2(n_2671),
.B(n_2753),
.C(n_2733),
.Y(n_3016)
);

AOI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2867),
.A2(n_2778),
.B1(n_2630),
.B2(n_2646),
.Y(n_3017)
);

BUFx2_ASAP7_75t_L g3018 ( 
.A(n_2810),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2837),
.A2(n_1539),
.B(n_1534),
.Y(n_3019)
);

OR2x2_ASAP7_75t_L g3020 ( 
.A(n_2790),
.B(n_2676),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2942),
.B(n_2778),
.Y(n_3021)
);

OAI21x1_ASAP7_75t_L g3022 ( 
.A1(n_2848),
.A2(n_1542),
.B(n_1539),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2815),
.B(n_2778),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2818),
.B(n_2676),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2835),
.Y(n_3025)
);

OAI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2862),
.A2(n_2197),
.B(n_2070),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2780),
.Y(n_3027)
);

OA21x2_ASAP7_75t_L g3028 ( 
.A1(n_2868),
.A2(n_2070),
.B(n_1986),
.Y(n_3028)
);

OR2x6_ASAP7_75t_L g3029 ( 
.A(n_2945),
.B(n_2646),
.Y(n_3029)
);

OAI21x1_ASAP7_75t_L g3030 ( 
.A1(n_2871),
.A2(n_1479),
.B(n_1446),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2839),
.B(n_2676),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2885),
.A2(n_2759),
.B(n_2715),
.Y(n_3032)
);

O2A1O1Ixp33_ASAP7_75t_L g3033 ( 
.A1(n_2880),
.A2(n_1941),
.B(n_1915),
.C(n_1905),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2894),
.B(n_2687),
.Y(n_3034)
);

BUFx6f_ASAP7_75t_L g3035 ( 
.A(n_2842),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2840),
.A2(n_2861),
.B(n_2858),
.Y(n_3036)
);

OAI21x1_ASAP7_75t_L g3037 ( 
.A1(n_2911),
.A2(n_1479),
.B(n_1446),
.Y(n_3037)
);

OAI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2916),
.A2(n_2841),
.B(n_2877),
.Y(n_3038)
);

OAI21xp5_ASAP7_75t_SL g3039 ( 
.A1(n_2809),
.A2(n_2646),
.B(n_2687),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2844),
.A2(n_2070),
.B(n_1986),
.Y(n_3040)
);

NOR2xp33_ASAP7_75t_L g3041 ( 
.A(n_2782),
.B(n_2845),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2828),
.Y(n_3042)
);

OAI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2877),
.A2(n_2113),
.B(n_2297),
.Y(n_3043)
);

NAND2x1p5_ASAP7_75t_L g3044 ( 
.A(n_2844),
.B(n_2687),
.Y(n_3044)
);

OAI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2806),
.A2(n_2113),
.B(n_2297),
.Y(n_3045)
);

AO21x1_ASAP7_75t_L g3046 ( 
.A1(n_2936),
.A2(n_48),
.B(n_49),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2844),
.A2(n_2113),
.B(n_2297),
.Y(n_3047)
);

AO31x2_ASAP7_75t_L g3048 ( 
.A1(n_2805),
.A2(n_2113),
.A3(n_2297),
.B(n_1976),
.Y(n_3048)
);

OAI21x1_ASAP7_75t_L g3049 ( 
.A1(n_2933),
.A2(n_1498),
.B(n_1446),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2834),
.Y(n_3050)
);

OAI21x1_ASAP7_75t_L g3051 ( 
.A1(n_2933),
.A2(n_1498),
.B(n_1562),
.Y(n_3051)
);

CKINVDCx5p33_ASAP7_75t_R g3052 ( 
.A(n_2789),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2872),
.B(n_2736),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2822),
.B(n_2696),
.Y(n_3054)
);

OAI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2927),
.A2(n_2297),
.B(n_1562),
.Y(n_3055)
);

O2A1O1Ixp5_ASAP7_75t_L g3056 ( 
.A1(n_2847),
.A2(n_1416),
.B(n_1408),
.C(n_2723),
.Y(n_3056)
);

NAND2xp33_ASAP7_75t_SL g3057 ( 
.A(n_2842),
.B(n_2723),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2805),
.A2(n_1562),
.B(n_1498),
.Y(n_3058)
);

AO21x1_ASAP7_75t_L g3059 ( 
.A1(n_2900),
.A2(n_51),
.B(n_52),
.Y(n_3059)
);

OAI21x1_ASAP7_75t_L g3060 ( 
.A1(n_2939),
.A2(n_1498),
.B(n_1562),
.Y(n_3060)
);

OAI21x1_ASAP7_75t_L g3061 ( 
.A1(n_2939),
.A2(n_1524),
.B(n_1416),
.Y(n_3061)
);

OAI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2804),
.A2(n_2856),
.B(n_2854),
.Y(n_3062)
);

A2O1A1Ixp33_ASAP7_75t_L g3063 ( 
.A1(n_2804),
.A2(n_2736),
.B(n_2723),
.C(n_54),
.Y(n_3063)
);

OAI21x1_ASAP7_75t_SL g3064 ( 
.A1(n_2940),
.A2(n_1524),
.B(n_2736),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_2872),
.A2(n_1976),
.B(n_1470),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2895),
.B(n_1524),
.Y(n_3066)
);

AO32x2_ASAP7_75t_L g3067 ( 
.A1(n_2856),
.A2(n_56),
.A3(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_3067)
);

AO31x2_ASAP7_75t_L g3068 ( 
.A1(n_2912),
.A2(n_2918),
.A3(n_2925),
.B(n_2829),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2872),
.A2(n_1976),
.B(n_1470),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2836),
.B(n_53),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_2801),
.B(n_56),
.Y(n_3071)
);

AOI22xp5_ASAP7_75t_L g3072 ( 
.A1(n_2909),
.A2(n_1470),
.B1(n_1474),
.B2(n_1464),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2872),
.B(n_1976),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2855),
.B(n_58),
.Y(n_3074)
);

OAI22x1_ASAP7_75t_L g3075 ( 
.A1(n_2884),
.A2(n_62),
.B1(n_58),
.B2(n_61),
.Y(n_3075)
);

A2O1A1Ixp33_ASAP7_75t_L g3076 ( 
.A1(n_2860),
.A2(n_64),
.B(n_61),
.C(n_63),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2893),
.B(n_63),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2945),
.A2(n_1470),
.B(n_1464),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2843),
.B(n_64),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2852),
.B(n_65),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_2853),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2865),
.B(n_66),
.Y(n_3082)
);

OAI21x1_ASAP7_75t_L g3083 ( 
.A1(n_2929),
.A2(n_1470),
.B(n_1464),
.Y(n_3083)
);

OAI21xp5_ASAP7_75t_L g3084 ( 
.A1(n_2886),
.A2(n_66),
.B(n_67),
.Y(n_3084)
);

OA21x2_ASAP7_75t_L g3085 ( 
.A1(n_2794),
.A2(n_68),
.B(n_69),
.Y(n_3085)
);

INVx4_ASAP7_75t_SL g3086 ( 
.A(n_2915),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2896),
.B(n_68),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2944),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_3088)
);

BUFx12f_ASAP7_75t_L g3089 ( 
.A(n_2842),
.Y(n_3089)
);

OAI21x1_ASAP7_75t_L g3090 ( 
.A1(n_2935),
.A2(n_2944),
.B(n_2924),
.Y(n_3090)
);

OR2x2_ASAP7_75t_L g3091 ( 
.A(n_2904),
.B(n_71),
.Y(n_3091)
);

OAI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2931),
.A2(n_72),
.B(n_73),
.Y(n_3092)
);

NOR2x1_ASAP7_75t_SL g3093 ( 
.A(n_2898),
.B(n_1003),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2820),
.B(n_74),
.Y(n_3094)
);

OAI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2799),
.A2(n_1478),
.B1(n_1502),
.B2(n_1474),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_L g3096 ( 
.A1(n_2863),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2811),
.B(n_77),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2850),
.A2(n_2906),
.B1(n_2910),
.B2(n_2905),
.Y(n_3098)
);

OAI21x1_ASAP7_75t_L g3099 ( 
.A1(n_2926),
.A2(n_1478),
.B(n_1474),
.Y(n_3099)
);

OAI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2921),
.A2(n_77),
.B(n_78),
.Y(n_3100)
);

OAI21x1_ASAP7_75t_L g3101 ( 
.A1(n_2937),
.A2(n_1502),
.B(n_1478),
.Y(n_3101)
);

AND2x4_ASAP7_75t_L g3102 ( 
.A(n_2919),
.B(n_296),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2919),
.A2(n_1502),
.B(n_1478),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2883),
.B(n_78),
.Y(n_3104)
);

OAI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2941),
.A2(n_2826),
.B1(n_2913),
.B2(n_2892),
.Y(n_3105)
);

INVx5_ASAP7_75t_L g3106 ( 
.A(n_2869),
.Y(n_3106)
);

INVx4_ASAP7_75t_L g3107 ( 
.A(n_2853),
.Y(n_3107)
);

NAND2x1_ASAP7_75t_L g3108 ( 
.A(n_2812),
.B(n_1502),
.Y(n_3108)
);

AOI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2831),
.A2(n_1513),
.B(n_1504),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2887),
.Y(n_3110)
);

OAI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2891),
.A2(n_80),
.B(n_81),
.Y(n_3111)
);

OAI21x1_ASAP7_75t_L g3112 ( 
.A1(n_2873),
.A2(n_1513),
.B(n_1504),
.Y(n_3112)
);

OAI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2849),
.A2(n_2873),
.B(n_2831),
.Y(n_3113)
);

OAI21x1_ASAP7_75t_L g3114 ( 
.A1(n_2914),
.A2(n_1513),
.B(n_1504),
.Y(n_3114)
);

OAI22xp5_ASAP7_75t_L g3115 ( 
.A1(n_2908),
.A2(n_84),
.B1(n_80),
.B2(n_82),
.Y(n_3115)
);

OR2x2_ASAP7_75t_L g3116 ( 
.A(n_2890),
.B(n_85),
.Y(n_3116)
);

OAI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2786),
.A2(n_85),
.B(n_86),
.Y(n_3117)
);

AO21x2_ASAP7_75t_L g3118 ( 
.A1(n_3036),
.A2(n_2953),
.B(n_3117),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_3107),
.Y(n_3119)
);

AO21x1_ASAP7_75t_L g3120 ( 
.A1(n_3088),
.A2(n_86),
.B(n_87),
.Y(n_3120)
);

A2O1A1Ixp33_ASAP7_75t_L g3121 ( 
.A1(n_3117),
.A2(n_91),
.B(n_87),
.C(n_88),
.Y(n_3121)
);

OR2x6_ASAP7_75t_L g3122 ( 
.A(n_3032),
.B(n_1003),
.Y(n_3122)
);

OAI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_3063),
.A2(n_91),
.B(n_93),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2954),
.Y(n_3124)
);

NAND3xp33_ASAP7_75t_SL g3125 ( 
.A(n_3059),
.B(n_93),
.C(n_94),
.Y(n_3125)
);

AOI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2955),
.A2(n_96),
.B(n_97),
.Y(n_3126)
);

NOR2xp33_ASAP7_75t_L g3127 ( 
.A(n_2982),
.B(n_96),
.Y(n_3127)
);

OAI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_3062),
.A2(n_97),
.B(n_98),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_SL g3129 ( 
.A(n_3098),
.B(n_3105),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_3055),
.A2(n_1513),
.B(n_1438),
.Y(n_3130)
);

AOI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_3062),
.A2(n_3088),
.B1(n_3105),
.B2(n_3084),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2973),
.Y(n_3132)
);

AO31x2_ASAP7_75t_L g3133 ( 
.A1(n_3001),
.A2(n_101),
.A3(n_99),
.B(n_100),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2963),
.B(n_100),
.Y(n_3134)
);

A2O1A1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_3084),
.A2(n_106),
.B(n_103),
.C(n_105),
.Y(n_3135)
);

OAI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2967),
.A2(n_3111),
.B(n_3100),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2969),
.B(n_103),
.Y(n_3137)
);

OAI21x1_ASAP7_75t_L g3138 ( 
.A1(n_2983),
.A2(n_302),
.B(n_301),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2946),
.B(n_107),
.Y(n_3139)
);

HB1xp67_ASAP7_75t_L g3140 ( 
.A(n_3068),
.Y(n_3140)
);

AOI221x1_ASAP7_75t_L g3141 ( 
.A1(n_3094),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.C(n_111),
.Y(n_3141)
);

CKINVDCx20_ASAP7_75t_R g3142 ( 
.A(n_3052),
.Y(n_3142)
);

AO31x2_ASAP7_75t_L g3143 ( 
.A1(n_3000),
.A2(n_112),
.A3(n_108),
.B(n_109),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_2998),
.B(n_112),
.Y(n_3144)
);

O2A1O1Ixp33_ASAP7_75t_L g3145 ( 
.A1(n_3076),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_3145)
);

A2O1A1Ixp33_ASAP7_75t_L g3146 ( 
.A1(n_3111),
.A2(n_116),
.B(n_113),
.C(n_114),
.Y(n_3146)
);

OAI21x1_ASAP7_75t_L g3147 ( 
.A1(n_3099),
.A2(n_305),
.B(n_303),
.Y(n_3147)
);

NAND3x1_ASAP7_75t_L g3148 ( 
.A(n_3008),
.B(n_116),
.C(n_117),
.Y(n_3148)
);

INVx1_ASAP7_75t_SL g3149 ( 
.A(n_3018),
.Y(n_3149)
);

O2A1O1Ixp33_ASAP7_75t_SL g3150 ( 
.A1(n_3094),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_3012),
.A2(n_1449),
.B(n_1448),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2946),
.B(n_120),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_3043),
.A2(n_1449),
.B(n_1448),
.Y(n_3153)
);

OAI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_3096),
.A2(n_1050),
.B1(n_125),
.B2(n_122),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_3043),
.A2(n_1449),
.B(n_1405),
.Y(n_3155)
);

OAI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_3100),
.A2(n_126),
.B(n_129),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2987),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2971),
.B(n_129),
.Y(n_3158)
);

A2O1A1Ixp33_ASAP7_75t_L g3159 ( 
.A1(n_2989),
.A2(n_133),
.B(n_130),
.C(n_131),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2971),
.B(n_130),
.Y(n_3160)
);

NAND3x1_ASAP7_75t_L g3161 ( 
.A(n_3041),
.B(n_133),
.C(n_134),
.Y(n_3161)
);

OAI21x1_ASAP7_75t_L g3162 ( 
.A1(n_3083),
.A2(n_314),
.B(n_313),
.Y(n_3162)
);

OAI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2949),
.A2(n_136),
.B(n_137),
.Y(n_3163)
);

AO31x2_ASAP7_75t_L g3164 ( 
.A1(n_3003),
.A2(n_136),
.A3(n_138),
.B(n_139),
.Y(n_3164)
);

INVx2_ASAP7_75t_SL g3165 ( 
.A(n_3106),
.Y(n_3165)
);

BUFx3_ASAP7_75t_L g3166 ( 
.A(n_3106),
.Y(n_3166)
);

NOR2xp33_ASAP7_75t_R g3167 ( 
.A(n_3106),
.B(n_140),
.Y(n_3167)
);

NAND3x1_ASAP7_75t_L g3168 ( 
.A(n_3017),
.B(n_140),
.C(n_141),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3025),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_3038),
.A2(n_1405),
.B(n_1050),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3042),
.Y(n_3171)
);

O2A1O1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_3115),
.A2(n_142),
.B(n_143),
.C(n_144),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2948),
.Y(n_3173)
);

OAI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2976),
.A2(n_1050),
.B1(n_143),
.B2(n_144),
.Y(n_3174)
);

AND2x2_ASAP7_75t_SL g3175 ( 
.A(n_2992),
.B(n_1050),
.Y(n_3175)
);

HB1xp67_ASAP7_75t_L g3176 ( 
.A(n_3068),
.Y(n_3176)
);

CKINVDCx16_ASAP7_75t_R g3177 ( 
.A(n_3089),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2952),
.A2(n_1405),
.B(n_145),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_3071),
.B(n_147),
.Y(n_3179)
);

INVx3_ASAP7_75t_L g3180 ( 
.A(n_3107),
.Y(n_3180)
);

AO31x2_ASAP7_75t_L g3181 ( 
.A1(n_2962),
.A2(n_3046),
.A3(n_2986),
.B(n_3047),
.Y(n_3181)
);

AOI21xp33_ASAP7_75t_L g3182 ( 
.A1(n_3098),
.A2(n_148),
.B(n_149),
.Y(n_3182)
);

NAND3xp33_ASAP7_75t_L g3183 ( 
.A(n_2961),
.B(n_148),
.C(n_149),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2956),
.B(n_2957),
.Y(n_3184)
);

NOR2xp67_ASAP7_75t_SL g3185 ( 
.A(n_3085),
.B(n_317),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2988),
.Y(n_3186)
);

AO31x2_ASAP7_75t_L g3187 ( 
.A1(n_2986),
.A2(n_150),
.A3(n_151),
.B(n_152),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2996),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_SL g3189 ( 
.A(n_2972),
.B(n_318),
.Y(n_3189)
);

INVx4_ASAP7_75t_L g3190 ( 
.A(n_3086),
.Y(n_3190)
);

AO32x2_ASAP7_75t_L g3191 ( 
.A1(n_2993),
.A2(n_150),
.A3(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_3191)
);

NAND3xp33_ASAP7_75t_L g3192 ( 
.A(n_3092),
.B(n_154),
.C(n_155),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_SL g3193 ( 
.A(n_2970),
.B(n_321),
.Y(n_3193)
);

CKINVDCx8_ASAP7_75t_R g3194 ( 
.A(n_3035),
.Y(n_3194)
);

AOI221xp5_ASAP7_75t_SL g3195 ( 
.A1(n_3075),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.C(n_162),
.Y(n_3195)
);

OAI21xp33_ASAP7_75t_SL g3196 ( 
.A1(n_3092),
.A2(n_160),
.B(n_163),
.Y(n_3196)
);

O2A1O1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_3077),
.A2(n_164),
.B(n_166),
.C(n_167),
.Y(n_3197)
);

AOI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_2975),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_3198)
);

INVx2_ASAP7_75t_SL g3199 ( 
.A(n_2958),
.Y(n_3199)
);

O2A1O1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_3016),
.A2(n_171),
.B(n_174),
.C(n_175),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_L g3201 ( 
.A1(n_3006),
.A2(n_325),
.B(n_324),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_2999),
.A2(n_174),
.B(n_176),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2999),
.A2(n_176),
.B(n_177),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_3035),
.Y(n_3204)
);

OAI22x1_ASAP7_75t_L g3205 ( 
.A1(n_3110),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2997),
.Y(n_3206)
);

OAI21x1_ASAP7_75t_L g3207 ( 
.A1(n_3019),
.A2(n_331),
.B(n_329),
.Y(n_3207)
);

INVx3_ASAP7_75t_L g3208 ( 
.A(n_2972),
.Y(n_3208)
);

AOI21x1_ASAP7_75t_L g3209 ( 
.A1(n_3053),
.A2(n_178),
.B(n_179),
.Y(n_3209)
);

HB1xp67_ASAP7_75t_L g3210 ( 
.A(n_3068),
.Y(n_3210)
);

AO31x2_ASAP7_75t_L g3211 ( 
.A1(n_2993),
.A2(n_180),
.A3(n_181),
.B(n_182),
.Y(n_3211)
);

OAI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_2985),
.A2(n_181),
.B(n_183),
.Y(n_3212)
);

OAI21x1_ASAP7_75t_L g3213 ( 
.A1(n_2974),
.A2(n_335),
.B(n_332),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_SL g3214 ( 
.A(n_2975),
.B(n_336),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_3029),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2979),
.B(n_183),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3026),
.A2(n_184),
.B(n_186),
.Y(n_3217)
);

AO32x2_ASAP7_75t_L g3218 ( 
.A1(n_3067),
.A2(n_184),
.A3(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_3002),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_3026),
.A2(n_188),
.B(n_190),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_3058),
.A2(n_192),
.B(n_193),
.Y(n_3221)
);

OR2x6_ASAP7_75t_L g3222 ( 
.A(n_3029),
.B(n_337),
.Y(n_3222)
);

OAI21x1_ASAP7_75t_L g3223 ( 
.A1(n_2977),
.A2(n_439),
.B(n_438),
.Y(n_3223)
);

OAI21x1_ASAP7_75t_L g3224 ( 
.A1(n_2981),
.A2(n_437),
.B(n_428),
.Y(n_3224)
);

AND2x6_ASAP7_75t_L g3225 ( 
.A(n_3102),
.B(n_193),
.Y(n_3225)
);

INVx5_ASAP7_75t_L g3226 ( 
.A(n_3035),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_3009),
.B(n_195),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3050),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_3058),
.A2(n_195),
.B(n_196),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3039),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_3230)
);

AOI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_2947),
.A2(n_199),
.B(n_200),
.Y(n_3231)
);

INVx4_ASAP7_75t_L g3232 ( 
.A(n_3086),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3023),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3010),
.B(n_201),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_SL g3235 ( 
.A1(n_3085),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_3235)
);

AO31x2_ASAP7_75t_L g3236 ( 
.A1(n_3093),
.A2(n_3078),
.A3(n_3040),
.B(n_3069),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3020),
.Y(n_3237)
);

AO31x2_ASAP7_75t_L g3238 ( 
.A1(n_3065),
.A2(n_207),
.A3(n_211),
.B(n_212),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3045),
.A2(n_3108),
.B(n_3073),
.Y(n_3239)
);

OAI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_3039),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3045),
.A2(n_216),
.B(n_217),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_2951),
.A2(n_217),
.B(n_218),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3013),
.B(n_220),
.Y(n_3243)
);

NAND3xp33_ASAP7_75t_L g3244 ( 
.A(n_3074),
.B(n_221),
.C(n_222),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_2984),
.A2(n_222),
.B(n_223),
.Y(n_3245)
);

AO21x2_ASAP7_75t_L g3246 ( 
.A1(n_2995),
.A2(n_224),
.B(n_225),
.Y(n_3246)
);

A2O1A1Ixp33_ASAP7_75t_L g3247 ( 
.A1(n_2984),
.A2(n_224),
.B(n_225),
.C(n_226),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2990),
.B(n_229),
.Y(n_3248)
);

BUFx6f_ASAP7_75t_L g3249 ( 
.A(n_2958),
.Y(n_3249)
);

AOI221x1_ASAP7_75t_L g3250 ( 
.A1(n_3097),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.C(n_234),
.Y(n_3250)
);

HB1xp67_ASAP7_75t_L g3251 ( 
.A(n_3024),
.Y(n_3251)
);

OAI21x1_ASAP7_75t_SL g3252 ( 
.A1(n_3120),
.A2(n_3007),
.B(n_3024),
.Y(n_3252)
);

OAI21x1_ASAP7_75t_L g3253 ( 
.A1(n_3151),
.A2(n_2964),
.B(n_2994),
.Y(n_3253)
);

OA21x2_ASAP7_75t_L g3254 ( 
.A1(n_3140),
.A2(n_3090),
.B(n_3113),
.Y(n_3254)
);

OAI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_3131),
.A2(n_3087),
.B1(n_3091),
.B2(n_2991),
.Y(n_3255)
);

AO21x2_ASAP7_75t_L g3256 ( 
.A1(n_3176),
.A2(n_3021),
.B(n_2994),
.Y(n_3256)
);

AOI21x1_ASAP7_75t_SL g3257 ( 
.A1(n_3158),
.A2(n_3160),
.B(n_3152),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_3129),
.B(n_3243),
.Y(n_3258)
);

INVx5_ASAP7_75t_L g3259 ( 
.A(n_3222),
.Y(n_3259)
);

AOI21xp33_ASAP7_75t_SL g3260 ( 
.A1(n_3177),
.A2(n_3070),
.B(n_3079),
.Y(n_3260)
);

OAI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3231),
.A2(n_3087),
.B(n_3080),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3233),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_3119),
.B(n_2960),
.Y(n_3263)
);

INVx6_ASAP7_75t_L g3264 ( 
.A(n_3226),
.Y(n_3264)
);

BUFx3_ASAP7_75t_L g3265 ( 
.A(n_3166),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_3210),
.Y(n_3266)
);

OAI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_3136),
.A2(n_3067),
.B1(n_3116),
.B2(n_3054),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3128),
.A2(n_3156),
.B1(n_3123),
.B2(n_3192),
.Y(n_3268)
);

AOI21x1_ASAP7_75t_L g3269 ( 
.A1(n_3209),
.A2(n_3103),
.B(n_3034),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_L g3270 ( 
.A(n_3248),
.B(n_3134),
.Y(n_3270)
);

AO21x1_ASAP7_75t_L g3271 ( 
.A1(n_3221),
.A2(n_3067),
.B(n_3034),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_L g3272 ( 
.A1(n_3125),
.A2(n_3104),
.B1(n_3082),
.B2(n_2978),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3214),
.A2(n_3102),
.B1(n_3057),
.B2(n_3004),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_3251),
.Y(n_3274)
);

AOI22xp5_ASAP7_75t_L g3275 ( 
.A1(n_3196),
.A2(n_2968),
.B1(n_3005),
.B2(n_3072),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3121),
.A2(n_3044),
.B1(n_2968),
.B2(n_3113),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_3124),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3132),
.Y(n_3278)
);

OAI21x1_ASAP7_75t_L g3279 ( 
.A1(n_3239),
.A2(n_2959),
.B(n_3044),
.Y(n_3279)
);

OAI22xp5_ASAP7_75t_L g3280 ( 
.A1(n_3247),
.A2(n_2980),
.B1(n_3027),
.B2(n_3031),
.Y(n_3280)
);

OAI21x1_ASAP7_75t_L g3281 ( 
.A1(n_3130),
.A2(n_3011),
.B(n_3014),
.Y(n_3281)
);

AOI221xp5_ASAP7_75t_L g3282 ( 
.A1(n_3150),
.A2(n_3081),
.B1(n_3027),
.B2(n_2980),
.C(n_3033),
.Y(n_3282)
);

BUFx3_ASAP7_75t_L g3283 ( 
.A(n_3165),
.Y(n_3283)
);

OAI21x1_ASAP7_75t_L g3284 ( 
.A1(n_3155),
.A2(n_3101),
.B(n_3112),
.Y(n_3284)
);

AO32x2_ASAP7_75t_L g3285 ( 
.A1(n_3199),
.A2(n_2950),
.A3(n_2960),
.B1(n_3048),
.B2(n_3028),
.Y(n_3285)
);

INVx4_ASAP7_75t_L g3286 ( 
.A(n_3190),
.Y(n_3286)
);

BUFx6f_ASAP7_75t_L g3287 ( 
.A(n_3204),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3184),
.B(n_2950),
.Y(n_3288)
);

INVx8_ASAP7_75t_L g3289 ( 
.A(n_3222),
.Y(n_3289)
);

OA21x2_ASAP7_75t_L g3290 ( 
.A1(n_3202),
.A2(n_3114),
.B(n_3056),
.Y(n_3290)
);

OAI21x1_ASAP7_75t_L g3291 ( 
.A1(n_3153),
.A2(n_3015),
.B(n_3109),
.Y(n_3291)
);

OA21x2_ASAP7_75t_L g3292 ( 
.A1(n_3203),
.A2(n_3022),
.B(n_3066),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3237),
.B(n_3086),
.Y(n_3293)
);

OA21x2_ASAP7_75t_L g3294 ( 
.A1(n_3170),
.A2(n_3066),
.B(n_3061),
.Y(n_3294)
);

AOI22xp33_ASAP7_75t_L g3295 ( 
.A1(n_3179),
.A2(n_2965),
.B1(n_3028),
.B2(n_3081),
.Y(n_3295)
);

OAI21x1_ASAP7_75t_L g3296 ( 
.A1(n_3223),
.A2(n_2966),
.B(n_3064),
.Y(n_3296)
);

HB1xp67_ASAP7_75t_L g3297 ( 
.A(n_3157),
.Y(n_3297)
);

INVx1_ASAP7_75t_SL g3298 ( 
.A(n_3149),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3169),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3171),
.Y(n_3300)
);

AO21x2_ASAP7_75t_L g3301 ( 
.A1(n_3118),
.A2(n_3095),
.B(n_2965),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3163),
.A2(n_3037),
.B1(n_3030),
.B2(n_3060),
.Y(n_3302)
);

OAI21x1_ASAP7_75t_L g3303 ( 
.A1(n_3224),
.A2(n_3051),
.B(n_3049),
.Y(n_3303)
);

AND2x4_ASAP7_75t_L g3304 ( 
.A(n_3119),
.B(n_3048),
.Y(n_3304)
);

OAI21x1_ASAP7_75t_L g3305 ( 
.A1(n_3138),
.A2(n_3048),
.B(n_234),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3186),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3188),
.Y(n_3307)
);

OAI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3229),
.A2(n_233),
.B(n_236),
.Y(n_3308)
);

AO21x2_ASAP7_75t_L g3309 ( 
.A1(n_3182),
.A2(n_237),
.B(n_238),
.Y(n_3309)
);

OAI21x1_ASAP7_75t_L g3310 ( 
.A1(n_3162),
.A2(n_3147),
.B(n_3201),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_L g3311 ( 
.A1(n_3213),
.A2(n_238),
.B(n_239),
.Y(n_3311)
);

OR2x6_ASAP7_75t_SL g3312 ( 
.A(n_3137),
.B(n_240),
.Y(n_3312)
);

OAI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3241),
.A2(n_3161),
.B(n_3217),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3206),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_3167),
.Y(n_3315)
);

BUFx2_ASAP7_75t_L g3316 ( 
.A(n_3208),
.Y(n_3316)
);

NAND2x1p5_ASAP7_75t_L g3317 ( 
.A(n_3190),
.B(n_3232),
.Y(n_3317)
);

OA21x2_ASAP7_75t_L g3318 ( 
.A1(n_3141),
.A2(n_240),
.B(n_241),
.Y(n_3318)
);

HB1xp67_ASAP7_75t_L g3319 ( 
.A(n_3173),
.Y(n_3319)
);

AO21x2_ASAP7_75t_L g3320 ( 
.A1(n_3220),
.A2(n_242),
.B(n_243),
.Y(n_3320)
);

OAI21x1_ASAP7_75t_L g3321 ( 
.A1(n_3242),
.A2(n_242),
.B(n_244),
.Y(n_3321)
);

OR2x2_ASAP7_75t_L g3322 ( 
.A(n_3219),
.B(n_245),
.Y(n_3322)
);

AOI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_3244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_3323)
);

OAI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3197),
.A2(n_248),
.B(n_249),
.Y(n_3324)
);

OA21x2_ASAP7_75t_L g3325 ( 
.A1(n_3195),
.A2(n_250),
.B(n_251),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3228),
.Y(n_3326)
);

INVx3_ASAP7_75t_L g3327 ( 
.A(n_3249),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3133),
.Y(n_3328)
);

BUFx12f_ASAP7_75t_L g3329 ( 
.A(n_3144),
.Y(n_3329)
);

AOI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_3200),
.A2(n_348),
.B(n_408),
.Y(n_3330)
);

INVx4_ASAP7_75t_L g3331 ( 
.A(n_3232),
.Y(n_3331)
);

OAI21x1_ASAP7_75t_L g3332 ( 
.A1(n_3178),
.A2(n_251),
.B(n_252),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3133),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_SL g3334 ( 
.A1(n_3175),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_3334)
);

AND2x4_ASAP7_75t_L g3335 ( 
.A(n_3180),
.B(n_253),
.Y(n_3335)
);

OAI21x1_ASAP7_75t_SL g3336 ( 
.A1(n_3212),
.A2(n_255),
.B(n_256),
.Y(n_3336)
);

BUFx3_ASAP7_75t_L g3337 ( 
.A(n_3249),
.Y(n_3337)
);

OA21x2_ASAP7_75t_L g3338 ( 
.A1(n_3245),
.A2(n_256),
.B(n_257),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3139),
.B(n_260),
.Y(n_3339)
);

OR2x6_ASAP7_75t_L g3340 ( 
.A(n_3122),
.B(n_261),
.Y(n_3340)
);

OR2x6_ASAP7_75t_L g3341 ( 
.A(n_3122),
.B(n_261),
.Y(n_3341)
);

OAI21x1_ASAP7_75t_L g3342 ( 
.A1(n_3180),
.A2(n_262),
.B(n_263),
.Y(n_3342)
);

O2A1O1Ixp33_ASAP7_75t_SL g3343 ( 
.A1(n_3146),
.A2(n_3135),
.B(n_3159),
.C(n_3230),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3215),
.B(n_264),
.Y(n_3344)
);

BUFx2_ASAP7_75t_L g3345 ( 
.A(n_3208),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3198),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_3346)
);

OAI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_3148),
.A2(n_3168),
.B(n_3183),
.Y(n_3347)
);

HB1xp67_ASAP7_75t_L g3348 ( 
.A(n_3164),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3234),
.B(n_266),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3216),
.B(n_267),
.Y(n_3350)
);

OA21x2_ASAP7_75t_L g3351 ( 
.A1(n_3250),
.A2(n_267),
.B(n_268),
.Y(n_3351)
);

CKINVDCx5p33_ASAP7_75t_R g3352 ( 
.A(n_3142),
.Y(n_3352)
);

OAI21x1_ASAP7_75t_L g3353 ( 
.A1(n_3207),
.A2(n_268),
.B(n_269),
.Y(n_3353)
);

AO21x1_ASAP7_75t_L g3354 ( 
.A1(n_3218),
.A2(n_269),
.B(n_272),
.Y(n_3354)
);

O2A1O1Ixp33_ASAP7_75t_SL g3355 ( 
.A1(n_3240),
.A2(n_273),
.B(n_274),
.C(n_277),
.Y(n_3355)
);

AOI221xp5_ASAP7_75t_L g3356 ( 
.A1(n_3172),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.C(n_283),
.Y(n_3356)
);

OAI21x1_ASAP7_75t_L g3357 ( 
.A1(n_3126),
.A2(n_285),
.B(n_286),
.Y(n_3357)
);

HB1xp67_ASAP7_75t_L g3358 ( 
.A(n_3164),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3133),
.Y(n_3359)
);

AO31x2_ASAP7_75t_L g3360 ( 
.A1(n_3154),
.A2(n_285),
.A3(n_286),
.B(n_338),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3164),
.Y(n_3361)
);

AOI211xp5_ASAP7_75t_SL g3362 ( 
.A1(n_3343),
.A2(n_3174),
.B(n_3189),
.C(n_3127),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_3268),
.A2(n_3235),
.B1(n_3225),
.B2(n_3205),
.Y(n_3363)
);

A2O1A1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_3313),
.A2(n_3145),
.B(n_3227),
.C(n_3185),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3297),
.Y(n_3365)
);

HB1xp67_ASAP7_75t_L g3366 ( 
.A(n_3266),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3288),
.B(n_3143),
.Y(n_3367)
);

BUFx8_ASAP7_75t_L g3368 ( 
.A(n_3349),
.Y(n_3368)
);

A2O1A1Ixp33_ASAP7_75t_L g3369 ( 
.A1(n_3347),
.A2(n_3193),
.B(n_3218),
.C(n_3191),
.Y(n_3369)
);

INVx3_ASAP7_75t_L g3370 ( 
.A(n_3264),
.Y(n_3370)
);

AO21x2_ASAP7_75t_L g3371 ( 
.A1(n_3266),
.A2(n_3358),
.B(n_3348),
.Y(n_3371)
);

NOR2x1_ASAP7_75t_SL g3372 ( 
.A(n_3256),
.B(n_3246),
.Y(n_3372)
);

INVx3_ASAP7_75t_L g3373 ( 
.A(n_3264),
.Y(n_3373)
);

OAI21x1_ASAP7_75t_L g3374 ( 
.A1(n_3279),
.A2(n_3218),
.B(n_3181),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3297),
.B(n_3143),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3268),
.A2(n_3191),
.B1(n_3194),
.B2(n_3226),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_3324),
.A2(n_3225),
.B1(n_3191),
.B2(n_3143),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3293),
.B(n_3181),
.Y(n_3378)
);

INVx3_ASAP7_75t_L g3379 ( 
.A(n_3264),
.Y(n_3379)
);

AOI21x1_ASAP7_75t_L g3380 ( 
.A1(n_3354),
.A2(n_3344),
.B(n_3316),
.Y(n_3380)
);

AO31x2_ASAP7_75t_L g3381 ( 
.A1(n_3271),
.A2(n_3211),
.A3(n_3181),
.B(n_3187),
.Y(n_3381)
);

AO31x2_ASAP7_75t_L g3382 ( 
.A1(n_3328),
.A2(n_3211),
.A3(n_3187),
.B(n_3238),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_3258),
.B(n_3225),
.Y(n_3383)
);

A2O1A1Ixp33_ASAP7_75t_L g3384 ( 
.A1(n_3308),
.A2(n_3225),
.B(n_3211),
.C(n_3187),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3277),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3277),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3299),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3299),
.Y(n_3388)
);

INVx3_ASAP7_75t_L g3389 ( 
.A(n_3286),
.Y(n_3389)
);

OAI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_3330),
.A2(n_3236),
.B(n_343),
.Y(n_3390)
);

OAI21x1_ASAP7_75t_SL g3391 ( 
.A1(n_3252),
.A2(n_345),
.B(n_347),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_3274),
.B(n_350),
.Y(n_3392)
);

AO31x2_ASAP7_75t_L g3393 ( 
.A1(n_3333),
.A2(n_351),
.A3(n_354),
.B(n_355),
.Y(n_3393)
);

CKINVDCx5p33_ASAP7_75t_R g3394 ( 
.A(n_3352),
.Y(n_3394)
);

HB1xp67_ASAP7_75t_L g3395 ( 
.A(n_3256),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3262),
.B(n_360),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_3343),
.A2(n_361),
.B(n_363),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3262),
.B(n_364),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3278),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3306),
.B(n_367),
.Y(n_3400)
);

BUFx6f_ASAP7_75t_L g3401 ( 
.A(n_3287),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3259),
.A2(n_373),
.B(n_375),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3307),
.B(n_378),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3314),
.B(n_380),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_3356),
.A2(n_381),
.B(n_383),
.C(n_384),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_3352),
.Y(n_3406)
);

OA21x2_ASAP7_75t_L g3407 ( 
.A1(n_3361),
.A2(n_389),
.B(n_390),
.Y(n_3407)
);

OA21x2_ASAP7_75t_L g3408 ( 
.A1(n_3359),
.A2(n_393),
.B(n_394),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3300),
.B(n_397),
.Y(n_3409)
);

CKINVDCx5p33_ASAP7_75t_R g3410 ( 
.A(n_3329),
.Y(n_3410)
);

HB1xp67_ASAP7_75t_L g3411 ( 
.A(n_3319),
.Y(n_3411)
);

AO31x2_ASAP7_75t_L g3412 ( 
.A1(n_3276),
.A2(n_404),
.A3(n_406),
.B(n_407),
.Y(n_3412)
);

BUFx5_ASAP7_75t_L g3413 ( 
.A(n_3304),
.Y(n_3413)
);

INVx4_ASAP7_75t_L g3414 ( 
.A(n_3289),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3326),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_SL g3416 ( 
.A(n_3259),
.B(n_3267),
.Y(n_3416)
);

AND2x2_ASAP7_75t_L g3417 ( 
.A(n_3283),
.B(n_3345),
.Y(n_3417)
);

OA21x2_ASAP7_75t_L g3418 ( 
.A1(n_3263),
.A2(n_3358),
.B(n_3253),
.Y(n_3418)
);

AO31x2_ASAP7_75t_L g3419 ( 
.A1(n_3331),
.A2(n_3280),
.A3(n_3255),
.B(n_3270),
.Y(n_3419)
);

AND2x4_ASAP7_75t_L g3420 ( 
.A(n_3265),
.B(n_3304),
.Y(n_3420)
);

AOI211x1_ASAP7_75t_L g3421 ( 
.A1(n_3267),
.A2(n_3261),
.B(n_3346),
.C(n_3339),
.Y(n_3421)
);

OAI21x1_ASAP7_75t_L g3422 ( 
.A1(n_3253),
.A2(n_3296),
.B(n_3254),
.Y(n_3422)
);

OAI21xp5_ASAP7_75t_L g3423 ( 
.A1(n_3338),
.A2(n_3318),
.B(n_3323),
.Y(n_3423)
);

OAI21x1_ASAP7_75t_L g3424 ( 
.A1(n_3254),
.A2(n_3281),
.B(n_3269),
.Y(n_3424)
);

AOI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_3259),
.A2(n_3351),
.B(n_3318),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3322),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3265),
.B(n_3298),
.Y(n_3427)
);

AO21x2_ASAP7_75t_L g3428 ( 
.A1(n_3301),
.A2(n_3320),
.B(n_3357),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3254),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3259),
.A2(n_3351),
.B(n_3318),
.Y(n_3430)
);

CKINVDCx11_ASAP7_75t_R g3431 ( 
.A(n_3312),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3270),
.B(n_3295),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3295),
.B(n_3301),
.Y(n_3433)
);

AO31x2_ASAP7_75t_L g3434 ( 
.A1(n_3350),
.A2(n_3285),
.A3(n_3338),
.B(n_3320),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3287),
.Y(n_3435)
);

AOI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3325),
.A2(n_3351),
.B1(n_3338),
.B2(n_3289),
.Y(n_3436)
);

CKINVDCx6p67_ASAP7_75t_R g3437 ( 
.A(n_3315),
.Y(n_3437)
);

OAI21x1_ASAP7_75t_L g3438 ( 
.A1(n_3317),
.A2(n_3284),
.B(n_3310),
.Y(n_3438)
);

AND2x4_ASAP7_75t_L g3439 ( 
.A(n_3337),
.B(n_3327),
.Y(n_3439)
);

AO21x2_ASAP7_75t_L g3440 ( 
.A1(n_3357),
.A2(n_3336),
.B(n_3260),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3302),
.B(n_3292),
.Y(n_3441)
);

AOI22xp33_ASAP7_75t_L g3442 ( 
.A1(n_3416),
.A2(n_3325),
.B1(n_3289),
.B2(n_3309),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3431),
.A2(n_3325),
.B1(n_3323),
.B2(n_3309),
.Y(n_3443)
);

INVx2_ASAP7_75t_SL g3444 ( 
.A(n_3427),
.Y(n_3444)
);

INVx4_ASAP7_75t_SL g3445 ( 
.A(n_3412),
.Y(n_3445)
);

CKINVDCx5p33_ASAP7_75t_R g3446 ( 
.A(n_3394),
.Y(n_3446)
);

BUFx2_ASAP7_75t_L g3447 ( 
.A(n_3414),
.Y(n_3447)
);

OAI21xp5_ASAP7_75t_SL g3448 ( 
.A1(n_3362),
.A2(n_3272),
.B(n_3334),
.Y(n_3448)
);

INVx4_ASAP7_75t_L g3449 ( 
.A(n_3437),
.Y(n_3449)
);

CKINVDCx11_ASAP7_75t_R g3450 ( 
.A(n_3406),
.Y(n_3450)
);

AOI22xp33_ASAP7_75t_L g3451 ( 
.A1(n_3432),
.A2(n_3272),
.B1(n_3341),
.B2(n_3340),
.Y(n_3451)
);

OAI21xp5_ASAP7_75t_SL g3452 ( 
.A1(n_3362),
.A2(n_3273),
.B(n_3282),
.Y(n_3452)
);

INVx4_ASAP7_75t_L g3453 ( 
.A(n_3410),
.Y(n_3453)
);

AOI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3376),
.A2(n_3355),
.B1(n_3341),
.B2(n_3340),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_3432),
.A2(n_3340),
.B1(n_3321),
.B2(n_3332),
.Y(n_3455)
);

OAI21xp5_ASAP7_75t_SL g3456 ( 
.A1(n_3363),
.A2(n_3364),
.B(n_3397),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3423),
.A2(n_3335),
.B1(n_3275),
.B2(n_3292),
.Y(n_3457)
);

AOI22xp33_ASAP7_75t_SL g3458 ( 
.A1(n_3376),
.A2(n_3335),
.B1(n_3311),
.B2(n_3342),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_SL g3459 ( 
.A1(n_3423),
.A2(n_3335),
.B1(n_3353),
.B2(n_3257),
.Y(n_3459)
);

NAND2xp33_ASAP7_75t_L g3460 ( 
.A(n_3369),
.B(n_3355),
.Y(n_3460)
);

INVx3_ASAP7_75t_L g3461 ( 
.A(n_3414),
.Y(n_3461)
);

OAI21xp5_ASAP7_75t_SL g3462 ( 
.A1(n_3363),
.A2(n_3360),
.B(n_3305),
.Y(n_3462)
);

INVx4_ASAP7_75t_L g3463 ( 
.A(n_3401),
.Y(n_3463)
);

AOI222xp33_ASAP7_75t_L g3464 ( 
.A1(n_3377),
.A2(n_3360),
.B1(n_3303),
.B2(n_3291),
.C1(n_3294),
.C2(n_3285),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_SL g3465 ( 
.A1(n_3425),
.A2(n_3294),
.B1(n_3292),
.B2(n_3290),
.Y(n_3465)
);

BUFx2_ASAP7_75t_L g3466 ( 
.A(n_3370),
.Y(n_3466)
);

CKINVDCx8_ASAP7_75t_R g3467 ( 
.A(n_3439),
.Y(n_3467)
);

AOI22xp33_ASAP7_75t_L g3468 ( 
.A1(n_3390),
.A2(n_3285),
.B1(n_3360),
.B2(n_3383),
.Y(n_3468)
);

OAI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_3421),
.A2(n_3384),
.B1(n_3436),
.B2(n_3430),
.Y(n_3469)
);

AOI22xp33_ASAP7_75t_SL g3470 ( 
.A1(n_3425),
.A2(n_3430),
.B1(n_3372),
.B2(n_3428),
.Y(n_3470)
);

INVxp67_ASAP7_75t_L g3471 ( 
.A(n_3440),
.Y(n_3471)
);

HB1xp67_ASAP7_75t_L g3472 ( 
.A(n_3371),
.Y(n_3472)
);

BUFx6f_ASAP7_75t_L g3473 ( 
.A(n_3408),
.Y(n_3473)
);

CKINVDCx11_ASAP7_75t_R g3474 ( 
.A(n_3435),
.Y(n_3474)
);

BUFx12f_ASAP7_75t_L g3475 ( 
.A(n_3368),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3411),
.Y(n_3476)
);

OAI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3405),
.A2(n_3380),
.B1(n_3390),
.B2(n_3433),
.Y(n_3477)
);

INVx2_ASAP7_75t_SL g3478 ( 
.A(n_3417),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3411),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_3368),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_SL g3481 ( 
.A1(n_3428),
.A2(n_3440),
.B1(n_3374),
.B2(n_3391),
.Y(n_3481)
);

OAI21xp5_ASAP7_75t_SL g3482 ( 
.A1(n_3402),
.A2(n_3441),
.B(n_3378),
.Y(n_3482)
);

AOI222xp33_ASAP7_75t_L g3483 ( 
.A1(n_3426),
.A2(n_3441),
.B1(n_3367),
.B2(n_3375),
.C1(n_3409),
.C2(n_3400),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_L g3484 ( 
.A(n_3370),
.B(n_3373),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3373),
.B(n_3379),
.Y(n_3485)
);

CKINVDCx5p33_ASAP7_75t_R g3486 ( 
.A(n_3389),
.Y(n_3486)
);

OAI21xp5_ASAP7_75t_SL g3487 ( 
.A1(n_3375),
.A2(n_3420),
.B(n_3389),
.Y(n_3487)
);

OAI22xp5_ASAP7_75t_SL g3488 ( 
.A1(n_3407),
.A2(n_3408),
.B1(n_3439),
.B2(n_3395),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3392),
.B(n_3400),
.Y(n_3489)
);

OAI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3409),
.A2(n_3403),
.B1(n_3404),
.B2(n_3398),
.Y(n_3490)
);

OAI222xp33_ASAP7_75t_L g3491 ( 
.A1(n_3403),
.A2(n_3404),
.B1(n_3396),
.B2(n_3398),
.C1(n_3395),
.C2(n_3365),
.Y(n_3491)
);

AOI211xp5_ASAP7_75t_SL g3492 ( 
.A1(n_3366),
.A2(n_3429),
.B(n_3419),
.C(n_3381),
.Y(n_3492)
);

CKINVDCx20_ASAP7_75t_R g3493 ( 
.A(n_3415),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3434),
.B(n_3419),
.Y(n_3494)
);

OAI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_3422),
.A2(n_3424),
.B(n_3438),
.Y(n_3495)
);

CKINVDCx6p67_ASAP7_75t_R g3496 ( 
.A(n_3366),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_L g3497 ( 
.A1(n_3385),
.A2(n_3386),
.B1(n_3387),
.B2(n_3388),
.Y(n_3497)
);

OAI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_3418),
.A2(n_3419),
.B1(n_3381),
.B2(n_3412),
.Y(n_3498)
);

OAI22xp33_ASAP7_75t_L g3499 ( 
.A1(n_3412),
.A2(n_3381),
.B1(n_3418),
.B2(n_3434),
.Y(n_3499)
);

INVxp67_ASAP7_75t_SL g3500 ( 
.A(n_3413),
.Y(n_3500)
);

OAI22xp33_ASAP7_75t_L g3501 ( 
.A1(n_3382),
.A2(n_3362),
.B1(n_3131),
.B2(n_3376),
.Y(n_3501)
);

OAI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3393),
.A2(n_3377),
.B1(n_3421),
.B2(n_3268),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3393),
.B(n_3378),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3416),
.A2(n_3431),
.B1(n_3423),
.B2(n_3432),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3432),
.B(n_3421),
.Y(n_3505)
);

INVxp67_ASAP7_75t_SL g3506 ( 
.A(n_3395),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3401),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3377),
.A2(n_3421),
.B1(n_3268),
.B2(n_3369),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3431),
.A2(n_3268),
.B1(n_3324),
.B2(n_3432),
.Y(n_3509)
);

OAI21xp5_ASAP7_75t_SL g3510 ( 
.A1(n_3362),
.A2(n_3268),
.B(n_3313),
.Y(n_3510)
);

CKINVDCx5p33_ASAP7_75t_R g3511 ( 
.A(n_3394),
.Y(n_3511)
);

OAI22xp5_ASAP7_75t_L g3512 ( 
.A1(n_3377),
.A2(n_3421),
.B1(n_3268),
.B2(n_3369),
.Y(n_3512)
);

OAI22xp5_ASAP7_75t_L g3513 ( 
.A1(n_3377),
.A2(n_3421),
.B1(n_3268),
.B2(n_3369),
.Y(n_3513)
);

CKINVDCx5p33_ASAP7_75t_R g3514 ( 
.A(n_3394),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3399),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3414),
.B(n_3437),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3377),
.A2(n_3421),
.B1(n_3268),
.B2(n_3369),
.Y(n_3517)
);

AOI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_3376),
.A2(n_3416),
.B1(n_3268),
.B2(n_3397),
.Y(n_3518)
);

AOI22xp33_ASAP7_75t_L g3519 ( 
.A1(n_3431),
.A2(n_3268),
.B1(n_3324),
.B2(n_3432),
.Y(n_3519)
);

AO21x2_ASAP7_75t_L g3520 ( 
.A1(n_3499),
.A2(n_3501),
.B(n_3472),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3466),
.B(n_3447),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3472),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_SL g3523 ( 
.A1(n_3508),
.A2(n_3513),
.B1(n_3512),
.B2(n_3517),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3503),
.B(n_3496),
.Y(n_3524)
);

OR2x2_ASAP7_75t_L g3525 ( 
.A(n_3476),
.B(n_3479),
.Y(n_3525)
);

AO21x2_ASAP7_75t_L g3526 ( 
.A1(n_3499),
.A2(n_3501),
.B(n_3506),
.Y(n_3526)
);

HB1xp67_ASAP7_75t_L g3527 ( 
.A(n_3445),
.Y(n_3527)
);

BUFx3_ASAP7_75t_L g3528 ( 
.A(n_3475),
.Y(n_3528)
);

AOI21x1_ASAP7_75t_L g3529 ( 
.A1(n_3469),
.A2(n_3505),
.B(n_3494),
.Y(n_3529)
);

INVx3_ASAP7_75t_L g3530 ( 
.A(n_3467),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3461),
.B(n_3484),
.Y(n_3531)
);

AO21x2_ASAP7_75t_L g3532 ( 
.A1(n_3506),
.A2(n_3498),
.B(n_3518),
.Y(n_3532)
);

BUFx2_ASAP7_75t_L g3533 ( 
.A(n_3449),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3456),
.A2(n_3510),
.B(n_3477),
.Y(n_3534)
);

OR2x6_ASAP7_75t_L g3535 ( 
.A(n_3462),
.B(n_3473),
.Y(n_3535)
);

BUFx3_ASAP7_75t_L g3536 ( 
.A(n_3480),
.Y(n_3536)
);

AND2x4_ASAP7_75t_L g3537 ( 
.A(n_3445),
.B(n_3500),
.Y(n_3537)
);

NAND3xp33_ASAP7_75t_L g3538 ( 
.A(n_3509),
.B(n_3519),
.C(n_3504),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3461),
.B(n_3485),
.Y(n_3539)
);

HB1xp67_ASAP7_75t_L g3540 ( 
.A(n_3445),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3515),
.B(n_3497),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3502),
.B(n_3509),
.Y(n_3542)
);

HB1xp67_ASAP7_75t_L g3543 ( 
.A(n_3444),
.Y(n_3543)
);

AO21x2_ASAP7_75t_L g3544 ( 
.A1(n_3471),
.A2(n_3495),
.B(n_3482),
.Y(n_3544)
);

BUFx2_ASAP7_75t_L g3545 ( 
.A(n_3449),
.Y(n_3545)
);

OR2x6_ASAP7_75t_L g3546 ( 
.A(n_3452),
.B(n_3448),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3519),
.B(n_3459),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3463),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3493),
.Y(n_3549)
);

INVx5_ASAP7_75t_SL g3550 ( 
.A(n_3507),
.Y(n_3550)
);

INVx3_ASAP7_75t_L g3551 ( 
.A(n_3453),
.Y(n_3551)
);

BUFx2_ASAP7_75t_L g3552 ( 
.A(n_3486),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3478),
.B(n_3459),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3488),
.Y(n_3554)
);

INVx6_ASAP7_75t_L g3555 ( 
.A(n_3453),
.Y(n_3555)
);

BUFx3_ASAP7_75t_L g3556 ( 
.A(n_3450),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3460),
.Y(n_3557)
);

AO21x2_ASAP7_75t_L g3558 ( 
.A1(n_3454),
.A2(n_3487),
.B(n_3470),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3474),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3458),
.B(n_3470),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3483),
.B(n_3490),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3481),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_3492),
.Y(n_3563)
);

BUFx2_ASAP7_75t_L g3564 ( 
.A(n_3516),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3451),
.B(n_3455),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3457),
.B(n_3481),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3489),
.Y(n_3567)
);

OR2x2_ASAP7_75t_L g3568 ( 
.A(n_3442),
.B(n_3468),
.Y(n_3568)
);

AO21x2_ASAP7_75t_L g3569 ( 
.A1(n_3491),
.A2(n_3465),
.B(n_3464),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3446),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3443),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3443),
.Y(n_3572)
);

OR2x6_ASAP7_75t_L g3573 ( 
.A(n_3465),
.B(n_3511),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3514),
.Y(n_3574)
);

AND2x4_ASAP7_75t_L g3575 ( 
.A(n_3445),
.B(n_3500),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3466),
.B(n_3447),
.Y(n_3576)
);

HB1xp67_ASAP7_75t_L g3577 ( 
.A(n_3445),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3472),
.Y(n_3578)
);

AOI21x1_ASAP7_75t_L g3579 ( 
.A1(n_3472),
.A2(n_3469),
.B(n_3508),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3472),
.Y(n_3580)
);

BUFx3_ASAP7_75t_L g3581 ( 
.A(n_3475),
.Y(n_3581)
);

NAND2x1p5_ASAP7_75t_L g3582 ( 
.A(n_3473),
.B(n_3425),
.Y(n_3582)
);

AOI22xp33_ASAP7_75t_L g3583 ( 
.A1(n_3508),
.A2(n_3512),
.B1(n_3517),
.B2(n_3513),
.Y(n_3583)
);

OR2x6_ASAP7_75t_L g3584 ( 
.A(n_3456),
.B(n_3397),
.Y(n_3584)
);

AO21x2_ASAP7_75t_L g3585 ( 
.A1(n_3499),
.A2(n_3501),
.B(n_3472),
.Y(n_3585)
);

OAI21x1_ASAP7_75t_L g3586 ( 
.A1(n_3498),
.A2(n_3469),
.B(n_3416),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3466),
.B(n_3447),
.Y(n_3587)
);

INVxp67_ASAP7_75t_L g3588 ( 
.A(n_3460),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3472),
.Y(n_3589)
);

INVx5_ASAP7_75t_SL g3590 ( 
.A(n_3584),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3582),
.Y(n_3591)
);

HB1xp67_ASAP7_75t_L g3592 ( 
.A(n_3582),
.Y(n_3592)
);

NAND2x1p5_ASAP7_75t_SL g3593 ( 
.A(n_3560),
.B(n_3566),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3582),
.Y(n_3594)
);

NOR2xp67_ASAP7_75t_L g3595 ( 
.A(n_3530),
.B(n_3588),
.Y(n_3595)
);

AND2x4_ASAP7_75t_L g3596 ( 
.A(n_3526),
.B(n_3520),
.Y(n_3596)
);

OR2x2_ASAP7_75t_L g3597 ( 
.A(n_3525),
.B(n_3541),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3521),
.B(n_3576),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3521),
.B(n_3576),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3587),
.B(n_3530),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3526),
.Y(n_3601)
);

OR2x2_ASAP7_75t_L g3602 ( 
.A(n_3525),
.B(n_3541),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3587),
.B(n_3530),
.Y(n_3603)
);

OR2x2_ASAP7_75t_L g3604 ( 
.A(n_3567),
.B(n_3526),
.Y(n_3604)
);

BUFx3_ASAP7_75t_L g3605 ( 
.A(n_3556),
.Y(n_3605)
);

BUFx2_ASAP7_75t_L g3606 ( 
.A(n_3520),
.Y(n_3606)
);

INVxp67_ASAP7_75t_SL g3607 ( 
.A(n_3556),
.Y(n_3607)
);

BUFx3_ASAP7_75t_L g3608 ( 
.A(n_3556),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3522),
.Y(n_3609)
);

NAND2x1_ASAP7_75t_L g3610 ( 
.A(n_3573),
.B(n_3584),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3530),
.B(n_3564),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_3520),
.B(n_3585),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3522),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3522),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3528),
.B(n_3581),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3585),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3564),
.B(n_3531),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_3528),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3531),
.B(n_3539),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3585),
.Y(n_3620)
);

HB1xp67_ASAP7_75t_L g3621 ( 
.A(n_3527),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3578),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3578),
.Y(n_3623)
);

BUFx2_ASAP7_75t_L g3624 ( 
.A(n_3533),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3524),
.B(n_3533),
.Y(n_3625)
);

AND2x4_ASAP7_75t_L g3626 ( 
.A(n_3537),
.B(n_3575),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3545),
.B(n_3550),
.Y(n_3627)
);

INVx3_ASAP7_75t_L g3628 ( 
.A(n_3569),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3578),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3523),
.B(n_3583),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3557),
.B(n_3554),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3580),
.Y(n_3632)
);

BUFx2_ASAP7_75t_L g3633 ( 
.A(n_3545),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3550),
.B(n_3553),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3569),
.Y(n_3635)
);

NAND2x1_ASAP7_75t_L g3636 ( 
.A(n_3573),
.B(n_3584),
.Y(n_3636)
);

INVx2_ASAP7_75t_SL g3637 ( 
.A(n_3537),
.Y(n_3637)
);

BUFx3_ASAP7_75t_L g3638 ( 
.A(n_3528),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3550),
.B(n_3553),
.Y(n_3639)
);

HB1xp67_ASAP7_75t_L g3640 ( 
.A(n_3540),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3569),
.Y(n_3641)
);

NOR2x1_ASAP7_75t_L g3642 ( 
.A(n_3573),
.B(n_3584),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3580),
.Y(n_3643)
);

INVx3_ASAP7_75t_L g3644 ( 
.A(n_3573),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3580),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3589),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3550),
.B(n_3552),
.Y(n_3647)
);

HB1xp67_ASAP7_75t_L g3648 ( 
.A(n_3577),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3550),
.B(n_3552),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3532),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3589),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3532),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3589),
.Y(n_3653)
);

NOR2x1_ASAP7_75t_L g3654 ( 
.A(n_3573),
.B(n_3584),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3549),
.B(n_3559),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3549),
.B(n_3559),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3549),
.B(n_3548),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3532),
.Y(n_3658)
);

AND2x4_ASAP7_75t_SL g3659 ( 
.A(n_3535),
.B(n_3543),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3560),
.Y(n_3660)
);

INVx3_ASAP7_75t_L g3661 ( 
.A(n_3536),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3537),
.Y(n_3662)
);

INVx3_ASAP7_75t_L g3663 ( 
.A(n_3536),
.Y(n_3663)
);

BUFx3_ASAP7_75t_L g3664 ( 
.A(n_3581),
.Y(n_3664)
);

NOR2xp33_ASAP7_75t_L g3665 ( 
.A(n_3581),
.B(n_3536),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_3548),
.B(n_3554),
.Y(n_3666)
);

INVxp67_ASAP7_75t_L g3667 ( 
.A(n_3557),
.Y(n_3667)
);

BUFx2_ASAP7_75t_L g3668 ( 
.A(n_3537),
.Y(n_3668)
);

BUFx6f_ASAP7_75t_L g3669 ( 
.A(n_3555),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3612),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3596),
.B(n_3558),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3606),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3596),
.B(n_3558),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3596),
.B(n_3558),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3606),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3612),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3612),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3612),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3596),
.B(n_3572),
.Y(n_3679)
);

INVxp67_ASAP7_75t_L g3680 ( 
.A(n_3611),
.Y(n_3680)
);

AND2x2_ASAP7_75t_SL g3681 ( 
.A(n_3635),
.B(n_3547),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3616),
.Y(n_3682)
);

AND2x2_ASAP7_75t_L g3683 ( 
.A(n_3628),
.B(n_3586),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3628),
.B(n_3586),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3616),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3628),
.B(n_3534),
.Y(n_3686)
);

BUFx2_ASAP7_75t_L g3687 ( 
.A(n_3616),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3628),
.B(n_3571),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3642),
.B(n_3535),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3620),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3620),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3642),
.B(n_3535),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3620),
.Y(n_3693)
);

BUFx3_ASAP7_75t_L g3694 ( 
.A(n_3601),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3654),
.B(n_3535),
.Y(n_3695)
);

OR2x2_ASAP7_75t_L g3696 ( 
.A(n_3601),
.B(n_3635),
.Y(n_3696)
);

INVxp67_ASAP7_75t_SL g3697 ( 
.A(n_3604),
.Y(n_3697)
);

HB1xp67_ASAP7_75t_L g3698 ( 
.A(n_3635),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3641),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3650),
.Y(n_3700)
);

HB1xp67_ASAP7_75t_L g3701 ( 
.A(n_3641),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3654),
.B(n_3535),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3641),
.B(n_3563),
.Y(n_3703)
);

BUFx3_ASAP7_75t_L g3704 ( 
.A(n_3650),
.Y(n_3704)
);

INVx3_ASAP7_75t_L g3705 ( 
.A(n_3650),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3600),
.B(n_3579),
.Y(n_3706)
);

INVxp67_ASAP7_75t_SL g3707 ( 
.A(n_3604),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3652),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3652),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_SL g3710 ( 
.A(n_3605),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3652),
.Y(n_3711)
);

OR2x2_ASAP7_75t_L g3712 ( 
.A(n_3593),
.B(n_3562),
.Y(n_3712)
);

HB1xp67_ASAP7_75t_L g3713 ( 
.A(n_3658),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3658),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3658),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3624),
.Y(n_3716)
);

INVx1_ASAP7_75t_SL g3717 ( 
.A(n_3611),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3600),
.B(n_3579),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3624),
.Y(n_3719)
);

INVx1_ASAP7_75t_SL g3720 ( 
.A(n_3633),
.Y(n_3720)
);

INVxp67_ASAP7_75t_L g3721 ( 
.A(n_3633),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3609),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3603),
.B(n_3544),
.Y(n_3723)
);

OR2x2_ASAP7_75t_L g3724 ( 
.A(n_3717),
.B(n_3593),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_3717),
.B(n_3607),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3717),
.B(n_3605),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3687),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3680),
.B(n_3605),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3680),
.B(n_3608),
.Y(n_3729)
);

OAI22xp5_ASAP7_75t_SL g3730 ( 
.A1(n_3712),
.A2(n_3546),
.B1(n_3610),
.B2(n_3636),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3687),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3706),
.B(n_3608),
.Y(n_3732)
);

INVxp67_ASAP7_75t_SL g3733 ( 
.A(n_3671),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3687),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3706),
.B(n_3608),
.Y(n_3735)
);

OR2x2_ASAP7_75t_L g3736 ( 
.A(n_3720),
.B(n_3593),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3698),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3706),
.B(n_3603),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3694),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3694),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3706),
.B(n_3598),
.Y(n_3741)
);

HB1xp67_ASAP7_75t_L g3742 ( 
.A(n_3698),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3701),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3701),
.Y(n_3744)
);

OAI221xp5_ASAP7_75t_L g3745 ( 
.A1(n_3712),
.A2(n_3538),
.B1(n_3546),
.B2(n_3610),
.C(n_3636),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3670),
.B(n_3661),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3718),
.B(n_3598),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3697),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3718),
.B(n_3599),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3694),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3694),
.Y(n_3751)
);

NAND3xp33_ASAP7_75t_SL g3752 ( 
.A(n_3712),
.B(n_3538),
.C(n_3542),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_3712),
.B(n_3638),
.Y(n_3753)
);

BUFx2_ASAP7_75t_L g3754 ( 
.A(n_3670),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3718),
.B(n_3599),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3697),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3694),
.Y(n_3757)
);

OR2x2_ASAP7_75t_L g3758 ( 
.A(n_3720),
.B(n_3597),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_3686),
.B(n_3595),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3718),
.B(n_3655),
.Y(n_3760)
);

HB1xp67_ASAP7_75t_L g3761 ( 
.A(n_3670),
.Y(n_3761)
);

INVx4_ASAP7_75t_L g3762 ( 
.A(n_3704),
.Y(n_3762)
);

AND2x2_ASAP7_75t_SL g3763 ( 
.A(n_3681),
.B(n_3630),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3720),
.B(n_3655),
.Y(n_3764)
);

NAND2x1p5_ASAP7_75t_L g3765 ( 
.A(n_3671),
.B(n_3673),
.Y(n_3765)
);

NAND2x1_ASAP7_75t_SL g3766 ( 
.A(n_3671),
.B(n_3661),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3670),
.Y(n_3767)
);

OAI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3686),
.A2(n_3546),
.B(n_3595),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3681),
.B(n_3546),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3681),
.B(n_3546),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3689),
.B(n_3656),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3689),
.B(n_3656),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3716),
.B(n_3597),
.Y(n_3773)
);

NAND2xp33_ASAP7_75t_R g3774 ( 
.A(n_3686),
.B(n_3644),
.Y(n_3774)
);

AND2x4_ASAP7_75t_L g3775 ( 
.A(n_3670),
.B(n_3661),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3742),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3752),
.B(n_3638),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3742),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3741),
.B(n_3617),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3741),
.B(n_3617),
.Y(n_3780)
);

OR2x2_ASAP7_75t_L g3781 ( 
.A(n_3736),
.B(n_3679),
.Y(n_3781)
);

AND2x4_ASAP7_75t_SL g3782 ( 
.A(n_3726),
.B(n_3618),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3747),
.B(n_3661),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3747),
.B(n_3663),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3766),
.Y(n_3785)
);

NOR2xp33_ASAP7_75t_L g3786 ( 
.A(n_3752),
.B(n_3638),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3761),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3761),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3749),
.B(n_3663),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3749),
.B(n_3663),
.Y(n_3790)
);

AND2x4_ASAP7_75t_L g3791 ( 
.A(n_3727),
.B(n_3676),
.Y(n_3791)
);

INVx3_ASAP7_75t_L g3792 ( 
.A(n_3762),
.Y(n_3792)
);

AND2x4_ASAP7_75t_SL g3793 ( 
.A(n_3726),
.B(n_3618),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3766),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3767),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3755),
.B(n_3738),
.Y(n_3796)
);

AND2x4_ASAP7_75t_SL g3797 ( 
.A(n_3732),
.B(n_3618),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3755),
.B(n_3738),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3760),
.B(n_3663),
.Y(n_3799)
);

OAI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3724),
.A2(n_3561),
.B1(n_3644),
.B2(n_3568),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3765),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3767),
.Y(n_3802)
);

NOR2x1_ASAP7_75t_L g3803 ( 
.A(n_3736),
.B(n_3696),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3763),
.B(n_3681),
.Y(n_3804)
);

INVx2_ASAP7_75t_SL g3805 ( 
.A(n_3727),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3760),
.B(n_3664),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3754),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3764),
.B(n_3664),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3764),
.B(n_3664),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3765),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3765),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3754),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3763),
.B(n_3681),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3727),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3779),
.B(n_3771),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3779),
.B(n_3771),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3805),
.Y(n_3817)
);

HB1xp67_ASAP7_75t_L g3818 ( 
.A(n_3807),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3780),
.B(n_3772),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3780),
.B(n_3772),
.Y(n_3820)
);

OR2x2_ASAP7_75t_L g3821 ( 
.A(n_3804),
.B(n_3724),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3805),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3805),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3807),
.Y(n_3824)
);

BUFx2_ASAP7_75t_L g3825 ( 
.A(n_3803),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3796),
.B(n_3725),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3803),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3796),
.B(n_3725),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3798),
.B(n_3625),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3812),
.Y(n_3830)
);

OR2x2_ASAP7_75t_L g3831 ( 
.A(n_3804),
.B(n_3813),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3798),
.B(n_3732),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3808),
.B(n_3625),
.Y(n_3833)
);

OR2x2_ASAP7_75t_L g3834 ( 
.A(n_3813),
.B(n_3758),
.Y(n_3834)
);

OR2x2_ASAP7_75t_L g3835 ( 
.A(n_3812),
.B(n_3758),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3808),
.B(n_3809),
.Y(n_3836)
);

AND2x4_ASAP7_75t_SL g3837 ( 
.A(n_3806),
.B(n_3618),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3787),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3809),
.B(n_3735),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3787),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3829),
.B(n_3615),
.Y(n_3841)
);

OR2x2_ASAP7_75t_L g3842 ( 
.A(n_3832),
.B(n_3815),
.Y(n_3842)
);

NOR2xp33_ASAP7_75t_L g3843 ( 
.A(n_3825),
.B(n_3618),
.Y(n_3843)
);

INVxp67_ASAP7_75t_SL g3844 ( 
.A(n_3825),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3829),
.B(n_3806),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3833),
.B(n_3735),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3820),
.B(n_3602),
.Y(n_3847)
);

OR2x2_ASAP7_75t_L g3848 ( 
.A(n_3835),
.B(n_3602),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3833),
.B(n_3665),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3836),
.B(n_3657),
.Y(n_3850)
);

NOR3x1_ASAP7_75t_L g3851 ( 
.A(n_3839),
.B(n_3768),
.C(n_3745),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3817),
.Y(n_3852)
);

OR2x6_ASAP7_75t_L g3853 ( 
.A(n_3827),
.B(n_3618),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3826),
.B(n_3783),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3826),
.B(n_3783),
.Y(n_3855)
);

AND2x4_ASAP7_75t_L g3856 ( 
.A(n_3822),
.B(n_3797),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3836),
.B(n_3657),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3823),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3828),
.B(n_3784),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3828),
.B(n_3784),
.Y(n_3860)
);

INVxp67_ASAP7_75t_L g3861 ( 
.A(n_3848),
.Y(n_3861)
);

OR2x2_ASAP7_75t_L g3862 ( 
.A(n_3846),
.B(n_3773),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3856),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3844),
.B(n_3763),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3845),
.B(n_3816),
.Y(n_3865)
);

OR2x2_ASAP7_75t_L g3866 ( 
.A(n_3855),
.B(n_3773),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3845),
.B(n_3816),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3844),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3856),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3854),
.B(n_3827),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3841),
.B(n_3819),
.Y(n_3871)
);

A2O1A1Ixp33_ASAP7_75t_L g3872 ( 
.A1(n_3843),
.A2(n_3686),
.B(n_3786),
.C(n_3777),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3854),
.B(n_3721),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3859),
.B(n_3721),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3856),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3853),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3849),
.B(n_3819),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3865),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3867),
.B(n_3850),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3871),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3873),
.B(n_3835),
.Y(n_3881)
);

INVx1_ASAP7_75t_SL g3882 ( 
.A(n_3877),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3863),
.B(n_3782),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3869),
.B(n_3857),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3875),
.B(n_3859),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3868),
.B(n_3753),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3873),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3866),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_L g3889 ( 
.A(n_3874),
.B(n_3710),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3885),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3879),
.Y(n_3891)
);

OAI322xp33_ASAP7_75t_L g3892 ( 
.A1(n_3889),
.A2(n_3777),
.A3(n_3786),
.B1(n_3800),
.B2(n_3688),
.C1(n_3759),
.C2(n_3679),
.Y(n_3892)
);

OAI22xp5_ASAP7_75t_L g3893 ( 
.A1(n_3882),
.A2(n_3710),
.B1(n_3571),
.B2(n_3562),
.Y(n_3893)
);

AND2x4_ASAP7_75t_L g3894 ( 
.A(n_3884),
.B(n_3860),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3882),
.B(n_3753),
.Y(n_3895)
);

NAND3xp33_ASAP7_75t_L g3896 ( 
.A(n_3881),
.B(n_3843),
.C(n_3872),
.Y(n_3896)
);

OAI322xp33_ASAP7_75t_L g3897 ( 
.A1(n_3886),
.A2(n_3800),
.A3(n_3688),
.B1(n_3679),
.B2(n_3769),
.C1(n_3770),
.C2(n_3781),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3894),
.B(n_3860),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3892),
.B(n_3874),
.Y(n_3899)
);

AOI22xp5_ASAP7_75t_L g3900 ( 
.A1(n_3891),
.A2(n_3730),
.B1(n_3649),
.B2(n_3647),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3890),
.B(n_3782),
.Y(n_3901)
);

AOI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3893),
.A2(n_3730),
.B1(n_3649),
.B2(n_3647),
.Y(n_3902)
);

AOI221xp5_ASAP7_75t_L g3903 ( 
.A1(n_3897),
.A2(n_3703),
.B1(n_3769),
.B2(n_3770),
.C(n_3745),
.Y(n_3903)
);

HB1xp67_ASAP7_75t_L g3904 ( 
.A(n_3895),
.Y(n_3904)
);

OAI22xp33_ASAP7_75t_SL g3905 ( 
.A1(n_3896),
.A2(n_3864),
.B1(n_3794),
.B2(n_3785),
.Y(n_3905)
);

OAI22xp33_ASAP7_75t_L g3906 ( 
.A1(n_3895),
.A2(n_3644),
.B1(n_3774),
.B2(n_3688),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3895),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3895),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3895),
.Y(n_3909)
);

AOI21xp33_ASAP7_75t_SL g3910 ( 
.A1(n_3895),
.A2(n_3864),
.B(n_3834),
.Y(n_3910)
);

INVx1_ASAP7_75t_SL g3911 ( 
.A(n_3898),
.Y(n_3911)
);

OAI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3900),
.A2(n_3861),
.B(n_3902),
.Y(n_3912)
);

OAI22xp5_ASAP7_75t_L g3913 ( 
.A1(n_3901),
.A2(n_3660),
.B1(n_3667),
.B2(n_3631),
.Y(n_3913)
);

NOR2xp33_ASAP7_75t_L g3914 ( 
.A(n_3910),
.B(n_3847),
.Y(n_3914)
);

A2O1A1Ixp33_ASAP7_75t_L g3915 ( 
.A1(n_3899),
.A2(n_3797),
.B(n_3793),
.C(n_3782),
.Y(n_3915)
);

O2A1O1Ixp33_ASAP7_75t_L g3916 ( 
.A1(n_3905),
.A2(n_3818),
.B(n_3870),
.C(n_3830),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3903),
.B(n_3728),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3906),
.B(n_3728),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3904),
.B(n_3729),
.Y(n_3919)
);

OR2x2_ASAP7_75t_L g3920 ( 
.A(n_3907),
.B(n_3781),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3908),
.B(n_3729),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3909),
.Y(n_3922)
);

OAI22xp33_ASAP7_75t_L g3923 ( 
.A1(n_3900),
.A2(n_3669),
.B1(n_3644),
.B2(n_3707),
.Y(n_3923)
);

AOI32xp33_ASAP7_75t_L g3924 ( 
.A1(n_3899),
.A2(n_3793),
.A3(n_3797),
.B1(n_3837),
.B2(n_3674),
.Y(n_3924)
);

O2A1O1Ixp33_ASAP7_75t_L g3925 ( 
.A1(n_3905),
.A2(n_3870),
.B(n_3830),
.C(n_3886),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3898),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3900),
.B(n_3837),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3900),
.B(n_3878),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_3898),
.B(n_3880),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_SL g3930 ( 
.A1(n_3899),
.A2(n_3674),
.B1(n_3671),
.B2(n_3673),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_L g3931 ( 
.A(n_3898),
.B(n_3862),
.Y(n_3931)
);

OAI32xp33_ASAP7_75t_L g3932 ( 
.A1(n_3898),
.A2(n_3834),
.A3(n_3821),
.B1(n_3696),
.B2(n_3883),
.Y(n_3932)
);

OAI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_3915),
.A2(n_3842),
.B(n_3887),
.Y(n_3933)
);

AOI221xp5_ASAP7_75t_L g3934 ( 
.A1(n_3932),
.A2(n_3793),
.B1(n_3858),
.B2(n_3852),
.C(n_3756),
.Y(n_3934)
);

AOI22xp5_ASAP7_75t_L g3935 ( 
.A1(n_3914),
.A2(n_3929),
.B1(n_3931),
.B2(n_3703),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3916),
.Y(n_3936)
);

INVxp67_ASAP7_75t_L g3937 ( 
.A(n_3919),
.Y(n_3937)
);

OAI21xp5_ASAP7_75t_SL g3938 ( 
.A1(n_3924),
.A2(n_3778),
.B(n_3776),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3925),
.A2(n_3888),
.B(n_3821),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3928),
.B(n_3666),
.Y(n_3940)
);

AOI21xp5_ASAP7_75t_L g3941 ( 
.A1(n_3927),
.A2(n_3831),
.B(n_3876),
.Y(n_3941)
);

OAI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3913),
.A2(n_3768),
.B(n_3824),
.Y(n_3942)
);

OAI211xp5_ASAP7_75t_L g3943 ( 
.A1(n_3930),
.A2(n_3840),
.B(n_3838),
.C(n_3776),
.Y(n_3943)
);

O2A1O1Ixp5_ASAP7_75t_L g3944 ( 
.A1(n_3912),
.A2(n_3778),
.B(n_3762),
.C(n_3707),
.Y(n_3944)
);

AOI31xp33_ASAP7_75t_L g3945 ( 
.A1(n_3920),
.A2(n_3840),
.A3(n_3814),
.B(n_3831),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3921),
.Y(n_3946)
);

O2A1O1Ixp33_ASAP7_75t_L g3947 ( 
.A1(n_3917),
.A2(n_3853),
.B(n_3792),
.C(n_3814),
.Y(n_3947)
);

OAI211xp5_ASAP7_75t_SL g3948 ( 
.A1(n_3918),
.A2(n_3792),
.B(n_3788),
.C(n_3795),
.Y(n_3948)
);

O2A1O1Ixp5_ASAP7_75t_L g3949 ( 
.A1(n_3923),
.A2(n_3762),
.B(n_3788),
.C(n_3802),
.Y(n_3949)
);

NOR3xp33_ASAP7_75t_L g3950 ( 
.A(n_3911),
.B(n_3792),
.C(n_3795),
.Y(n_3950)
);

AOI21xp33_ASAP7_75t_SL g3951 ( 
.A1(n_3926),
.A2(n_3853),
.B(n_3802),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3922),
.B(n_3851),
.Y(n_3952)
);

OAI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3917),
.A2(n_3669),
.B1(n_3719),
.B2(n_3716),
.Y(n_3953)
);

AOI222xp33_ASAP7_75t_L g3954 ( 
.A1(n_3912),
.A2(n_3674),
.B1(n_3673),
.B2(n_3703),
.C1(n_3699),
.C2(n_3748),
.Y(n_3954)
);

AOI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3914),
.A2(n_3703),
.B1(n_3669),
.B2(n_3789),
.Y(n_3955)
);

OAI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3915),
.A2(n_3756),
.B(n_3748),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3924),
.B(n_3792),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3932),
.A2(n_3810),
.B(n_3801),
.Y(n_3958)
);

AOI22xp5_ASAP7_75t_L g3959 ( 
.A1(n_3940),
.A2(n_3719),
.B1(n_3716),
.B2(n_3669),
.Y(n_3959)
);

BUFx2_ASAP7_75t_L g3960 ( 
.A(n_3956),
.Y(n_3960)
);

O2A1O1Ixp5_ASAP7_75t_L g3961 ( 
.A1(n_3943),
.A2(n_3762),
.B(n_3811),
.C(n_3810),
.Y(n_3961)
);

AOI221xp5_ASAP7_75t_L g3962 ( 
.A1(n_3953),
.A2(n_3791),
.B1(n_3785),
.B2(n_3794),
.C(n_3811),
.Y(n_3962)
);

NOR2xp33_ASAP7_75t_L g3963 ( 
.A(n_3955),
.B(n_3716),
.Y(n_3963)
);

NAND3xp33_ASAP7_75t_SL g3964 ( 
.A(n_3934),
.B(n_3719),
.C(n_3801),
.Y(n_3964)
);

OAI211xp5_ASAP7_75t_SL g3965 ( 
.A1(n_3935),
.A2(n_3794),
.B(n_3785),
.C(n_3801),
.Y(n_3965)
);

NAND2xp33_ASAP7_75t_R g3966 ( 
.A(n_3951),
.B(n_3791),
.Y(n_3966)
);

AOI222xp33_ASAP7_75t_L g3967 ( 
.A1(n_3936),
.A2(n_3674),
.B1(n_3673),
.B2(n_3699),
.C1(n_3672),
.C2(n_3675),
.Y(n_3967)
);

AOI211xp5_ASAP7_75t_L g3968 ( 
.A1(n_3938),
.A2(n_3811),
.B(n_3810),
.C(n_3743),
.Y(n_3968)
);

OAI221xp5_ASAP7_75t_L g3969 ( 
.A1(n_3942),
.A2(n_3719),
.B1(n_3744),
.B2(n_3737),
.C(n_3743),
.Y(n_3969)
);

AOI31xp33_ASAP7_75t_L g3970 ( 
.A1(n_3939),
.A2(n_3941),
.A3(n_3952),
.B(n_3933),
.Y(n_3970)
);

AOI221xp5_ASAP7_75t_L g3971 ( 
.A1(n_3945),
.A2(n_3947),
.B1(n_3948),
.B2(n_3950),
.C(n_3958),
.Y(n_3971)
);

AOI321xp33_ASAP7_75t_L g3972 ( 
.A1(n_3946),
.A2(n_3791),
.A3(n_3734),
.B1(n_3731),
.B2(n_3737),
.C(n_3744),
.Y(n_3972)
);

AOI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3937),
.A2(n_3669),
.B1(n_3790),
.B2(n_3789),
.Y(n_3973)
);

OAI211xp5_ASAP7_75t_L g3974 ( 
.A1(n_3957),
.A2(n_3734),
.B(n_3731),
.C(n_3750),
.Y(n_3974)
);

OAI21xp33_ASAP7_75t_L g3975 ( 
.A1(n_3954),
.A2(n_3790),
.B(n_3799),
.Y(n_3975)
);

OAI211xp5_ASAP7_75t_SL g3976 ( 
.A1(n_3944),
.A2(n_3699),
.B(n_3696),
.C(n_3757),
.Y(n_3976)
);

AOI222xp33_ASAP7_75t_L g3977 ( 
.A1(n_3949),
.A2(n_3672),
.B1(n_3675),
.B2(n_3676),
.C1(n_3733),
.C2(n_3678),
.Y(n_3977)
);

OAI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3955),
.A2(n_3669),
.B1(n_3660),
.B2(n_3799),
.Y(n_3978)
);

AOI22xp33_ASAP7_75t_L g3979 ( 
.A1(n_3940),
.A2(n_3684),
.B1(n_3683),
.B2(n_3660),
.Y(n_3979)
);

NAND3xp33_ASAP7_75t_SL g3980 ( 
.A(n_3934),
.B(n_3740),
.C(n_3739),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3947),
.A2(n_3791),
.B(n_3750),
.C(n_3757),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3939),
.A2(n_3740),
.B(n_3739),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_SL g3983 ( 
.A1(n_3978),
.A2(n_3733),
.B1(n_3757),
.B2(n_3751),
.Y(n_3983)
);

AOI321xp33_ASAP7_75t_L g3984 ( 
.A1(n_3968),
.A2(n_3751),
.A3(n_3750),
.B1(n_3740),
.B2(n_3739),
.C(n_3675),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3982),
.A2(n_3751),
.B(n_3672),
.Y(n_3985)
);

NAND2xp33_ASAP7_75t_L g3986 ( 
.A(n_3975),
.B(n_3696),
.Y(n_3986)
);

AND3x1_ASAP7_75t_L g3987 ( 
.A(n_3971),
.B(n_3666),
.C(n_3689),
.Y(n_3987)
);

NOR3xp33_ASAP7_75t_L g3988 ( 
.A(n_3970),
.B(n_3551),
.C(n_3574),
.Y(n_3988)
);

OR3x1_ASAP7_75t_L g3989 ( 
.A(n_3964),
.B(n_3682),
.C(n_3693),
.Y(n_3989)
);

O2A1O1Ixp33_ASAP7_75t_L g3990 ( 
.A1(n_3981),
.A2(n_3676),
.B(n_3677),
.C(n_3678),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3959),
.B(n_3551),
.Y(n_3991)
);

NOR4xp25_ASAP7_75t_L g3992 ( 
.A(n_3965),
.B(n_3676),
.C(n_3682),
.D(n_3693),
.Y(n_3992)
);

AOI211xp5_ASAP7_75t_SL g3993 ( 
.A1(n_3974),
.A2(n_3689),
.B(n_3695),
.C(n_3692),
.Y(n_3993)
);

AOI21xp33_ASAP7_75t_SL g3994 ( 
.A1(n_3966),
.A2(n_3676),
.B(n_3702),
.Y(n_3994)
);

AOI221xp5_ASAP7_75t_L g3995 ( 
.A1(n_3969),
.A2(n_3775),
.B1(n_3746),
.B2(n_3682),
.C(n_3690),
.Y(n_3995)
);

AOI221x1_ASAP7_75t_L g3996 ( 
.A1(n_3980),
.A2(n_3775),
.B1(n_3746),
.B2(n_3690),
.C(n_3693),
.Y(n_3996)
);

O2A1O1Ixp33_ASAP7_75t_L g3997 ( 
.A1(n_3961),
.A2(n_3677),
.B(n_3678),
.C(n_3713),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3973),
.B(n_3555),
.Y(n_3998)
);

OAI211xp5_ASAP7_75t_L g3999 ( 
.A1(n_3962),
.A2(n_3678),
.B(n_3677),
.C(n_3713),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3994),
.B(n_3972),
.Y(n_4000)
);

OAI221xp5_ASAP7_75t_L g4001 ( 
.A1(n_3993),
.A2(n_3979),
.B1(n_3963),
.B2(n_3960),
.C(n_3976),
.Y(n_4001)
);

NAND3xp33_ASAP7_75t_L g4002 ( 
.A(n_3986),
.B(n_3967),
.C(n_3977),
.Y(n_4002)
);

OR3x1_ASAP7_75t_L g4003 ( 
.A(n_3998),
.B(n_3690),
.C(n_3711),
.Y(n_4003)
);

NAND4xp25_ASAP7_75t_L g4004 ( 
.A(n_3988),
.B(n_3775),
.C(n_3746),
.D(n_3695),
.Y(n_4004)
);

NOR2x1_ASAP7_75t_L g4005 ( 
.A(n_3989),
.B(n_3704),
.Y(n_4005)
);

NAND4xp25_ASAP7_75t_SL g4006 ( 
.A(n_3995),
.B(n_3702),
.C(n_3695),
.D(n_3692),
.Y(n_4006)
);

NOR4xp25_ASAP7_75t_L g4007 ( 
.A(n_3984),
.B(n_3677),
.C(n_3714),
.D(n_3711),
.Y(n_4007)
);

NOR2xp67_ASAP7_75t_SL g4008 ( 
.A(n_3985),
.B(n_3555),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3983),
.B(n_3746),
.Y(n_4009)
);

NAND5xp2_ASAP7_75t_L g4010 ( 
.A(n_3997),
.B(n_3702),
.C(n_3695),
.D(n_3692),
.E(n_3714),
.Y(n_4010)
);

INVx2_ASAP7_75t_L g4011 ( 
.A(n_3987),
.Y(n_4011)
);

NAND3xp33_ASAP7_75t_L g4012 ( 
.A(n_3991),
.B(n_3775),
.C(n_3692),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3990),
.Y(n_4013)
);

OAI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3999),
.A2(n_3992),
.B(n_3996),
.Y(n_4014)
);

AOI311xp33_ASAP7_75t_L g4015 ( 
.A1(n_4001),
.A2(n_3711),
.A3(n_3714),
.B(n_3722),
.C(n_3613),
.Y(n_4015)
);

NAND3xp33_ASAP7_75t_SL g4016 ( 
.A(n_4014),
.B(n_3702),
.C(n_3684),
.Y(n_4016)
);

NAND4xp25_ASAP7_75t_SL g4017 ( 
.A(n_4012),
.B(n_3684),
.C(n_3683),
.D(n_3691),
.Y(n_4017)
);

OAI211xp5_ASAP7_75t_L g4018 ( 
.A1(n_4009),
.A2(n_3691),
.B(n_3685),
.C(n_3683),
.Y(n_4018)
);

AOI211x1_ASAP7_75t_SL g4019 ( 
.A1(n_4002),
.A2(n_3685),
.B(n_3691),
.C(n_3709),
.Y(n_4019)
);

AOI221xp5_ASAP7_75t_L g4020 ( 
.A1(n_4006),
.A2(n_3685),
.B1(n_3691),
.B2(n_3704),
.C(n_3709),
.Y(n_4020)
);

NOR3xp33_ASAP7_75t_L g4021 ( 
.A(n_4000),
.B(n_3551),
.C(n_3570),
.Y(n_4021)
);

AOI22xp5_ASAP7_75t_L g4022 ( 
.A1(n_4004),
.A2(n_3634),
.B1(n_3639),
.B2(n_3627),
.Y(n_4022)
);

AOI211xp5_ASAP7_75t_L g4023 ( 
.A1(n_4010),
.A2(n_3683),
.B(n_3684),
.C(n_3723),
.Y(n_4023)
);

NOR3xp33_ASAP7_75t_L g4024 ( 
.A(n_4011),
.B(n_3551),
.C(n_3574),
.Y(n_4024)
);

NOR2x2_ASAP7_75t_L g4025 ( 
.A(n_4008),
.B(n_3570),
.Y(n_4025)
);

OAI21xp33_ASAP7_75t_SL g4026 ( 
.A1(n_4005),
.A2(n_3685),
.B(n_3723),
.Y(n_4026)
);

OAI221xp5_ASAP7_75t_L g4027 ( 
.A1(n_4007),
.A2(n_3704),
.B1(n_3708),
.B2(n_3709),
.C(n_3715),
.Y(n_4027)
);

XNOR2x1_ASAP7_75t_L g4028 ( 
.A(n_4013),
.B(n_3634),
.Y(n_4028)
);

NOR3xp33_ASAP7_75t_SL g4029 ( 
.A(n_4003),
.B(n_3722),
.C(n_3643),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_4008),
.B(n_3555),
.Y(n_4030)
);

AOI311xp33_ASAP7_75t_L g4031 ( 
.A1(n_4001),
.A2(n_3722),
.A3(n_3653),
.B(n_3651),
.C(n_3622),
.Y(n_4031)
);

NAND3xp33_ASAP7_75t_L g4032 ( 
.A(n_4002),
.B(n_3709),
.C(n_3708),
.Y(n_4032)
);

INVx2_ASAP7_75t_SL g4033 ( 
.A(n_4028),
.Y(n_4033)
);

AO22x1_ASAP7_75t_L g4034 ( 
.A1(n_4024),
.A2(n_3627),
.B1(n_3639),
.B2(n_3723),
.Y(n_4034)
);

NOR2x1_ASAP7_75t_L g4035 ( 
.A(n_4032),
.B(n_3704),
.Y(n_4035)
);

AOI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_4021),
.A2(n_4022),
.B1(n_4016),
.B2(n_4030),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_4025),
.Y(n_4037)
);

NOR3xp33_ASAP7_75t_L g4038 ( 
.A(n_4026),
.B(n_3723),
.C(n_3708),
.Y(n_4038)
);

OAI22x1_ASAP7_75t_L g4039 ( 
.A1(n_4017),
.A2(n_3640),
.B1(n_3621),
.B2(n_3648),
.Y(n_4039)
);

INVx1_ASAP7_75t_SL g4040 ( 
.A(n_4019),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_4023),
.B(n_3708),
.Y(n_4041)
);

OAI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_4027),
.A2(n_3715),
.B1(n_3700),
.B2(n_3637),
.Y(n_4042)
);

NOR2x1_ASAP7_75t_L g4043 ( 
.A(n_4018),
.B(n_3705),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_4029),
.B(n_3700),
.Y(n_4044)
);

AOI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_4020),
.A2(n_3715),
.B1(n_3700),
.B2(n_3705),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_4031),
.B(n_3619),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_4015),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_4028),
.Y(n_4048)
);

INVxp67_ASAP7_75t_L g4049 ( 
.A(n_4028),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_4034),
.Y(n_4050)
);

OR2x2_ASAP7_75t_L g4051 ( 
.A(n_4042),
.B(n_3700),
.Y(n_4051)
);

NOR3xp33_ASAP7_75t_L g4052 ( 
.A(n_4049),
.B(n_4033),
.C(n_4048),
.Y(n_4052)
);

NOR2x1_ASAP7_75t_L g4053 ( 
.A(n_4035),
.B(n_3705),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_4039),
.Y(n_4054)
);

INVx3_ASAP7_75t_L g4055 ( 
.A(n_4037),
.Y(n_4055)
);

NOR5xp2_ASAP7_75t_L g4056 ( 
.A(n_4047),
.B(n_3592),
.C(n_3623),
.D(n_3629),
.E(n_3653),
.Y(n_4056)
);

NAND4xp25_ASAP7_75t_SL g4057 ( 
.A(n_4036),
.B(n_3715),
.C(n_3700),
.D(n_3662),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_4046),
.B(n_3715),
.Y(n_4058)
);

NOR4xp75_ASAP7_75t_L g4059 ( 
.A(n_4041),
.B(n_3705),
.C(n_3637),
.D(n_3529),
.Y(n_4059)
);

NOR3xp33_ASAP7_75t_L g4060 ( 
.A(n_4040),
.B(n_3705),
.C(n_3565),
.Y(n_4060)
);

OAI211xp5_ASAP7_75t_SL g4061 ( 
.A1(n_4054),
.A2(n_4044),
.B(n_4043),
.C(n_4038),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_4060),
.B(n_4045),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_4052),
.B(n_3548),
.Y(n_4063)
);

NOR2xp67_ASAP7_75t_L g4064 ( 
.A(n_4057),
.B(n_3705),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4053),
.Y(n_4065)
);

O2A1O1Ixp5_ASAP7_75t_L g4066 ( 
.A1(n_4058),
.A2(n_3591),
.B(n_3594),
.C(n_3662),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_4063),
.B(n_4059),
.Y(n_4067)
);

BUFx2_ASAP7_75t_L g4068 ( 
.A(n_4065),
.Y(n_4068)
);

NAND2x1p5_ASAP7_75t_L g4069 ( 
.A(n_4064),
.B(n_4055),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4068),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_4067),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_4070),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_4072),
.A2(n_4050),
.B1(n_4071),
.B2(n_4061),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4073),
.B(n_4051),
.Y(n_4074)
);

AOI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_4074),
.A2(n_4062),
.B1(n_4069),
.B2(n_4056),
.Y(n_4075)
);

XOR2xp5_ASAP7_75t_L g4076 ( 
.A(n_4075),
.B(n_4066),
.Y(n_4076)
);

AOI221xp5_ASAP7_75t_L g4077 ( 
.A1(n_4076),
.A2(n_3629),
.B1(n_3609),
.B2(n_3613),
.C(n_3614),
.Y(n_4077)
);

OAI332xp33_ASAP7_75t_L g4078 ( 
.A1(n_4077),
.A2(n_3662),
.A3(n_3594),
.B1(n_3591),
.B2(n_3632),
.B3(n_3614),
.C1(n_3622),
.C2(n_3623),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_4078),
.Y(n_4079)
);

OAI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_4079),
.A2(n_3591),
.B(n_3594),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4080),
.Y(n_4081)
);

AOI22xp33_ASAP7_75t_L g4082 ( 
.A1(n_4081),
.A2(n_3668),
.B1(n_3626),
.B2(n_3646),
.Y(n_4082)
);

OAI221xp5_ASAP7_75t_R g4083 ( 
.A1(n_4082),
.A2(n_3590),
.B1(n_3668),
.B2(n_3659),
.C(n_3626),
.Y(n_4083)
);

OAI221xp5_ASAP7_75t_R g4084 ( 
.A1(n_4082),
.A2(n_3590),
.B1(n_3659),
.B2(n_3626),
.C(n_3645),
.Y(n_4084)
);

AOI22xp5_ASAP7_75t_L g4085 ( 
.A1(n_4083),
.A2(n_3626),
.B1(n_3659),
.B2(n_3590),
.Y(n_4085)
);

AOI211xp5_ASAP7_75t_L g4086 ( 
.A1(n_4085),
.A2(n_4084),
.B(n_3643),
.C(n_3632),
.Y(n_4086)
);


endmodule