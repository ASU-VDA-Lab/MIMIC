module fake_jpeg_11848_n_99 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_99);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_26),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_13),
.B1(n_22),
.B2(n_20),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_13),
.B1(n_11),
.B2(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_17),
.B1(n_21),
.B2(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_36),
.B1(n_28),
.B2(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_39),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_18),
.B1(n_14),
.B2(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_34),
.B1(n_38),
.B2(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_10),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_34),
.Y(n_55)
);

A2O1A1O1Ixp25_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_48),
.B(n_51),
.C(n_52),
.D(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_51),
.B1(n_45),
.B2(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_35),
.B1(n_30),
.B2(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_72)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_59),
.B1(n_64),
.B2(n_45),
.Y(n_67)
);

AOI221xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.C(n_73),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_63),
.B(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_56),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_52),
.B(n_31),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_38),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_61),
.C(n_55),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_57),
.C(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_61),
.C(n_25),
.Y(n_80)
);

OAI221xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_74),
.B1(n_81),
.B2(n_73),
.C(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_90),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_82),
.B1(n_83),
.B2(n_78),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_89),
.B(n_4),
.C(n_5),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_66),
.B(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_7),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_7),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

NOR2xp67_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_92),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_5),
.C(n_6),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_96),
.Y(n_99)
);


endmodule