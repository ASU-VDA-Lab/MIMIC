module fake_jpeg_10824_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_31),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_16),
.B(n_35),
.C(n_34),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_52),
.B(n_49),
.C(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_13),
.B1(n_33),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_56),
.B1(n_42),
.B2(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_1),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_36),
.B1(n_11),
.B2(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_42),
.B2(n_48),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_74),
.B1(n_79),
.B2(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_23),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_4),
.B(n_5),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_80),
.C(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_7),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_7),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_24),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_92),
.SN(n_92)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_10),
.Y(n_88)
);

AO22x2_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_27),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_81),
.C(n_86),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_98),
.C(n_99),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_91),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_96),
.B(n_89),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_94),
.C(n_92),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_101),
.Y(n_102)
);

AOI211xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_100),
.B(n_92),
.C(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_90),
.C(n_95),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_85),
.Y(n_106)
);


endmodule