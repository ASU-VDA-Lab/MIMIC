module fake_ariane_1551_n_185 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_185);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_185;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_174;
wire n_100;
wire n_132;
wire n_62;
wire n_147;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_82;
wire n_178;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_101;
wire n_94;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_87;
wire n_81;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVxp33_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_8),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_53),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_0),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_101),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_73),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_65),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_54),
.B1(n_85),
.B2(n_84),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_74),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_75),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_115),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_93),
.Y(n_127)
);

NOR2xp67_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_91),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_113),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_69),
.B(n_57),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_81),
.B(n_77),
.C(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_80),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_83),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_104),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_131),
.B(n_136),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_124),
.B(n_129),
.Y(n_148)
);

OAI21x1_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_124),
.B(n_129),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_133),
.Y(n_150)
);

AO21x2_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_6),
.B(n_7),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_9),
.B(n_11),
.Y(n_154)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_138),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_153),
.B(n_154),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_151),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_171),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_176),
.Y(n_177)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.C(n_38),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AO22x2_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_47),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_50),
.B(n_51),
.Y(n_185)
);


endmodule