module fake_netlist_6_819_n_1861 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1861);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1861;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_116),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_11),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_89),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_44),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_119),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_6),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_174),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_106),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_70),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_84),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_28),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_136),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_93),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_95),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_83),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_44),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_151),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_158),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_54),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_109),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_38),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_186),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_118),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_50),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_144),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_65),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_124),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_107),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_75),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_182),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_178),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_150),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_33),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_112),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_8),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_139),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_87),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_101),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_143),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_30),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_61),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_40),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_52),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_130),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_96),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_59),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_64),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_39),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_131),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_3),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_53),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_33),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_66),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_61),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_42),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_35),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_54),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_1),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_43),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_20),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_169),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_195),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_20),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_69),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_180),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_164),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_155),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_137),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_62),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_86),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_114),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_120),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_42),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_17),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_36),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_52),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_71),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_176),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_73),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_88),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_38),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_103),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_59),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_50),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_15),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_123),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_135),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_45),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_77),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_162),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_35),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_53),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_172),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_152),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_41),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_60),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_41),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_115),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_185),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_6),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_142),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_17),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_10),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_43),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_32),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_51),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_110),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_19),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_188),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_133),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_128),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_19),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_105),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_196),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_125),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_166),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_111),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_80),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_27),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_7),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_9),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_56),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_92),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_51),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_10),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_39),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_16),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_72),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_190),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_99),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_13),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_12),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_141),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_108),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_7),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_138),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_173),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_82),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_5),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_49),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_117),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_145),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_159),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_168),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_56),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_94),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_270),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_347),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_244),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_245),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_270),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_251),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_254),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_270),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_331),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_328),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_341),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_293),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_203),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_270),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_300),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_206),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_256),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_236),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_220),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_231),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_257),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_255),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_238),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_255),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_260),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_241),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_202),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_259),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_268),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_217),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_248),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_275),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_252),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_204),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_269),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_276),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_279),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_236),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_322),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_278),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_285),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_280),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_283),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_307),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_289),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_236),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_294),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_296),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_329),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_303),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_326),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_354),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_309),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_364),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_217),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_240),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_287),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_377),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_318),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_323),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_288),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_389),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_325),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_292),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_295),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_330),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_233),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_297),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_353),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_357),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_365),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_370),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_380),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_348),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_348),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_298),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_234),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_211),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_299),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_313),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_211),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_357),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_314),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_357),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_367),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_315),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_229),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_240),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_209),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_401),
.A2(n_215),
.B1(n_391),
.B2(n_369),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_243),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_243),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_473),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_431),
.B(n_249),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_394),
.B(n_402),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_435),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_393),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_216),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_249),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_411),
.A2(n_422),
.B(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_393),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_439),
.A2(n_277),
.B1(n_337),
.B2(n_214),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_223),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_461),
.B(n_229),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_444),
.B(n_247),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_397),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_400),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_422),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

CKINVDCx11_ASAP7_75t_R g523 ( 
.A(n_451),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_412),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_459),
.B(n_253),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_414),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_461),
.B(n_247),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_395),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_405),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_484),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_415),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_404),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_433),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_403),
.B(n_199),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_418),
.B(n_216),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_410),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_406),
.B(n_352),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_419),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_496),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_485),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_433),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_395),
.B(n_374),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_420),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_427),
.Y(n_553)
);

AND3x1_ASAP7_75t_L g554 ( 
.A(n_462),
.B(n_383),
.C(n_222),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_396),
.B(n_362),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_396),
.B(n_383),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_429),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_464),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_398),
.B(n_375),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_485),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

INVx6_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_492),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_409),
.B(n_208),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_491),
.B(n_199),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_436),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

CKINVDCx11_ASAP7_75t_R g572 ( 
.A(n_440),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_488),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_441),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_398),
.B(n_213),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_442),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_448),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_416),
.B(n_200),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_449),
.A2(n_350),
.B1(n_339),
.B2(n_366),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_511),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_525),
.B(n_399),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_520),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_501),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_514),
.B(n_399),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_507),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_531),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_514),
.B(n_413),
.Y(n_593)
);

BUFx6f_ASAP7_75t_SL g594 ( 
.A(n_566),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_507),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_533),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_555),
.B(n_413),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_520),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_526),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_545),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

AND3x2_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_503),
.C(n_530),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_501),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_554),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_425),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_508),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_526),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_561),
.B(n_425),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_512),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_520),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_512),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_499),
.B(n_432),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_535),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_542),
.B(n_479),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_SL g618 ( 
.A(n_566),
.B(n_432),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_518),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_542),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_500),
.B(n_434),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_551),
.B(n_434),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_515),
.B(n_479),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_516),
.B(n_437),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_575),
.B(n_437),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_567),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_543),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_515),
.B(n_480),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_509),
.B(n_216),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_564),
.B(n_481),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_564),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_R g637 ( 
.A(n_530),
.B(n_445),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_521),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_499),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_509),
.B(n_216),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_550),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_510),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_445),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_510),
.B(n_446),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_510),
.A2(n_453),
.B1(n_455),
.B2(n_452),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_550),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_550),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_550),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_519),
.A2(n_538),
.B1(n_569),
.B2(n_446),
.Y(n_651)
);

INVx8_ASAP7_75t_L g652 ( 
.A(n_509),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_521),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_564),
.B(n_481),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_524),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_558),
.B(n_463),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_557),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_503),
.B(n_463),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_509),
.B(n_216),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_521),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_515),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_528),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_527),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_527),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_539),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_557),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_557),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_564),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_537),
.B(n_467),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_497),
.B(n_467),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_528),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_547),
.B(n_470),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_536),
.Y(n_675)
);

BUFx6f_ASAP7_75t_SL g676 ( 
.A(n_536),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_531),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_529),
.A2(n_466),
.B1(n_469),
.B2(n_465),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_506),
.B(n_470),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_513),
.B(n_482),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_557),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_557),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_549),
.A2(n_571),
.B1(n_574),
.B2(n_570),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_532),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_537),
.B(n_498),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_528),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_576),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_522),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_537),
.B(n_471),
.Y(n_691)
);

AO21x2_ASAP7_75t_L g692 ( 
.A1(n_504),
.A2(n_227),
.B(n_226),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_534),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_577),
.B(n_471),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_548),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_534),
.B(n_474),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_534),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_532),
.B(n_474),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_578),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_546),
.B(n_483),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_546),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_546),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_578),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_578),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_578),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_578),
.B(n_483),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_556),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_581),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_562),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_562),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_541),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_573),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_573),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_509),
.A2(n_493),
.B1(n_490),
.B2(n_486),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_580),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

BUFx6f_ASAP7_75t_SL g722 ( 
.A(n_509),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_560),
.B(n_443),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_572),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_563),
.Y(n_725)
);

INVx6_ASAP7_75t_L g726 ( 
.A(n_540),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_563),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_568),
.A2(n_235),
.B(n_230),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_568),
.A2(n_351),
.B1(n_316),
.B2(n_349),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_621),
.B(n_265),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_621),
.A2(n_486),
.B1(n_487),
.B2(n_493),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_629),
.B(n_487),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_588),
.B(n_490),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_661),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_593),
.B(n_489),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_640),
.B(n_265),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_592),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_640),
.B(n_265),
.Y(n_738)
);

NOR2x1_ASAP7_75t_L g739 ( 
.A(n_597),
.B(n_239),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_635),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_592),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_617),
.B(n_423),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_725),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_643),
.B(n_265),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_661),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_643),
.B(n_242),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_609),
.B(n_552),
.C(n_541),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_696),
.B(n_263),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_656),
.B(n_447),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_617),
.B(n_628),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_717),
.B(n_645),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_635),
.B(n_482),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_669),
.B(n_691),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_630),
.B(n_552),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_589),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_680),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_728),
.A2(n_335),
.B1(n_384),
.B2(n_360),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_596),
.B(n_267),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_709),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_606),
.B(n_200),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_633),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_709),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_633),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_596),
.B(n_599),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_675),
.B(n_450),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_627),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_712),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_712),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_599),
.B(n_271),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_583),
.B(n_201),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_613),
.B(n_335),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_637),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_713),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_627),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_713),
.Y(n_775)
);

OAI221xp5_ASAP7_75t_L g776 ( 
.A1(n_647),
.A2(n_458),
.B1(n_472),
.B2(n_478),
.C(n_475),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_646),
.B(n_201),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_697),
.B(n_237),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_601),
.B(n_602),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_625),
.B(n_205),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_674),
.B(n_205),
.Y(n_781)
);

AO22x2_ASAP7_75t_L g782 ( 
.A1(n_670),
.A2(n_286),
.B1(n_291),
.B2(n_304),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_715),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_605),
.A2(n_454),
.B1(n_457),
.B2(n_468),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_688),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_695),
.B(n_207),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_675),
.B(n_207),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_602),
.B(n_607),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_715),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_L g790 ( 
.A(n_651),
.B(n_595),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_708),
.B(n_246),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_687),
.B(n_210),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_607),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_680),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_610),
.B(n_308),
.Y(n_795)
);

BUFx4f_ASAP7_75t_L g796 ( 
.A(n_635),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_SL g797 ( 
.A(n_636),
.B(n_668),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_605),
.A2(n_266),
.B1(n_262),
.B2(n_261),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_610),
.B(n_311),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_589),
.B(n_480),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_612),
.B(n_324),
.Y(n_801)
);

NOR3xp33_ASAP7_75t_L g802 ( 
.A(n_658),
.B(n_559),
.C(n_553),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_612),
.B(n_343),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_SL g804 ( 
.A1(n_711),
.A2(n_553),
.B1(n_559),
.B2(n_385),
.Y(n_804)
);

OAI221xp5_ASAP7_75t_L g805 ( 
.A1(n_678),
.A2(n_363),
.B1(n_355),
.B2(n_359),
.C(n_381),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_614),
.B(n_565),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_639),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_702),
.B(n_250),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_SL g809 ( 
.A1(n_711),
.A2(n_372),
.B1(n_369),
.B2(n_371),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_688),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_716),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_687),
.B(n_335),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_623),
.B(n_210),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_723),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_635),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_595),
.B(n_212),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_690),
.B(n_335),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_716),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_619),
.B(n_565),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_619),
.B(n_258),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_620),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_728),
.A2(n_384),
.B1(n_371),
.B2(n_372),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_652),
.B(n_264),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_724),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_719),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_620),
.B(n_272),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_723),
.B(n_523),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_582),
.B(n_384),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_644),
.A2(n_332),
.B(n_273),
.C(n_274),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_644),
.B(n_281),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_655),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_655),
.B(n_282),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_636),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_663),
.B(n_284),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_719),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_664),
.B(n_290),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_724),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_720),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_720),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_594),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_664),
.A2(n_426),
.B(n_428),
.C(n_336),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_654),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_665),
.A2(n_345),
.B(n_306),
.C(n_310),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_690),
.B(n_384),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_728),
.A2(n_385),
.B1(n_386),
.B2(n_391),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_636),
.B(n_212),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_654),
.B(n_683),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_710),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_668),
.B(n_586),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_584),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_685),
.B(n_718),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_668),
.B(n_618),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_654),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_693),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_654),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_639),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_679),
.B(n_218),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_729),
.B(n_218),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_721),
.B(n_301),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_721),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_594),
.B(n_219),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_L g862 ( 
.A(n_680),
.B(n_344),
.C(n_338),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_700),
.B(n_0),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_587),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_677),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_727),
.B(n_219),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_L g867 ( 
.A1(n_594),
.A2(n_386),
.B1(n_334),
.B2(n_333),
.C(n_327),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_727),
.B(n_221),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_705),
.B(n_221),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_586),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_603),
.B(n_224),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_694),
.B(n_698),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_694),
.B(n_302),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_676),
.B(n_224),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_705),
.B(n_225),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_587),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_692),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_604),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_L g879 ( 
.A(n_652),
.B(n_305),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_698),
.B(n_312),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_582),
.Y(n_881)
);

BUFx12f_ASAP7_75t_SL g882 ( 
.A(n_752),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_749),
.B(n_686),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_740),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_749),
.B(n_692),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_754),
.B(n_604),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_766),
.Y(n_887)
);

BUFx4f_ASAP7_75t_L g888 ( 
.A(n_740),
.Y(n_888)
);

AO22x1_ASAP7_75t_L g889 ( 
.A1(n_858),
.A2(n_684),
.B1(n_228),
.B2(n_225),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_796),
.B(n_706),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_781),
.B(n_692),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_833),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_774),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_735),
.B(n_676),
.Y(n_894)
);

NOR2x1p5_ASAP7_75t_L g895 ( 
.A(n_833),
.B(n_684),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_740),
.B(n_652),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_785),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_743),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_751),
.A2(n_676),
.B1(n_701),
.B2(n_707),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_862),
.B(n_361),
.C(n_232),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_865),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_850),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_864),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_742),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_872),
.A2(n_741),
.B(n_737),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_822),
.A2(n_616),
.B1(n_624),
.B2(n_600),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_714),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_864),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_SL g909 ( 
.A1(n_779),
.A2(n_701),
.B(n_707),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_847),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_SL g911 ( 
.A(n_786),
.B(n_228),
.C(n_232),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_750),
.B(n_660),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_735),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_815),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_848),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_730),
.A2(n_814),
.B(n_805),
.C(n_822),
.Y(n_916)
);

INVx4_ASAP7_75t_SL g917 ( 
.A(n_828),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_793),
.B(n_660),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_878),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_772),
.B(n_732),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_796),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_755),
.B(n_699),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_785),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_860),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_821),
.B(n_831),
.Y(n_925)
);

AOI221xp5_ASAP7_75t_SL g926 ( 
.A1(n_845),
.A2(n_659),
.B1(n_641),
.B2(n_634),
.C(n_600),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_761),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_755),
.B(n_800),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_800),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_876),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_851),
.B(n_671),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_763),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_759),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_842),
.Y(n_934)
);

BUFx8_ASAP7_75t_SL g935 ( 
.A(n_824),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_731),
.B(n_361),
.C(n_356),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_853),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_733),
.B(n_714),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_828),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_753),
.A2(n_704),
.B1(n_703),
.B2(n_699),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_855),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_847),
.B(n_703),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_762),
.Y(n_943)
);

INVx3_ASAP7_75t_SL g944 ( 
.A(n_837),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_770),
.B(n_714),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_SL g946 ( 
.A(n_770),
.B(n_780),
.C(n_857),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_856),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_752),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_SL g949 ( 
.A(n_784),
.B(n_858),
.C(n_867),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_734),
.B(n_672),
.Y(n_950)
);

NAND2x1p5_ASAP7_75t_L g951 ( 
.A(n_856),
.B(n_810),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_752),
.B(n_745),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_739),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_753),
.B(n_704),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_767),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_780),
.B(n_673),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_767),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_810),
.B(n_590),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_764),
.B(n_673),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_877),
.B(n_632),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_788),
.B(n_673),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_790),
.B(n_632),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_768),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_816),
.B(n_585),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_SL g965 ( 
.A1(n_863),
.A2(n_373),
.B1(n_356),
.B2(n_358),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_756),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_863),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_768),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_849),
.B(n_726),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_863),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_737),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_773),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_773),
.Y(n_973)
);

INVxp33_ASAP7_75t_L g974 ( 
.A(n_804),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_757),
.B(n_598),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_775),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_813),
.B(n_608),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_797),
.B(n_642),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_775),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_854),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_783),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_827),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_783),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_870),
.Y(n_984)
);

INVxp67_ASAP7_75t_SL g985 ( 
.A(n_881),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_857),
.B(n_590),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_789),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_794),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_787),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_789),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_811),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_811),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_854),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_818),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_746),
.B(n_598),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_818),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_881),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_825),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_845),
.A2(n_631),
.B(n_608),
.C(n_616),
.Y(n_999)
);

INVxp33_ASAP7_75t_L g1000 ( 
.A(n_871),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_741),
.B(n_642),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_813),
.B(n_590),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_SL g1003 ( 
.A1(n_782),
.A2(n_373),
.B1(n_392),
.B2(n_390),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_828),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_825),
.B(n_648),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_880),
.A2(n_666),
.B1(n_649),
.B2(n_657),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_835),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_820),
.B(n_826),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_838),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_838),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_830),
.B(n_832),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_839),
.Y(n_1012)
);

AND2x6_ASAP7_75t_L g1013 ( 
.A(n_839),
.B(n_650),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_792),
.Y(n_1014)
);

NOR2x1p5_ASAP7_75t_L g1015 ( 
.A(n_834),
.B(n_358),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_871),
.A2(n_378),
.B1(n_368),
.B2(n_379),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_806),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_782),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_852),
.B(n_657),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_819),
.B(n_666),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_782),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_828),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_840),
.B(n_667),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_836),
.B(n_667),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_760),
.B(n_615),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_758),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_748),
.B(n_611),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_828),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_795),
.B(n_611),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_769),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_799),
.A2(n_390),
.B1(n_368),
.B2(n_378),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_777),
.B(n_681),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_801),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_803),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_730),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_798),
.B(n_615),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_771),
.A2(n_744),
.B(n_736),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_866),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_817),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_817),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_812),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_812),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_873),
.B(n_681),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_884),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_919),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_931),
.A2(n_807),
.B(n_652),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_913),
.B(n_861),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_910),
.A2(n_771),
.B1(n_874),
.B2(n_861),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_910),
.B(n_913),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_SL g1050 ( 
.A(n_947),
.B(n_726),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_920),
.B(n_874),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_920),
.B(n_802),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_883),
.B(n_859),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1026),
.B(n_1030),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_884),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_971),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_985),
.A2(n_879),
.B(n_823),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1026),
.B(n_868),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_946),
.A2(n_843),
.B(n_829),
.C(n_778),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_985),
.A2(n_949),
.B1(n_891),
.B2(n_965),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_949),
.A2(n_736),
.B1(n_738),
.B2(n_744),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_SL g1062 ( 
.A(n_945),
.B(n_747),
.C(n_841),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_965),
.A2(n_738),
.B1(n_809),
.B2(n_846),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_946),
.B(n_1000),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_945),
.B(n_869),
.Y(n_1065)
);

OAI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_894),
.A2(n_776),
.B(n_875),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1008),
.A2(n_662),
.B(n_808),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_911),
.A2(n_791),
.B1(n_726),
.B2(n_844),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_901),
.Y(n_1069)
);

AO21x1_ASAP7_75t_L g1070 ( 
.A1(n_885),
.A2(n_844),
.B(n_682),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_901),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_916),
.A2(n_638),
.B(n_624),
.C(n_631),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_911),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_919),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_960),
.A2(n_622),
.B(n_662),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_935),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_904),
.B(n_379),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1003),
.A2(n_970),
.B1(n_1018),
.B2(n_1021),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_907),
.B(n_382),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1000),
.B(n_382),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_915),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_1011),
.A2(n_638),
.B(n_641),
.C(n_659),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_886),
.B(n_1038),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1033),
.B(n_387),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_966),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_935),
.Y(n_1086)
);

OA22x2_ASAP7_75t_L g1087 ( 
.A1(n_967),
.A2(n_392),
.B1(n_388),
.B2(n_387),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_975),
.A2(n_689),
.B(n_653),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_1031),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_1002),
.A2(n_722),
.B(n_626),
.C(n_689),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_944),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_R g1092 ( 
.A(n_984),
.B(n_726),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_944),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_914),
.Y(n_1094)
);

AO32x1_ASAP7_75t_L g1095 ( 
.A1(n_1018),
.A2(n_2),
.A3(n_4),
.B1(n_8),
.B2(n_12),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_966),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_882),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_986),
.A2(n_689),
.B(n_653),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1001),
.A2(n_1020),
.B(n_954),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1003),
.A2(n_722),
.B1(n_346),
.B2(n_342),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1034),
.B(n_626),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_895),
.Y(n_1102)
);

AND2x2_ASAP7_75t_SL g1103 ( 
.A(n_970),
.B(n_888),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_914),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_934),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_884),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_SL g1107 ( 
.A(n_982),
.B(n_936),
.C(n_938),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_924),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_928),
.B(n_340),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_977),
.B(n_626),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_925),
.A2(n_722),
.B1(n_639),
.B2(n_16),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_884),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_974),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_1113)
);

AO32x1_ASAP7_75t_L g1114 ( 
.A1(n_1035),
.A2(n_14),
.A3(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_961),
.A2(n_540),
.B(n_74),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_898),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_889),
.B(n_21),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1036),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_896),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_902),
.Y(n_1120)
);

CKINVDCx8_ASAP7_75t_R g1121 ( 
.A(n_921),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_892),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_937),
.B(n_24),
.Y(n_1123)
);

OAI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1014),
.A2(n_1016),
.B1(n_989),
.B2(n_936),
.C(n_938),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_903),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_929),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_988),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_SL g1128 ( 
.A(n_948),
.B(n_26),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_908),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_974),
.B(n_29),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_927),
.B(n_540),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_892),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_932),
.B(n_540),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_887),
.A2(n_29),
.B(n_31),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_999),
.A2(n_192),
.B(n_81),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1036),
.A2(n_79),
.B1(n_167),
.B2(n_157),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_948),
.B(n_31),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_888),
.B(n_76),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1024),
.A2(n_85),
.B(n_154),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1031),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_1140)
);

AOI222xp33_ASAP7_75t_L g1141 ( 
.A1(n_952),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.C1(n_55),
.C2(n_57),
.Y(n_1141)
);

CKINVDCx11_ASAP7_75t_R g1142 ( 
.A(n_921),
.Y(n_1142)
);

NOR2x1_ASAP7_75t_SL g1143 ( 
.A(n_896),
.B(n_90),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_952),
.B(n_46),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_929),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_928),
.B(n_57),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_941),
.B(n_58),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_956),
.A2(n_58),
.B(n_60),
.C(n_62),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_921),
.B(n_113),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_947),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_906),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1017),
.B(n_63),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_943),
.Y(n_1153)
);

OR2x6_ASAP7_75t_L g1154 ( 
.A(n_921),
.B(n_97),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_906),
.A2(n_98),
.B1(n_126),
.B2(n_134),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_959),
.B(n_187),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_997),
.A2(n_147),
.B1(n_148),
.B2(n_999),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_953),
.B(n_942),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_962),
.B(n_1025),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_909),
.A2(n_1025),
.B(n_1037),
.C(n_1041),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_900),
.B(n_899),
.C(n_893),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_930),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1023),
.B(n_896),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_954),
.A2(n_912),
.B(n_900),
.C(n_978),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_997),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_L g1166 ( 
.A(n_890),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1015),
.A2(n_1032),
.B1(n_1019),
.B2(n_1023),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_968),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1042),
.A2(n_950),
.B(n_964),
.C(n_1019),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_933),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_997),
.Y(n_1171)
);

AOI31xp67_ASAP7_75t_L g1172 ( 
.A1(n_1156),
.A2(n_1024),
.A3(n_1043),
.B(n_940),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1135),
.A2(n_960),
.B(n_926),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1057),
.A2(n_1029),
.B(n_1043),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1081),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1047),
.B(n_969),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1163),
.B(n_922),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1080),
.B(n_957),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1163),
.B(n_922),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1070),
.A2(n_1160),
.A3(n_1157),
.B(n_1060),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1054),
.B(n_990),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1121),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1067),
.A2(n_995),
.B(n_1027),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_L g1184 ( 
.A(n_1064),
.B(n_950),
.C(n_918),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1077),
.B(n_992),
.Y(n_1185)
);

AND3x4_ASAP7_75t_L g1186 ( 
.A(n_1086),
.B(n_993),
.C(n_976),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1060),
.A2(n_1020),
.B(n_1001),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1122),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1083),
.B(n_994),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1075),
.A2(n_1005),
.B(n_958),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1046),
.A2(n_939),
.B(n_1022),
.Y(n_1191)
);

AO21x1_ASAP7_75t_L g1192 ( 
.A1(n_1157),
.A2(n_1135),
.B(n_1151),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1063),
.A2(n_991),
.B1(n_1012),
.B2(n_987),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1169),
.A2(n_973),
.A3(n_979),
.B(n_1007),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1098),
.A2(n_981),
.B(n_983),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1063),
.A2(n_1009),
.B1(n_972),
.B2(n_998),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1155),
.A2(n_951),
.B(n_1006),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1071),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1051),
.B(n_996),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1142),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1072),
.A2(n_1040),
.B(n_1039),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1158),
.B(n_963),
.Y(n_1202)
);

AOI221x1_ASAP7_75t_L g1203 ( 
.A1(n_1078),
.A2(n_1028),
.B1(n_897),
.B2(n_923),
.C(n_980),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1045),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1094),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_SL g1206 ( 
.A(n_1141),
.B(n_951),
.C(n_1010),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1069),
.B(n_955),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1141),
.A2(n_923),
.B1(n_980),
.B2(n_1004),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1132),
.B(n_917),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1061),
.A2(n_1013),
.B(n_1028),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1123),
.B(n_1013),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1061),
.A2(n_1013),
.A3(n_1111),
.B(n_1088),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1085),
.B(n_1074),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1130),
.A2(n_1013),
.B1(n_1113),
.B2(n_1117),
.C(n_1124),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1066),
.A2(n_1059),
.B(n_1164),
.C(n_1065),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1161),
.A2(n_1062),
.B(n_1048),
.C(n_1167),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1126),
.B(n_1119),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1146),
.B(n_1144),
.Y(n_1218)
);

AOI221x1_ASAP7_75t_L g1219 ( 
.A1(n_1078),
.A2(n_1111),
.B1(n_1048),
.B2(n_1118),
.C(n_1155),
.Y(n_1219)
);

OAI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1134),
.A2(n_1084),
.B(n_1058),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1110),
.A2(n_1139),
.B(n_1101),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1145),
.B(n_1096),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1137),
.B(n_1126),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1049),
.B(n_1108),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1154),
.B(n_1055),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1082),
.A2(n_1152),
.B(n_1115),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1089),
.A2(n_1140),
.B(n_1107),
.C(n_1073),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1104),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1068),
.A2(n_1148),
.B(n_1153),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1147),
.B(n_1100),
.C(n_1136),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1079),
.B(n_1116),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1127),
.B(n_1105),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1044),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1168),
.B(n_1103),
.Y(n_1234)
);

NOR2x1_ASAP7_75t_L g1235 ( 
.A(n_1055),
.B(n_1112),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1131),
.A2(n_1133),
.B(n_1125),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1166),
.A2(n_1119),
.B1(n_1170),
.B2(n_1129),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1120),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1162),
.B(n_1109),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1150),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1143),
.A2(n_1114),
.A3(n_1095),
.B(n_1112),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1097),
.Y(n_1242)
);

AOI221x1_ASAP7_75t_L g1243 ( 
.A1(n_1095),
.A2(n_1114),
.B1(n_1171),
.B2(n_1165),
.C(n_1087),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1092),
.B(n_1171),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1165),
.B(n_1171),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1138),
.A2(n_1154),
.B(n_1119),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1093),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1154),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1044),
.B(n_1106),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1087),
.A2(n_1119),
.B(n_1128),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1050),
.A2(n_1106),
.B(n_1114),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1102),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1149),
.A2(n_1095),
.B(n_1106),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1076),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1047),
.B(n_913),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1122),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1075),
.A2(n_905),
.B(n_1099),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1054),
.B(n_913),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1070),
.A2(n_1160),
.A3(n_1157),
.B(n_1060),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1047),
.B(n_913),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1121),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1045),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1047),
.B(n_910),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1135),
.A2(n_1160),
.B(n_1090),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1066),
.A2(n_946),
.B(n_945),
.C(n_781),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1159),
.A2(n_910),
.B1(n_913),
.B2(n_945),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1054),
.B(n_913),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1155),
.A2(n_1135),
.B(n_1160),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1047),
.B(n_910),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1052),
.A2(n_945),
.B(n_751),
.C(n_786),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1057),
.A2(n_1067),
.B(n_1053),
.Y(n_1271)
);

AO22x2_ASAP7_75t_L g1272 ( 
.A1(n_1078),
.A2(n_946),
.B1(n_1063),
.B2(n_1060),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1135),
.A2(n_1160),
.B(n_1090),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1057),
.A2(n_1067),
.B(n_1053),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1135),
.A2(n_1160),
.B(n_1090),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1060),
.A2(n_910),
.B1(n_757),
.B2(n_913),
.Y(n_1276)
);

O2A1O1Ixp5_ASAP7_75t_L g1277 ( 
.A1(n_1052),
.A2(n_945),
.B(n_751),
.C(n_786),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1069),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1044),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1060),
.A2(n_910),
.B1(n_757),
.B2(n_913),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1138),
.B(n_945),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1075),
.A2(n_905),
.B(n_1099),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1075),
.A2(n_905),
.B(n_1099),
.Y(n_1283)
);

AND2x6_ASAP7_75t_L g1284 ( 
.A(n_1165),
.B(n_921),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1054),
.B(n_591),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1075),
.A2(n_905),
.B(n_1099),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1160),
.A2(n_946),
.B(n_1060),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1121),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1081),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1163),
.B(n_884),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1080),
.B(n_742),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1047),
.B(n_910),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1047),
.B(n_786),
.C(n_781),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1075),
.A2(n_905),
.B(n_1099),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1056),
.Y(n_1295)
);

INVx3_ASAP7_75t_SL g1296 ( 
.A(n_1091),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1159),
.A2(n_910),
.B1(n_913),
.B2(n_945),
.Y(n_1297)
);

AO32x2_ASAP7_75t_L g1298 ( 
.A1(n_1060),
.A2(n_1078),
.A3(n_1111),
.B1(n_1018),
.B2(n_1157),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1080),
.B(n_742),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1075),
.A2(n_905),
.B(n_1099),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1054),
.B(n_913),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1060),
.A2(n_910),
.B1(n_757),
.B2(n_913),
.Y(n_1302)
);

NOR2x1_ASAP7_75t_SL g1303 ( 
.A(n_1154),
.B(n_1119),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_1094),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1080),
.B(n_742),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1278),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1257),
.A2(n_1283),
.B(n_1282),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1203),
.A2(n_1287),
.B(n_1226),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1285),
.B(n_1278),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1265),
.A2(n_1293),
.B(n_1215),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1208),
.A2(n_1268),
.B1(n_1293),
.B2(n_1230),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1270),
.A2(n_1277),
.B(n_1287),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1286),
.A2(n_1300),
.B(n_1294),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1218),
.B(n_1291),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1246),
.B(n_1217),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1209),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1216),
.B(n_1266),
.Y(n_1318)
);

BUFx4f_ASAP7_75t_SL g1319 ( 
.A(n_1188),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_1242),
.B(n_1247),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1227),
.A2(n_1302),
.B(n_1280),
.C(n_1276),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1175),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1193),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_1191),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1221),
.A2(n_1174),
.B(n_1183),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1281),
.A2(n_1192),
.B(n_1197),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1297),
.B(n_1281),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1230),
.A2(n_1220),
.B(n_1214),
.C(n_1208),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1219),
.A2(n_1187),
.B(n_1184),
.Y(n_1330)
);

BUFx5_ASAP7_75t_L g1331 ( 
.A(n_1284),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1201),
.A2(n_1210),
.B(n_1187),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1184),
.A2(n_1229),
.B(n_1302),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1210),
.A2(n_1251),
.B(n_1236),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1194),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1194),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1264),
.A2(n_1273),
.B(n_1275),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1276),
.A2(n_1280),
.B(n_1206),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1272),
.B(n_1220),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1255),
.A2(n_1260),
.B1(n_1258),
.B2(n_1267),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1295),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1289),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1238),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1299),
.A2(n_1305),
.B1(n_1231),
.B2(n_1234),
.C(n_1301),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1253),
.A2(n_1193),
.B(n_1196),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1243),
.A2(n_1237),
.A3(n_1303),
.B(n_1172),
.Y(n_1346)
);

OR2x6_ASAP7_75t_L g1347 ( 
.A(n_1225),
.B(n_1248),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1292),
.B(n_1176),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1264),
.A2(n_1275),
.B(n_1273),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1181),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1173),
.A2(n_1199),
.B(n_1202),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1225),
.A2(n_1224),
.B1(n_1200),
.B2(n_1239),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1250),
.A2(n_1245),
.B(n_1211),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1186),
.A2(n_1225),
.B1(n_1189),
.B2(n_1223),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1173),
.A2(n_1178),
.B(n_1185),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1207),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1212),
.A2(n_1180),
.A3(n_1259),
.B(n_1194),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1180),
.A2(n_1259),
.B(n_1240),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1235),
.A2(n_1249),
.B(n_1244),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1180),
.A2(n_1259),
.B(n_1212),
.Y(n_1360)
);

AO32x2_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1241),
.A3(n_1212),
.B1(n_1233),
.B2(n_1279),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1304),
.Y(n_1362)
);

OR2x6_ASAP7_75t_L g1363 ( 
.A(n_1217),
.B(n_1200),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1298),
.A2(n_1241),
.B(n_1205),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1198),
.B(n_1232),
.Y(n_1365)
);

OAI221xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1298),
.A2(n_1254),
.B1(n_1204),
.B2(n_1262),
.C(n_1252),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1241),
.A2(n_1290),
.B(n_1213),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1182),
.Y(n_1368)
);

INVxp33_ASAP7_75t_L g1369 ( 
.A(n_1182),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1290),
.A2(n_1209),
.B(n_1182),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1261),
.A2(n_1288),
.B(n_1256),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1261),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1261),
.B(n_1288),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1288),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1296),
.A2(n_1293),
.B(n_946),
.C(n_1277),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1268),
.A2(n_1274),
.B(n_1271),
.Y(n_1376)
);

AO32x2_ASAP7_75t_L g1377 ( 
.A1(n_1276),
.A2(n_1060),
.A3(n_1078),
.B1(n_1302),
.B2(n_1280),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1246),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1182),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1182),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1218),
.B(n_1291),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1218),
.B(n_1291),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1208),
.A2(n_1268),
.B1(n_1293),
.B2(n_1230),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1182),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1293),
.A2(n_946),
.B1(n_1272),
.B2(n_1141),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1386)
);

OR2x6_ASAP7_75t_L g1387 ( 
.A(n_1246),
.B(n_1225),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1388)
);

AO32x2_ASAP7_75t_L g1389 ( 
.A1(n_1276),
.A2(n_1060),
.A3(n_1078),
.B1(n_1302),
.B2(n_1280),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1265),
.A2(n_946),
.B(n_1216),
.C(n_1293),
.Y(n_1390)
);

OAI221xp5_ASAP7_75t_L g1391 ( 
.A1(n_1293),
.A2(n_949),
.B1(n_1265),
.B2(n_946),
.C(n_913),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1203),
.A2(n_1287),
.B(n_1226),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1228),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1265),
.A2(n_946),
.B(n_1216),
.C(n_1293),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1194),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_SL g1396 ( 
.A1(n_1265),
.A2(n_946),
.B(n_1216),
.C(n_1227),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1293),
.A2(n_946),
.B1(n_1272),
.B2(n_1141),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1257),
.A2(n_1283),
.B(n_1282),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1303),
.A2(n_1246),
.B(n_1192),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1175),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1175),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1209),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1175),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1268),
.A2(n_1274),
.B(n_1271),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1218),
.B(n_1291),
.Y(n_1406)
);

AOI21xp33_ASAP7_75t_L g1407 ( 
.A1(n_1293),
.A2(n_1230),
.B(n_1265),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1200),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1182),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1281),
.A2(n_946),
.B1(n_552),
.B2(n_553),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1188),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1257),
.A2(n_1283),
.B(n_1282),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1218),
.B(n_1291),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1416)
);

BUFx10_ASAP7_75t_L g1417 ( 
.A(n_1182),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1182),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1222),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1246),
.B(n_1225),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1175),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1208),
.A2(n_1281),
.B1(n_1293),
.B2(n_1219),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1218),
.B(n_1291),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1200),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1175),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1265),
.B(n_1060),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1203),
.A2(n_1287),
.B(n_1226),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1268),
.A2(n_1274),
.B(n_1271),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1293),
.B(n_609),
.C(n_949),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1315),
.B(n_1381),
.Y(n_1431)
);

NOR2xp67_ASAP7_75t_L g1432 ( 
.A(n_1350),
.B(n_1309),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1347),
.B(n_1363),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1382),
.B(n_1406),
.Y(n_1434)
);

BUFx4f_ASAP7_75t_SL g1435 ( 
.A(n_1408),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1371),
.B(n_1306),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1323),
.B(n_1340),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1415),
.B(n_1423),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1356),
.B(n_1419),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1337),
.A2(n_1312),
.B(n_1326),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1430),
.A2(n_1394),
.B(n_1390),
.C(n_1329),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1385),
.A2(n_1397),
.B1(n_1366),
.B2(n_1323),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1312),
.A2(n_1326),
.B(n_1349),
.Y(n_1443)
);

AOI21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1339),
.A2(n_1327),
.B(n_1386),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1339),
.A2(n_1327),
.B(n_1386),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1340),
.B(n_1310),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1407),
.A2(n_1383),
.B(n_1311),
.C(n_1333),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1347),
.B(n_1363),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1385),
.A2(n_1397),
.B1(n_1366),
.B2(n_1391),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1376),
.A2(n_1429),
.B(n_1405),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1348),
.B(n_1355),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1391),
.A2(n_1422),
.B1(n_1410),
.B2(n_1411),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1362),
.B(n_1306),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1355),
.B(n_1371),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1390),
.B(n_1394),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1422),
.A2(n_1410),
.B1(n_1411),
.B2(n_1399),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1313),
.B(n_1328),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1380),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1376),
.A2(n_1429),
.B(n_1405),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_SL g1460 ( 
.A1(n_1388),
.A2(n_1427),
.B(n_1426),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1319),
.Y(n_1461)
);

BUFx8_ASAP7_75t_L g1462 ( 
.A(n_1424),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1375),
.A2(n_1420),
.B(n_1387),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1416),
.A2(n_1426),
.B1(n_1412),
.B2(n_1321),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1318),
.B(n_1330),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1321),
.A2(n_1344),
.B1(n_1318),
.B2(n_1333),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1319),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1325),
.A2(n_1324),
.B(n_1334),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1413),
.B(n_1344),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1396),
.A2(n_1354),
.B(n_1352),
.C(n_1393),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1393),
.B(n_1367),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1417),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1342),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1474)
);

AOI21x1_ASAP7_75t_SL g1475 ( 
.A1(n_1335),
.A2(n_1395),
.B(n_1336),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1341),
.B(n_1343),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1354),
.A2(n_1428),
.B1(n_1308),
.B2(n_1392),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1368),
.Y(n_1478)
);

O2A1O1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1400),
.A2(n_1368),
.B(n_1365),
.C(n_1372),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1332),
.A2(n_1370),
.B(n_1320),
.C(n_1359),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1351),
.B(n_1338),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1387),
.B(n_1420),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1338),
.B(n_1316),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1387),
.B(n_1420),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1374),
.A2(n_1370),
.B(n_1401),
.C(n_1421),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1402),
.A2(n_1425),
.B(n_1404),
.C(n_1373),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1307),
.A2(n_1398),
.B(n_1314),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1317),
.B(n_1403),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1369),
.B(n_1418),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1379),
.A2(n_1384),
.B(n_1409),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1345),
.B(n_1358),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1345),
.B(n_1360),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1417),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1357),
.B(n_1353),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1361),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1331),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1364),
.B(n_1357),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1361),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1331),
.A2(n_1377),
.B(n_1389),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1346),
.B(n_1331),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1414),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1346),
.B(n_1377),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1346),
.B(n_1323),
.Y(n_1503)
);

O2A1O1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1396),
.A2(n_946),
.B(n_1265),
.C(n_1227),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1378),
.A2(n_1246),
.B(n_1265),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1315),
.B(n_1381),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1347),
.B(n_1363),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1315),
.B(n_1381),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1323),
.B(n_1340),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1315),
.B(n_1381),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1385),
.A2(n_1208),
.B1(n_1397),
.B2(n_1268),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1430),
.A2(n_945),
.B(n_1281),
.C(n_1293),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1376),
.A2(n_1429),
.B(n_1405),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1413),
.Y(n_1514)
);

BUFx8_ASAP7_75t_L g1515 ( 
.A(n_1408),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1322),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1315),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1315),
.B(n_1381),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1385),
.A2(n_1208),
.B1(n_1397),
.B2(n_1268),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1396),
.A2(n_946),
.B(n_1265),
.C(n_1227),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1323),
.B(n_1340),
.Y(n_1521)
);

O2A1O1Ixp5_ASAP7_75t_L g1522 ( 
.A1(n_1310),
.A2(n_1192),
.B(n_1287),
.C(n_1407),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1306),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_SL g1524 ( 
.A(n_1387),
.B(n_1420),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1376),
.A2(n_1429),
.B(n_1405),
.Y(n_1525)
);

OAI31xp33_ASAP7_75t_L g1526 ( 
.A1(n_1430),
.A2(n_1293),
.A3(n_945),
.B(n_609),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1376),
.A2(n_1429),
.B(n_1405),
.Y(n_1527)
);

OAI31xp33_ASAP7_75t_L g1528 ( 
.A1(n_1430),
.A2(n_1293),
.A3(n_945),
.B(n_609),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1323),
.B(n_1340),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1396),
.A2(n_946),
.B(n_1265),
.C(n_1227),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1315),
.B(n_1381),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1450),
.A2(n_1525),
.B(n_1513),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1454),
.B(n_1451),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1436),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1487),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1450),
.A2(n_1525),
.B(n_1513),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1459),
.B(n_1527),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1463),
.B(n_1482),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1462),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1471),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1481),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1477),
.B(n_1499),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1432),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1473),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1523),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1484),
.B(n_1505),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1511),
.A2(n_1519),
.B1(n_1449),
.B2(n_1442),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1501),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1492),
.B(n_1494),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1453),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1483),
.B(n_1474),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1492),
.B(n_1502),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1497),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1483),
.B(n_1500),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_R g1556 ( 
.A(n_1446),
.B(n_1433),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1491),
.A2(n_1522),
.B(n_1447),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1500),
.B(n_1480),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1437),
.B(n_1509),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1437),
.B(n_1509),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1495),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1529),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1498),
.B(n_1521),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1468),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1443),
.B(n_1440),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1455),
.A2(n_1446),
.B(n_1465),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1496),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1441),
.A2(n_1530),
.B(n_1504),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1440),
.B(n_1465),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1468),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1448),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1511),
.A2(n_1519),
.B1(n_1449),
.B2(n_1464),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1439),
.B(n_1476),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1512),
.A2(n_1486),
.B(n_1466),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1431),
.B(n_1434),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1448),
.B(n_1507),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1438),
.B(n_1531),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1506),
.B(n_1508),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1485),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1570),
.B(n_1466),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1570),
.B(n_1456),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1535),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1456),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1547),
.A2(n_1528),
.B1(n_1526),
.B2(n_1442),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1517),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1575),
.A2(n_1469),
.B1(n_1452),
.B2(n_1464),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1569),
.B(n_1470),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1518),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1534),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1533),
.B(n_1510),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1540),
.B(n_1478),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1561),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1540),
.Y(n_1595)
);

AOI31xp33_ASAP7_75t_L g1596 ( 
.A1(n_1547),
.A2(n_1461),
.A3(n_1467),
.B(n_1457),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1548),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1520),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1541),
.B(n_1475),
.Y(n_1599)
);

OAI322xp33_ASAP7_75t_L g1600 ( 
.A1(n_1569),
.A2(n_1479),
.A3(n_1490),
.B1(n_1445),
.B2(n_1444),
.C1(n_1514),
.C2(n_1460),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1565),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1488),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1533),
.B(n_1489),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1555),
.B(n_1532),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1458),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1592),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1585),
.A2(n_1573),
.B1(n_1575),
.B2(n_1560),
.C(n_1562),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_SL g1608 ( 
.A(n_1588),
.B(n_1539),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1593),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1601),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1593),
.Y(n_1611)
);

OAI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1585),
.A2(n_1573),
.B1(n_1575),
.B2(n_1560),
.C(n_1562),
.Y(n_1612)
);

OAI33xp33_ASAP7_75t_L g1613 ( 
.A1(n_1599),
.A2(n_1566),
.A3(n_1554),
.B1(n_1549),
.B2(n_1559),
.B3(n_1580),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1593),
.Y(n_1614)
);

NAND2xp33_ASAP7_75t_R g1615 ( 
.A(n_1588),
.B(n_1575),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1594),
.Y(n_1616)
);

AOI33xp33_ASAP7_75t_L g1617 ( 
.A1(n_1587),
.A2(n_1550),
.A3(n_1558),
.B1(n_1563),
.B2(n_1551),
.B3(n_1544),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

OAI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1598),
.A2(n_1559),
.B(n_1543),
.C(n_1557),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1600),
.A2(n_1536),
.B1(n_1532),
.B2(n_1546),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1594),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_R g1622 ( 
.A(n_1592),
.B(n_1539),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1594),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1603),
.B(n_1545),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1595),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_R g1626 ( 
.A(n_1592),
.B(n_1539),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1605),
.A2(n_1571),
.B(n_1564),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1584),
.A2(n_1546),
.B1(n_1536),
.B2(n_1532),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1586),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1595),
.Y(n_1630)
);

BUFx12f_ASAP7_75t_L g1631 ( 
.A(n_1586),
.Y(n_1631)
);

AOI31xp33_ASAP7_75t_L g1632 ( 
.A1(n_1602),
.A2(n_1556),
.A3(n_1572),
.B(n_1577),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1602),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1538),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1584),
.A2(n_1546),
.B1(n_1536),
.B2(n_1538),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1600),
.A2(n_1537),
.B(n_1546),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1590),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1581),
.A2(n_1557),
.B1(n_1552),
.B2(n_1538),
.Y(n_1638)
);

AOI322xp5_ASAP7_75t_L g1639 ( 
.A1(n_1582),
.A2(n_1579),
.A3(n_1578),
.B1(n_1576),
.B2(n_1563),
.C1(n_1558),
.C2(n_1574),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1599),
.B(n_1552),
.C(n_1558),
.Y(n_1640)
);

AO21x2_ASAP7_75t_L g1641 ( 
.A1(n_1583),
.A2(n_1571),
.B(n_1564),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1610),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1622),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1641),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1641),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1611),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1622),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1614),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1616),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1621),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1623),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1610),
.Y(n_1654)
);

INVx4_ASAP7_75t_SL g1655 ( 
.A(n_1634),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1625),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1636),
.A2(n_1537),
.B(n_1596),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1610),
.Y(n_1658)
);

INVx4_ASAP7_75t_SL g1659 ( 
.A(n_1634),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1630),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1606),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1632),
.B(n_1568),
.Y(n_1662)
);

INVx4_ASAP7_75t_SL g1663 ( 
.A(n_1634),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1618),
.B(n_1637),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1653),
.B(n_1633),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1645),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1643),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1642),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1642),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1653),
.B(n_1610),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1655),
.B(n_1610),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1654),
.B(n_1628),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1568),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1654),
.B(n_1604),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1647),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1645),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1654),
.B(n_1604),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1644),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1639),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1658),
.B(n_1655),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1644),
.B(n_1631),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1655),
.B(n_1635),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1660),
.B(n_1617),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1646),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1649),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1655),
.B(n_1627),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1648),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1643),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

CKINVDCx16_ASAP7_75t_R g1693 ( 
.A(n_1648),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1655),
.B(n_1638),
.Y(n_1694)
);

AND4x1_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1608),
.C(n_1617),
.D(n_1620),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1659),
.B(n_1638),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1664),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1660),
.B(n_1591),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1664),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1646),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1650),
.B(n_1651),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_SL g1702 ( 
.A(n_1662),
.B(n_1613),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1659),
.B(n_1597),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1681),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1693),
.B(n_1435),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1669),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1669),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1670),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_SL g1709 ( 
.A1(n_1690),
.A2(n_1699),
.B(n_1684),
.C(n_1686),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1683),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1681),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1699),
.B(n_1651),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1670),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1674),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1693),
.B(n_1643),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1678),
.Y(n_1718)
);

AND2x4_ASAP7_75t_SL g1719 ( 
.A(n_1673),
.B(n_1661),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1695),
.B(n_1657),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1688),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1702),
.A2(n_1685),
.B1(n_1696),
.B2(n_1694),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1688),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1701),
.Y(n_1724)
);

OAI21xp33_ASAP7_75t_L g1725 ( 
.A1(n_1702),
.A2(n_1657),
.B(n_1620),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1685),
.B(n_1659),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1695),
.B(n_1659),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.B(n_1659),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1665),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1673),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.B(n_1663),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1681),
.B(n_1663),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1683),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1697),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1701),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1697),
.B(n_1665),
.Y(n_1736)
);

BUFx12f_ASAP7_75t_L g1737 ( 
.A(n_1697),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1663),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1684),
.B(n_1589),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1698),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1682),
.B(n_1624),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1686),
.B(n_1652),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1712),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1716),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1719),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1704),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1712),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1726),
.B(n_1683),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1707),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1737),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1671),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1711),
.B(n_1682),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1704),
.B(n_1675),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1729),
.B(n_1672),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1737),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1708),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1731),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1713),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1728),
.B(n_1671),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1720),
.A2(n_1694),
.B1(n_1696),
.B2(n_1675),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1734),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1722),
.A2(n_1596),
.B1(n_1612),
.B2(n_1607),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1734),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1710),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1710),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1720),
.A2(n_1725),
.B1(n_1727),
.B2(n_1728),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1731),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1732),
.B(n_1671),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1758),
.B(n_1709),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1764),
.A2(n_1727),
.B1(n_1615),
.B2(n_1732),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1746),
.Y(n_1773)
);

NAND2x1p5_ASAP7_75t_L g1774 ( 
.A(n_1751),
.B(n_1738),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1748),
.B(n_1705),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1764),
.A2(n_1709),
.B(n_1738),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1745),
.A2(n_1615),
.B1(n_1741),
.B2(n_1736),
.Y(n_1777)
);

AOI21xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1768),
.A2(n_1676),
.B(n_1733),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1762),
.A2(n_1753),
.B(n_1756),
.C(n_1751),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1744),
.A2(n_1742),
.B(n_1719),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1758),
.B(n_1733),
.Y(n_1781)
);

OAI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1756),
.A2(n_1675),
.B(n_1694),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1754),
.B(n_1742),
.C(n_1735),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1745),
.A2(n_1739),
.B1(n_1666),
.B2(n_1696),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1746),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1769),
.A2(n_1666),
.B1(n_1640),
.B2(n_1676),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1746),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1755),
.A2(n_1769),
.B1(n_1666),
.B2(n_1747),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1763),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1748),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1752),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1752),
.B(n_1724),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1761),
.B(n_1770),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1775),
.B(n_1761),
.Y(n_1794)
);

NOR3xp33_ASAP7_75t_L g1795 ( 
.A(n_1779),
.B(n_1747),
.C(n_1743),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1773),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1790),
.B(n_1770),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1793),
.B(n_1755),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1785),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1774),
.Y(n_1800)
);

NOR2x1_ASAP7_75t_L g1801 ( 
.A(n_1776),
.B(n_1763),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1791),
.B(n_1743),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1774),
.B(n_1782),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1780),
.B(n_1766),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1787),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1789),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1771),
.B(n_1763),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1788),
.B(n_1765),
.Y(n_1808)
);

OAI211xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1801),
.A2(n_1776),
.B(n_1772),
.C(n_1781),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1795),
.A2(n_1788),
.B(n_1778),
.C(n_1786),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1803),
.A2(n_1783),
.B1(n_1777),
.B2(n_1784),
.C(n_1792),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1797),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1804),
.A2(n_1767),
.B1(n_1676),
.B2(n_1730),
.Y(n_1813)
);

AOI211xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1807),
.A2(n_1730),
.B(n_1765),
.C(n_1767),
.Y(n_1814)
);

OAI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1808),
.A2(n_1765),
.B(n_1767),
.C(n_1757),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_SL g1816 ( 
.A(n_1808),
.B(n_1676),
.C(n_1626),
.Y(n_1816)
);

NOR3xp33_ASAP7_75t_L g1817 ( 
.A(n_1800),
.B(n_1802),
.C(n_1798),
.Y(n_1817)
);

OAI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1794),
.A2(n_1730),
.B1(n_1691),
.B2(n_1668),
.Y(n_1818)
);

OAI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1796),
.A2(n_1691),
.B1(n_1668),
.B2(n_1740),
.Y(n_1819)
);

XOR2x2_ASAP7_75t_L g1820 ( 
.A(n_1806),
.B(n_1462),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1815),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1809),
.A2(n_1805),
.B(n_1799),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_1817),
.B(n_1750),
.C(n_1749),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1812),
.B(n_1816),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1820),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1814),
.B(n_1749),
.Y(n_1826)
);

OAI322xp33_ASAP7_75t_L g1827 ( 
.A1(n_1810),
.A2(n_1760),
.A3(n_1759),
.B1(n_1757),
.B2(n_1750),
.C1(n_1691),
.C2(n_1723),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1826),
.Y(n_1828)
);

NAND2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1824),
.B(n_1515),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1822),
.A2(n_1811),
.B(n_1813),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1827),
.B(n_1818),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1821),
.B(n_1819),
.Y(n_1832)
);

NAND2x1_ASAP7_75t_L g1833 ( 
.A(n_1823),
.B(n_1759),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1825),
.B(n_1760),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1826),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_R g1836 ( 
.A(n_1828),
.B(n_1515),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1829),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1830),
.A2(n_1717),
.B(n_1715),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1834),
.Y(n_1839)
);

OAI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1833),
.A2(n_1668),
.B1(n_1718),
.B2(n_1721),
.Y(n_1840)
);

AO22x1_ASAP7_75t_L g1841 ( 
.A1(n_1832),
.A2(n_1673),
.B1(n_1668),
.B2(n_1472),
.Y(n_1841)
);

NAND4xp75_ASAP7_75t_L g1842 ( 
.A(n_1839),
.B(n_1835),
.C(n_1831),
.D(n_1689),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1840),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1837),
.B(n_1668),
.Y(n_1844)
);

NAND4xp75_ASAP7_75t_L g1845 ( 
.A(n_1838),
.B(n_1689),
.C(n_1703),
.D(n_1677),
.Y(n_1845)
);

XNOR2xp5_ASAP7_75t_L g1846 ( 
.A(n_1842),
.B(n_1841),
.Y(n_1846)
);

NOR3xp33_ASAP7_75t_L g1847 ( 
.A(n_1843),
.B(n_1836),
.C(n_1493),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1846),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1847),
.A2(n_1844),
.B1(n_1845),
.B2(n_1673),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1848),
.Y(n_1850)
);

INVx3_ASAP7_75t_SL g1851 ( 
.A(n_1849),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1850),
.Y(n_1852)
);

CKINVDCx20_ASAP7_75t_R g1853 ( 
.A(n_1851),
.Y(n_1853)
);

AO22x2_ASAP7_75t_L g1854 ( 
.A1(n_1852),
.A2(n_1692),
.B1(n_1687),
.B2(n_1667),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1853),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1855),
.A2(n_1673),
.B1(n_1672),
.B2(n_1687),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1856),
.B(n_1854),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1679),
.B(n_1667),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1858),
.A2(n_1689),
.B1(n_1703),
.B2(n_1680),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1667),
.B1(n_1700),
.B2(n_1679),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1679),
.B(n_1700),
.C(n_1667),
.Y(n_1861)
);


endmodule