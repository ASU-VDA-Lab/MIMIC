module real_jpeg_33143_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_0),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_0),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_2),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

CKINVDCx11_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_67),
.B1(n_69),
.B2(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_73),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_3),
.A2(n_73),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_3),
.A2(n_73),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_6),
.A2(n_29),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_29),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

AOI22x1_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_29),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_6),
.B(n_328),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g400 ( 
.A1(n_6),
.A2(n_401),
.A3(n_408),
.B1(n_411),
.B2(n_417),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_6),
.B(n_149),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_7),
.Y(n_407)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_7),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_8),
.Y(n_59)
);

AO22x2_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_59),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22x1_ASAP7_75t_R g156 ( 
.A1(n_8),
.A2(n_59),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_8),
.A2(n_59),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_9),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_9),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_12),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_13),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_13),
.A2(n_107),
.B1(n_253),
.B2(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_13),
.A2(n_253),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_13),
.A2(n_253),
.B1(n_429),
.B2(n_432),
.Y(n_428)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_289),
.B(n_542),
.Y(n_17)
);

O2A1O1Ixp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_268),
.B(n_284),
.C(n_285),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_227),
.B(n_267),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_21),
.B(n_536),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_199),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_22),
.B(n_199),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_145),
.C(n_163),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_23),
.A2(n_145),
.B1(n_146),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_23),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_64),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_24),
.B(n_65),
.C(n_111),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_24),
.A2(n_202),
.B1(n_225),
.B2(n_226),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_55),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_25),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_35),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_26),
.A2(n_35),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_26),
.B(n_62),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_28),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_29),
.B(n_63),
.Y(n_305)
);

AOI32xp33_ASAP7_75t_L g318 ( 
.A1(n_29),
.A2(n_319),
.A3(n_322),
.B1(n_326),
.B2(n_327),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_29),
.B(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_29),
.B(n_113),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_29),
.B(n_303),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_30),
.Y(n_362)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_35),
.B(n_56),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_35),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_35),
.Y(n_276)
);

NOR2x1p5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_41),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_43),
.Y(n_208)
);

AO22x2_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_44),
.Y(n_348)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_45),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_45),
.B(n_249),
.Y(n_375)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_48),
.Y(n_223)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_50),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_55),
.A2(n_204),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_55),
.B(n_248),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_57),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_111),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_74),
.B(n_101),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_74),
.B(n_218),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_74),
.A2(n_218),
.B(n_280),
.Y(n_279)
);

AO21x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_82),
.B(n_90),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_82),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_84),
.Y(n_345)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_97),
.B2(n_100),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_101),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2x1p5_ASAP7_75t_SL g244 ( 
.A(n_102),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_103),
.Y(n_280)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NAND2x1_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_110),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_111),
.A2(n_213),
.B1(n_214),
.B2(n_224),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_111),
.B(n_214),
.C(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_111),
.A2(n_224),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g491 ( 
.A(n_111),
.B(n_374),
.C(n_377),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_124),
.B(n_139),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_139),
.Y(n_154)
);

NAND2x1p5_ASAP7_75t_L g195 ( 
.A(n_112),
.B(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_112),
.B(n_189),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_112),
.B(n_332),
.Y(n_385)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_125),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_122),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_118),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_118),
.Y(n_431)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_120),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_124),
.B(n_332),
.Y(n_331)
);

NAND2x1_ASAP7_75t_L g424 ( 
.A(n_124),
.B(n_139),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.B1(n_134),
.B2(n_136),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_128),
.Y(n_321)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_136),
.Y(n_421)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21x1_ASAP7_75t_SL g259 ( 
.A1(n_146),
.A2(n_147),
.B(n_153),
.Y(n_259)
);

NAND2x1p5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_149),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_149),
.B(n_311),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_151),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_152),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_154),
.B(n_331),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_155),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_155),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_155),
.B(n_231),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_159),
.Y(n_419)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_162),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_163),
.B(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_185),
.B(n_196),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_164),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_164),
.B(n_197),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_164),
.B(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_164),
.A2(n_186),
.B1(n_318),
.B2(n_392),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_164),
.A2(n_186),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_169),
.B(n_178),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_169),
.A2(n_301),
.B(n_367),
.Y(n_484)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_170),
.B(n_179),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_170),
.B(n_428),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_174),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_174),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_175),
.Y(n_368)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_176),
.Y(n_450)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_185),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_187),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_194),
.B(n_195),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_195),
.B(n_331),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_195),
.B(n_424),
.Y(n_485)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_196),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_196),
.B(n_539),
.Y(n_542)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_200),
.Y(n_283)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_202),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_212),
.Y(n_202)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_209),
.B(n_210),
.Y(n_203)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_210),
.B(n_257),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_211),
.B(n_375),
.Y(n_482)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_216),
.B(n_310),
.Y(n_473)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_282),
.C(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_264),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_228),
.B(n_264),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_258),
.C(n_260),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_229),
.B(n_518),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_243),
.C(n_246),
.Y(n_229)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_230),
.Y(n_514)
);

XOR2x2_ASAP7_75t_SL g478 ( 
.A(n_232),
.B(n_479),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

AND2x4_ASAP7_75t_SL g426 ( 
.A(n_233),
.B(n_427),
.Y(n_426)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_237),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_238),
.A2(n_364),
.B(n_367),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_238),
.B(n_445),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_244),
.B(n_247),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_245),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_259),
.B(n_262),
.Y(n_518)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_268),
.B(n_285),
.Y(n_534)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_281),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_281),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_275),
.C(n_277),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_278),
.B(n_507),
.C(n_508),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_279),
.B(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_287),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_287),
.B(n_288),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_533),
.B(n_537),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_524),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_467),
.B(n_523),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_380),
.B(n_466),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_337),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_295),
.B(n_337),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_316),
.C(n_330),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_296),
.B(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_308),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_299),
.Y(n_448)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_301),
.B(n_427),
.Y(n_442)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_339)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_330),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_373),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_372),
.Y(n_338)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_339),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_340),
.B(n_495),
.C(n_496),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_340),
.B(n_495),
.C(n_496),
.Y(n_528)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_363),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_342),
.B(n_363),
.Y(n_476)
);

OAI31xp33_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_346),
.A3(n_349),
.B(n_353),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_358),
.B(n_362),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx2_ASAP7_75t_R g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_373),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_389),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_395),
.B(n_465),
.Y(n_380)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_393),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_382),
.B(n_393),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.C(n_390),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_383),
.A2(n_384),
.B1(n_387),
.B2(n_388),
.Y(n_463)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_424),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_463),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_458),
.B(n_464),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_438),
.B(n_457),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_425),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_398),
.B(n_425),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_422),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_399),
.A2(n_400),
.B1(n_422),
.B2(n_423),
.Y(n_455)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx4f_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_435),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_426),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_460),
.C(n_461),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_453),
.B(n_456),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_443),
.B(n_452),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_442),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_449),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NOR2x1_ASAP7_75t_L g456 ( 
.A(n_454),
.B(n_455),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_462),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_500),
.C(n_516),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_493),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_469),
.B(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_486),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_470),
.B(n_486),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_477),
.Y(n_470)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_471),
.Y(n_502)
);

MAJx2_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_474),
.C(n_476),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_473),
.A2(n_474),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_473),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_475),
.Y(n_490)
);

XNOR2x1_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_488),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.Y(n_477)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_478),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_482),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

XOR2x2_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_485),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_491),
.C(n_492),
.Y(n_486)
);

XNOR2x1_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_499),
.Y(n_498)
);

XOR2x1_ASAP7_75t_SL g499 ( 
.A(n_491),
.B(n_492),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_498),
.Y(n_493)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_529),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_505),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_501),
.B(n_505),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.C(n_504),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_509),
.Y(n_505)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_513),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_510),
.Y(n_521)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_513),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_519),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_519),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_521),
.C(n_522),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_531),
.C(n_532),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_529),
.C(n_530),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_535),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_538),
.A2(n_540),
.B(n_541),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_539),
.Y(n_538)
);


endmodule