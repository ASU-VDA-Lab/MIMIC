module fake_jpeg_20742_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_26),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_17),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_19),
.B1(n_25),
.B2(n_35),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_64),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_30),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_36),
.Y(n_74)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_73),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_67),
.B(n_98),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_25),
.B1(n_41),
.B2(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_68),
.A2(n_77),
.B1(n_104),
.B2(n_71),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_36),
.CI(n_39),
.CON(n_73),
.SN(n_73)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_80),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_41),
.B1(n_44),
.B2(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_84),
.B1(n_85),
.B2(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_41),
.B1(n_22),
.B2(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_40),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_21),
.B(n_20),
.C(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_99),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_38),
.B1(n_39),
.B2(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_39),
.B(n_40),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_37),
.B(n_43),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_40),
.C(n_37),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_93),
.C(n_37),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_40),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_59),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_43),
.Y(n_129)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_40),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_43),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_22),
.B1(n_39),
.B2(n_26),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_38),
.A3(n_63),
.B1(n_58),
.B2(n_50),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_43),
.C(n_16),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_108),
.A2(n_125),
.B(n_78),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_95),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_55),
.B1(n_54),
.B2(n_63),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_123),
.B1(n_67),
.B2(n_98),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_118),
.B(n_131),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_37),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_65),
.A2(n_33),
.B1(n_43),
.B2(n_37),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_103),
.B1(n_99),
.B2(n_86),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_33),
.B1(n_43),
.B2(n_28),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_73),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_27),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_133),
.A2(n_72),
.B1(n_88),
.B2(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_75),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_18),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_92),
.C(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_147),
.C(n_158),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_143),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_145),
.B1(n_152),
.B2(n_127),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_82),
.B1(n_81),
.B2(n_34),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_116),
.B1(n_128),
.B2(n_108),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_83),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_166),
.B1(n_117),
.B2(n_132),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_95),
.B1(n_102),
.B2(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_87),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_87),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_31),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_78),
.C(n_70),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_32),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_79),
.B(n_18),
.C(n_16),
.D(n_31),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_126),
.B(n_18),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_79),
.B1(n_29),
.B2(n_28),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_126),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_89),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_125),
.B1(n_123),
.B2(n_113),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_185),
.B1(n_162),
.B2(n_148),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_122),
.B1(n_127),
.B2(n_131),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_178),
.B1(n_189),
.B2(n_152),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_111),
.B1(n_124),
.B2(n_114),
.Y(n_178)
);

AOI221xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_160),
.B1(n_156),
.B2(n_143),
.C(n_162),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_184),
.Y(n_213)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_132),
.B1(n_130),
.B2(n_117),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_106),
.C(n_130),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_147),
.C(n_138),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_171),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_194),
.B(n_161),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_155),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_31),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_159),
.B1(n_139),
.B2(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_201),
.B(n_203),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_209),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_221),
.C(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_207),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_156),
.B(n_146),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_187),
.B(n_170),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_167),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_210),
.A2(n_219),
.B(n_223),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_164),
.B1(n_149),
.B2(n_34),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_149),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_16),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_194),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_191),
.B1(n_170),
.B2(n_196),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_1),
.B(n_2),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_197),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_34),
.C(n_32),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_172),
.B(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_185),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_187),
.A2(n_180),
.B(n_182),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_231),
.C(n_221),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_232),
.B(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_176),
.C(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_217),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_243),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_194),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_245),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_206),
.B1(n_204),
.B2(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_200),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_168),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_208),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_257),
.C(n_263),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_204),
.B(n_216),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_262),
.B(n_244),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_202),
.B1(n_223),
.B2(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_224),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_168),
.B1(n_218),
.B2(n_219),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_175),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_234),
.B1(n_241),
.B2(n_230),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_184),
.B1(n_175),
.B2(n_11),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_226),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_8),
.B(n_13),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_34),
.C(n_8),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_274),
.B1(n_259),
.B2(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_232),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_231),
.C(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_249),
.C(n_263),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_230),
.B(n_238),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_6),
.B(n_13),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_260),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_270),
.C(n_271),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_274),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_229),
.B(n_250),
.C(n_249),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_289),
.C(n_266),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_251),
.B(n_229),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_265),
.B(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_7),
.C(n_12),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_6),
.C(n_8),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_267),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_282),
.B1(n_286),
.B2(n_4),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_287),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_297),
.C(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_278),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_271),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_299),
.B(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_2),
.B(n_3),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_294),
.C(n_299),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_291),
.B(n_292),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_4),
.B(n_2),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_311),
.B(n_3),
.Y(n_312)
);


endmodule