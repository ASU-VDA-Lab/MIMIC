module real_jpeg_18850_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g58 ( 
.A(n_0),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_508),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_1),
.B(n_509),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_2),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_2),
.B(n_134),
.Y(n_223)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_3),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_3),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_175),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_3),
.B(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_4),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_5),
.B(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_5),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_5),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_5),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_5),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_5),
.B(n_255),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_6),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_6),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_7),
.B(n_69),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_7),
.B(n_180),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_7),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_7),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_7),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_7),
.B(n_421),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_8),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_8),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_8),
.B(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_8),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_8),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_8),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_8),
.B(n_469),
.Y(n_468)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_9),
.Y(n_257)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_9),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_10),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g308 ( 
.A(n_10),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g371 ( 
.A(n_10),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_10),
.B(n_115),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g410 ( 
.A(n_10),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_10),
.B(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_11),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_12),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_12),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_12),
.Y(n_401)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_14),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_15),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_15),
.B(n_132),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_15),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_15),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_15),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_15),
.B(n_444),
.Y(n_443)
);

AND2x2_ASAP7_75t_SL g455 ( 
.A(n_15),
.B(n_456),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_16),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_16),
.Y(n_423)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_17),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_163),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_162),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_140),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_23),
.B(n_140),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_72),
.C(n_102),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_24),
.B(n_72),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_51),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_25),
.B(n_52),
.C(n_64),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_26),
.B(n_49),
.C(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.C(n_35),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_28),
.B(n_35),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_29),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_32),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_32),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_33),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_33),
.Y(n_125)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_34),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_35),
.B(n_189),
.C(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_35),
.A2(n_36),
.B1(n_189),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_46),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_46),
.A2(n_50),
.B1(n_135),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_46),
.A2(n_50),
.B1(n_193),
.B2(n_194),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_50),
.B(n_129),
.C(n_135),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_50),
.B(n_188),
.C(n_193),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_64),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_53),
.B(n_56),
.C(n_60),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_56),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_56),
.A2(n_63),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_56),
.B(n_92),
.C(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_56),
.A2(n_63),
.B1(n_207),
.B2(n_208),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_57),
.B(n_136),
.Y(n_135)
);

NAND2x1_ASAP7_75t_L g151 ( 
.A(n_57),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_59),
.B(n_113),
.Y(n_331)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.C(n_68),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_60),
.B(n_114),
.C(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_62),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_65),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_77),
.C(n_83),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_75),
.B1(n_83),
.B2(n_84),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_65),
.B(n_308),
.C(n_311),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_65),
.A2(n_75),
.B1(n_308),
.B2(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_67),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_86),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_73),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_76),
.B(n_86),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_131),
.C(n_133),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_83),
.A2(n_84),
.B1(n_133),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_84),
.B(n_223),
.Y(n_428)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_85),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_85),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_96),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_90),
.Y(n_310)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_92),
.A2(n_122),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_97),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_103),
.B(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_123),
.C(n_128),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_104),
.B(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_120),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_105),
.B(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_107),
.B(n_120),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.C(n_116),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_114),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_133),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_174),
.B(n_178),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_133),
.A2(n_171),
.B1(n_174),
.B2(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_133),
.B(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_134),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_135),
.Y(n_197)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_150),
.A2(n_151),
.B1(n_226),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_221),
.C(n_226),
.Y(n_220)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_154),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx11_ASAP7_75t_SL g161 ( 
.A(n_156),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_500),
.B(n_504),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_241),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_230),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_166),
.B(n_230),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_R g166 ( 
.A(n_167),
.B(n_198),
.C(n_201),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_167),
.B(n_199),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_186),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_168),
.B(n_187),
.C(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_183),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_169),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_171),
.B(n_420),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_172),
.B(n_183),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_174),
.B(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_174),
.A2(n_205),
.B1(n_305),
.B2(n_306),
.Y(n_364)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_177),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_182),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_182),
.A2(n_334),
.B1(n_486),
.B2(n_487),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_201),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_215),
.C(n_219),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_202),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.C(n_212),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_203),
.B(n_206),
.Y(n_323)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_211),
.Y(n_342)
);

XOR2x1_ASAP7_75t_L g322 ( 
.A(n_212),
.B(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_289)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.C(n_224),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_223),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_239),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_233),
.B(n_235),
.C(n_239),
.Y(n_503)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_387),
.Y(n_241)
);

A2O1A1O1Ixp25_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_324),
.B(n_377),
.C(n_378),
.D(n_386),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_244),
.B(n_379),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_294),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_245),
.B(n_294),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_287),
.Y(n_245)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_246),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_271),
.C(n_283),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.C(n_261),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_249),
.B(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_251),
.A2(n_252),
.B1(n_261),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_252),
.A2(n_253),
.B(n_258),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.C(n_266),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_263),
.Y(n_302)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_266),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_267),
.B(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_283),
.B1(n_284),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.C(n_280),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_276),
.Y(n_317)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_279),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_281),
.B(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_290),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_299),
.C(n_321),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_296),
.B1(n_322),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_316),
.C(n_318),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_307),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_301),
.B(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_303),
.A2(n_304),
.B1(n_307),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_311),
.B(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_349),
.B(n_376),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_346),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_346),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.C(n_343),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_343),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.C(n_333),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_332),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.C(n_340),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_335),
.A2(n_340),
.B1(n_341),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_335),
.Y(n_488)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_352),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.C(n_360),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_353),
.A2(n_354),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_357),
.B(n_360),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_365),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_361),
.B(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_364),
.B(n_365),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.C(n_374),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_366),
.A2(n_367),
.B1(n_374),
.B2(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2x1_ASAP7_75t_L g436 ( 
.A(n_371),
.B(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_374),
.Y(n_438)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_384),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.C(n_383),
.Y(n_380)
);

NAND4xp25_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.C(n_390),
.D(n_391),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_494),
.B(n_499),
.Y(n_391)
);

AOI21x1_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_482),
.B(n_493),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_439),
.B(n_481),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_424),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_395),
.B(n_424),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_409),
.C(n_418),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_396),
.B(n_478),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_408),
.C(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_408),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_409),
.A2(n_418),
.B1(n_419),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_415),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_415),
.Y(n_452)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_433),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_425),
.B(n_434),
.C(n_436),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_429),
.C(n_431),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_427)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_428),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_430),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_475),
.B(n_480),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_462),
.B(n_474),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_451),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_442),
.B(n_451),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_447),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_447),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_455),
.C(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_467),
.B(n_473),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_466),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_476),
.B(n_477),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_492),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_492),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_490),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_489),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_489),
.C(n_490),
.Y(n_495)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_496),
.Y(n_499)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_500),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

NOR2x1_ASAP7_75t_R g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_503),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);


endmodule