module fake_jpeg_762_n_65 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_20),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_27),
.C(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_38),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_1),
.C(n_2),
.Y(n_38)
);

XNOR2x2_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_19),
.Y(n_39)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_3),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_18),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_11),
.B(n_17),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_52),
.B(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_44),
.B1(n_6),
.B2(n_7),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_4),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_12),
.C(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_47),
.B(n_8),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_60),
.C(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_59),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OAI221xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_54),
.B1(n_15),
.B2(n_16),
.C(n_9),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_7),
.Y(n_65)
);


endmodule