module real_jpeg_23747_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_1),
.A2(n_82),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_1),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_93),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_93),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_93),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_85),
.B(n_87),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_77),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_26),
.C(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_67),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_41),
.B1(n_186),
.B2(n_193),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_71),
.Y(n_176)
);

INVx8_ASAP7_75t_SL g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_8),
.A2(n_69),
.B1(n_92),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_56),
.Y(n_141)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_114),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_52),
.B1(n_94),
.B2(n_95),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_22),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_24),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_24),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_24),
.B(n_89),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_25),
.B(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_31),
.A2(n_32),
.B1(n_62),
.B2(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_62),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_32),
.A2(n_63),
.A3(n_65),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_32),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_35),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_35),
.A2(n_146),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_35),
.A2(n_145),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_35),
.A2(n_144),
.B1(n_145),
.B2(n_166),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_48),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_41),
.A2(n_48),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_41),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_41),
.A2(n_183),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_42),
.B(n_49),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_42),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_51),
.Y(n_178)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.C(n_73),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_70),
.B(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_68),
.B1(n_72),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_67),
.B1(n_128),
.B2(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_65),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_79),
.B(n_88),
.C(n_109),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g137 ( 
.A(n_64),
.B(n_89),
.CON(n_137),
.SN(n_137)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_78),
.C(n_102),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_84),
.B2(n_90),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_77),
.B1(n_91),
.B2(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_86),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_89),
.B(n_194),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_115),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_120),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_209),
.B(n_213),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_160),
.B(n_208),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_147),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_134),
.B(n_147),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.C(n_143),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_135),
.B(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_142),
.B(n_143),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_155),
.C(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_159),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_154),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_203),
.B(n_207),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_179),
.B(n_202),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_189),
.B(n_201),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_188),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_196),
.B(n_200),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);


endmodule