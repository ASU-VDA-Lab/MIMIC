module fake_jpeg_23546_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_0),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_50),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_25),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_22),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_35),
.B1(n_30),
.B2(n_24),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_35),
.B1(n_24),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_59),
.B1(n_71),
.B2(n_27),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g101 ( 
.A(n_55),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_35),
.B1(n_18),
.B2(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_16),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_30),
.B1(n_23),
.B2(n_20),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_19),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_19),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_58),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_107),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_26),
.B1(n_31),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_98),
.B1(n_52),
.B2(n_66),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_22),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_72),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_26),
.B1(n_27),
.B2(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_104),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_49),
.B(n_22),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_14),
.B(n_11),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_28),
.B(n_3),
.C(n_4),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_51),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_117),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_129),
.B1(n_95),
.B2(n_93),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_122),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_80),
.B(n_84),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_55),
.B1(n_50),
.B2(n_52),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_131),
.B1(n_95),
.B2(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_136),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_63),
.C(n_42),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_88),
.B(n_81),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_128),
.C(n_137),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_42),
.C(n_63),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_66),
.B1(n_48),
.B2(n_56),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_1),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_108),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_48),
.B1(n_56),
.B2(n_28),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_135),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_2),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_85),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_157),
.CI(n_120),
.CON(n_170),
.SN(n_170)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_146),
.B(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_114),
.B(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_157),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_83),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_91),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_161),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_133),
.B1(n_115),
.B2(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_172),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_159),
.C(n_142),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_176),
.B1(n_160),
.B2(n_113),
.Y(n_190)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_150),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_114),
.B1(n_109),
.B2(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_147),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_169),
.A2(n_151),
.B1(n_152),
.B2(n_145),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_167),
.B1(n_181),
.B2(n_171),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_194),
.Y(n_208)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_123),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_140),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.C(n_191),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_175),
.A3(n_179),
.B1(n_177),
.B2(n_170),
.Y(n_189)
);

AOI321xp33_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_166),
.A3(n_148),
.B1(n_178),
.B2(n_168),
.C(n_118),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_189),
.A3(n_195),
.B1(n_196),
.B2(n_191),
.C1(n_187),
.C2(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_154),
.C(n_156),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_196),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_138),
.B1(n_134),
.B2(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_164),
.B1(n_177),
.B2(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_123),
.B1(n_184),
.B2(n_183),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_180),
.C(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_209),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_89),
.B(n_83),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_118),
.B(n_89),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_91),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_208),
.B(n_204),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_201),
.B(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_216),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_143),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_64),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_206),
.C(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_117),
.C(n_74),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_227),
.B(n_220),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_225),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_64),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_2),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_224),
.B(n_222),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_219),
.C(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_231),
.C(n_6),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_211),
.C(n_218),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_212),
.B1(n_7),
.B2(n_8),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_234),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_225),
.Y(n_234)
);

AOI31xp33_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_7),
.A3(n_9),
.B(n_10),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_235),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_10),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_240),
.Y(n_242)
);


endmodule