module fake_ariane_2133_n_1757 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1757);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1757;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_53),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_33),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_108),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_28),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_27),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_49),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_34),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_21),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_111),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_49),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_20),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_115),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_92),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_76),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_39),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_59),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_128),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_36),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_130),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_109),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_39),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_41),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_83),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_6),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_35),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_25),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_72),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_117),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_19),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_37),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_46),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_123),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_85),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_12),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_112),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_77),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_31),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_132),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_81),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_71),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_9),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_7),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_35),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_103),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_129),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_17),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_48),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_4),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_2),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_97),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_60),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_59),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_101),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_9),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_32),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_65),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_27),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_126),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_43),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_38),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_125),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_30),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_70),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_138),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_12),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_96),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_94),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_154),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_17),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_98),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_119),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_42),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_116),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_54),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_7),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_102),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_16),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_38),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_139),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_24),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_3),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_88),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_41),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_46),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_69),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_24),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_152),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_21),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_75),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_121),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_16),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_144),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_118),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_30),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_4),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_53),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_99),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_106),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_84),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_37),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_50),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_13),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_48),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_11),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_14),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_34),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_104),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_0),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_89),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_124),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_40),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_20),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_10),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_54),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_148),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_100),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_180),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_0),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_210),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_210),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_200),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_205),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_169),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_174),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_203),
.B(n_1),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_210),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_210),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_218),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_210),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_210),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_210),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_173),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_173),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_159),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_166),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_203),
.B(n_3),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_159),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_169),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_171),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_161),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_161),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_192),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_212),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_162),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_231),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_169),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_182),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_182),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_242),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_275),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_238),
.B(n_5),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_169),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_244),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_178),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_250),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_178),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_306),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_268),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_230),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_285),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_181),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_238),
.B(n_5),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_169),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_181),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_158),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_186),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_160),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_188),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_198),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_189),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_174),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_191),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_202),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_196),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_186),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_217),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_217),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_222),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_245),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_179),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_201),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

CKINVDCx6p67_ASAP7_75t_R g391 ( 
.A(n_363),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_245),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_336),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_333),
.B(n_263),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_263),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_276),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_321),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_321),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_213),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_340),
.B(n_276),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_326),
.A2(n_286),
.B(n_283),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_337),
.A2(n_286),
.B(n_283),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_351),
.B(n_230),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_340),
.B(n_213),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_312),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_337),
.A2(n_303),
.B(n_183),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_342),
.B(n_303),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_342),
.B(n_190),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_319),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_316),
.B(n_299),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_344),
.Y(n_438)
);

NAND2x1_ASAP7_75t_L g439 ( 
.A(n_344),
.B(n_190),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_316),
.B(n_179),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_365),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_348),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_430),
.A2(n_363),
.B1(n_319),
.B2(n_335),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_436),
.A2(n_324),
.B1(n_354),
.B2(n_366),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_383),
.C(n_382),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_414),
.B(n_371),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_361),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_314),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_414),
.B(n_373),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_372),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

NOR2x1p5_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_443),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_436),
.A2(n_314),
.B1(n_300),
.B2(n_322),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

BUFx6f_ASAP7_75t_SL g480 ( 
.A(n_391),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_422),
.A2(n_385),
.B1(n_384),
.B2(n_383),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_375),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_451),
.B(n_377),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_447),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_391),
.B(n_313),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

BUFx4f_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_419),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_447),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_451),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_SL g494 ( 
.A(n_394),
.B(n_409),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_422),
.A2(n_385),
.B1(n_384),
.B2(n_382),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_447),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_419),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_396),
.B(n_265),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_447),
.B(n_387),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_451),
.B(n_369),
.Y(n_504)
);

BUFx6f_ASAP7_75t_SL g505 ( 
.A(n_431),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_157),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_451),
.B(n_353),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_439),
.B(n_348),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_394),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_394),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_322),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_447),
.B(n_163),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_451),
.B(n_431),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_451),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_431),
.B(n_379),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_395),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_396),
.B(n_198),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_450),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_376),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_422),
.A2(n_413),
.B1(n_408),
.B2(n_396),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_396),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_434),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_434),
.B(n_386),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_409),
.B(n_198),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_422),
.A2(n_253),
.B1(n_288),
.B2(n_226),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_442),
.C(n_429),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_429),
.B(n_198),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_434),
.B(n_352),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_410),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_429),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_374),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_434),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_446),
.B(n_352),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_446),
.B(n_374),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_410),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_439),
.A2(n_272),
.B1(n_292),
.B2(n_183),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

BUFx4f_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_455),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_442),
.B(n_208),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_399),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_395),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_417),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_443),
.A2(n_298),
.B1(n_204),
.B2(n_290),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_417),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_446),
.B(n_378),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_455),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_415),
.B(n_378),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_417),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_442),
.A2(n_318),
.B1(n_320),
.B2(n_327),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_455),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_388),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_417),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_446),
.B(n_215),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_415),
.B(n_164),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_418),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_446),
.B(n_170),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_444),
.B(n_194),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_441),
.B(n_219),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_388),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_443),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_455),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_441),
.B(n_444),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_388),
.B(n_259),
.C(n_224),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_441),
.B(n_176),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_423),
.B(n_164),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_454),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_390),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_454),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_399),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_454),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_441),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_454),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_418),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_408),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_408),
.A2(n_278),
.B1(n_209),
.B2(n_233),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_456),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_413),
.A2(n_253),
.B1(n_235),
.B2(n_288),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_456),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_399),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_418),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_423),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_456),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_SL g606 ( 
.A(n_511),
.B(n_541),
.C(n_513),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_459),
.A2(n_425),
.B1(n_454),
.B2(n_438),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_469),
.B(n_393),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_491),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_470),
.B(n_444),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_475),
.B(n_423),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_459),
.A2(n_500),
.B1(n_510),
.B2(n_573),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_570),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_570),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_560),
.A2(n_413),
.B1(n_408),
.B2(n_454),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_522),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_604),
.A2(n_420),
.B(n_397),
.C(n_390),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_469),
.B(n_418),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_462),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_469),
.B(n_393),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_546),
.B(n_445),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_558),
.B(n_334),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_525),
.B(n_445),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_491),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_508),
.B(n_418),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_508),
.B(n_527),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_462),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_508),
.B(n_390),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_530),
.B(n_445),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_527),
.B(n_392),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_527),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_449),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_581),
.B(n_392),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_573),
.B(n_449),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_466),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_500),
.A2(n_425),
.B1(n_454),
.B2(n_438),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_579),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_587),
.B(n_449),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_558),
.B(n_397),
.C(n_392),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_579),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_587),
.B(n_452),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_550),
.B(n_452),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_465),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_563),
.B(n_452),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_528),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_581),
.B(n_397),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_463),
.B(n_420),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_581),
.B(n_420),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_534),
.B(n_424),
.C(n_421),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_560),
.A2(n_413),
.B1(n_408),
.B2(n_456),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_589),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_583),
.A2(n_424),
.B(n_421),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_466),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_465),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_589),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_542),
.B(n_421),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_575),
.A2(n_398),
.B1(n_400),
.B2(n_411),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_480),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_542),
.B(n_424),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_457),
.B(n_456),
.C(n_400),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_565),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_521),
.B(n_523),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_580),
.A2(n_398),
.B1(n_411),
.B2(n_401),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_565),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_565),
.B(n_448),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_490),
.B(n_456),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_560),
.A2(n_413),
.B1(n_408),
.B2(n_456),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_490),
.B(n_399),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_559),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_559),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_565),
.B(n_448),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_597),
.B(n_401),
.C(n_448),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_490),
.B(n_399),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_580),
.B(n_498),
.Y(n_678)
);

INVxp33_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_561),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_561),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_554),
.B(n_399),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_500),
.A2(n_448),
.B1(n_453),
.B2(n_260),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_488),
.B(n_476),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_560),
.A2(n_413),
.B1(n_453),
.B2(n_248),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_538),
.B(n_453),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_514),
.B(n_453),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_471),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_585),
.B(n_399),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_476),
.B(n_338),
.Y(n_691)
);

NAND2x1_ASAP7_75t_L g692 ( 
.A(n_500),
.B(n_403),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_554),
.B(n_399),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_566),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_505),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_566),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_510),
.B(n_399),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_557),
.B(n_416),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_473),
.B(n_416),
.Y(n_699)
);

BUFx6f_ASAP7_75t_SL g700 ( 
.A(n_510),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_494),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_471),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_599),
.A2(n_500),
.B1(n_533),
.B2(n_597),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_567),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_484),
.B(n_416),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_584),
.A2(n_206),
.B1(n_224),
.B2(n_226),
.C(n_235),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_557),
.B(n_416),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_500),
.A2(n_247),
.B1(n_258),
.B2(n_232),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_567),
.B(n_416),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_557),
.B(n_416),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_571),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_480),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_483),
.Y(n_714)
);

BUFx6f_ASAP7_75t_SL g715 ( 
.A(n_510),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_461),
.B(n_403),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_557),
.B(n_416),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_483),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_556),
.B(n_577),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_572),
.A2(n_309),
.B(n_280),
.C(n_297),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_596),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_475),
.B(n_341),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_574),
.B(n_416),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_574),
.B(n_416),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_595),
.B(n_194),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_SL g727 ( 
.A(n_532),
.B(n_220),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_467),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_535),
.B(n_343),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_595),
.B(n_404),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_603),
.B(n_404),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_603),
.B(n_407),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_500),
.B(n_407),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_467),
.B(n_412),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_467),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_489),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_467),
.B(n_345),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_507),
.B(n_227),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_482),
.B(n_412),
.Y(n_739)
);

BUFx12f_ASAP7_75t_SL g740 ( 
.A(n_552),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_591),
.B(n_412),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_495),
.B(n_206),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_493),
.B(n_274),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_489),
.B(n_274),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_591),
.B(n_405),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_499),
.B(n_501),
.Y(n_746)
);

BUFx8_ASAP7_75t_L g747 ( 
.A(n_505),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_591),
.B(n_405),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_591),
.B(n_405),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_499),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_505),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_584),
.B(n_350),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_501),
.B(n_277),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_502),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_L g755 ( 
.A1(n_552),
.A2(n_277),
.B1(n_280),
.B2(n_282),
.C(n_309),
.Y(n_755)
);

AOI22x1_ASAP7_75t_L g756 ( 
.A1(n_598),
.A2(n_282),
.B1(n_297),
.B2(n_437),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_504),
.B(n_228),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_526),
.B(n_356),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_576),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_503),
.A2(n_258),
.B1(n_214),
.B2(n_211),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_502),
.B(n_234),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_461),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_598),
.B(n_236),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_509),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_509),
.B(n_239),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_512),
.B(n_240),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_512),
.B(n_243),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_591),
.B(n_405),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_517),
.B(n_246),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_517),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_531),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_601),
.B(n_405),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_531),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_601),
.B(n_405),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_539),
.B(n_359),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_539),
.B(n_249),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_551),
.B(n_252),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_493),
.B(n_519),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_699),
.A2(n_528),
.B(n_518),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_610),
.B(n_551),
.Y(n_780)
);

NAND2x1_ASAP7_75t_L g781 ( 
.A(n_633),
.B(n_553),
.Y(n_781)
);

BUFx4f_ASAP7_75t_L g782 ( 
.A(n_662),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_706),
.A2(n_486),
.B(n_553),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_612),
.A2(n_588),
.B(n_592),
.C(n_594),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_683),
.B(n_601),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_649),
.A2(n_592),
.B(n_588),
.Y(n_786)
);

O2A1O1Ixp5_ASAP7_75t_L g787 ( 
.A1(n_651),
.A2(n_598),
.B(n_497),
.C(n_537),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_672),
.A2(n_594),
.B(n_468),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_672),
.A2(n_468),
.B(n_464),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_624),
.B(n_362),
.Y(n_790)
);

OR2x2_ASAP7_75t_SL g791 ( 
.A(n_722),
.B(n_606),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_656),
.A2(n_472),
.B(n_464),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_677),
.A2(n_474),
.B(n_472),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_610),
.B(n_519),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_622),
.B(n_460),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_622),
.B(n_460),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_633),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_611),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_683),
.B(n_601),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_607),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_682),
.A2(n_478),
.B(n_477),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_693),
.A2(n_479),
.B(n_478),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_690),
.A2(n_485),
.B(n_481),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_607),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_614),
.A2(n_605),
.B(n_602),
.C(n_485),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_608),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_667),
.A2(n_605),
.B(n_602),
.C(n_487),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_670),
.A2(n_492),
.B(n_487),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_669),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_678),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_660),
.A2(n_549),
.B(n_547),
.C(n_548),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_670),
.A2(n_496),
.B(n_492),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_637),
.B(n_460),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_641),
.B(n_645),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_666),
.A2(n_524),
.B(n_516),
.C(n_586),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_652),
.A2(n_516),
.B(n_496),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_683),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_497),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_608),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_626),
.B(n_497),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_658),
.B(n_364),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_647),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_621),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_775),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_703),
.A2(n_537),
.B1(n_600),
.B2(n_578),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_621),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_636),
.A2(n_524),
.B(n_520),
.Y(n_827)
);

BUFx12f_ASAP7_75t_L g828 ( 
.A(n_713),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_675),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_666),
.B(n_537),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_665),
.B(n_578),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_752),
.B(n_691),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_629),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_683),
.B(n_601),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_764),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_668),
.B(n_578),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_758),
.B(n_164),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_600),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_704),
.B(n_600),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_629),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_686),
.A2(n_248),
.B1(n_296),
.B2(n_576),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_762),
.B(n_520),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_751),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_673),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_704),
.B(n_590),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_636),
.A2(n_650),
.B(n_623),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_618),
.B(n_248),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_L g849 ( 
.A(n_723),
.B(n_254),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_661),
.B(n_529),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_681),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_704),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_676),
.A2(n_529),
.B(n_586),
.C(n_582),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_650),
.A2(n_548),
.B(n_582),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_743),
.B(n_536),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_743),
.B(n_609),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_662),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_694),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_704),
.B(n_590),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_747),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_687),
.A2(n_547),
.B(n_569),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_710),
.A2(n_545),
.B(n_569),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_724),
.A2(n_545),
.B(n_564),
.Y(n_863)
);

OAI321xp33_ASAP7_75t_L g864 ( 
.A1(n_707),
.A2(n_432),
.A3(n_437),
.B1(n_435),
.B2(n_296),
.C(n_433),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_685),
.B(n_536),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_743),
.B(n_540),
.Y(n_866)
);

NAND2x1_ASAP7_75t_L g867 ( 
.A(n_674),
.B(n_540),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_696),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_618),
.B(n_296),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_705),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_738),
.B(n_544),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_725),
.A2(n_549),
.B(n_564),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_646),
.A2(n_562),
.B(n_555),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_740),
.Y(n_874)
);

CKINVDCx10_ASAP7_75t_R g875 ( 
.A(n_700),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_720),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_738),
.B(n_544),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_734),
.B(n_590),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_747),
.Y(n_879)
);

BUFx8_ASAP7_75t_L g880 ( 
.A(n_700),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_688),
.B(n_555),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_701),
.B(n_562),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_688),
.B(n_257),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_741),
.A2(n_515),
.B(n_506),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_619),
.A2(n_632),
.B(n_630),
.C(n_615),
.Y(n_885)
);

BUFx12f_ASAP7_75t_L g886 ( 
.A(n_737),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_735),
.B(n_628),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_741),
.A2(n_576),
.B(n_437),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_648),
.A2(n_177),
.B(n_184),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_625),
.A2(n_172),
.B(n_185),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_261),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_751),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_638),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_631),
.A2(n_167),
.B(n_168),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_698),
.A2(n_165),
.B(n_187),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_628),
.B(n_266),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_698),
.A2(n_711),
.B(n_708),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_708),
.A2(n_711),
.B(n_746),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_728),
.B(n_269),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_620),
.A2(n_576),
.B(n_437),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_620),
.A2(n_627),
.B(n_634),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_712),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_679),
.B(n_271),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_627),
.A2(n_281),
.B(n_195),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_718),
.A2(n_284),
.B(n_197),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_630),
.A2(n_287),
.B(n_199),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_717),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_744),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_635),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_697),
.B(n_405),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_662),
.B(n_432),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_739),
.A2(n_435),
.B(n_432),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_632),
.A2(n_616),
.B(n_655),
.C(n_659),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_613),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_SL g916 ( 
.A1(n_653),
.A2(n_432),
.B(n_435),
.C(n_10),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_640),
.B(n_289),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_642),
.A2(n_308),
.B1(n_307),
.B2(n_301),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_638),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_613),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_644),
.B(n_435),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_763),
.B(n_576),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_727),
.B(n_193),
.C(n_207),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_664),
.A2(n_697),
.B(n_757),
.C(n_721),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_730),
.A2(n_273),
.B(n_223),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_731),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_732),
.A2(n_279),
.B(n_225),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_291),
.B(n_216),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_757),
.B(n_576),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_736),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_716),
.A2(n_576),
.B(n_405),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_613),
.A2(n_293),
.B1(n_221),
.B2(n_229),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_679),
.B(n_6),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_695),
.B(n_237),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_674),
.A2(n_302),
.B(n_241),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_695),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_617),
.B(n_251),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_729),
.Y(n_939)
);

AOI21xp33_ASAP7_75t_L g940 ( 
.A1(n_742),
.A2(n_709),
.B(n_733),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_750),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_684),
.B(n_405),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_639),
.A2(n_433),
.B(n_428),
.C(n_427),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_680),
.A2(n_305),
.B(n_264),
.Y(n_944)
);

OAI21xp33_ASAP7_75t_L g945 ( 
.A1(n_761),
.A2(n_255),
.B(n_256),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_778),
.Y(n_946)
);

O2A1O1Ixp5_ASAP7_75t_L g947 ( 
.A1(n_765),
.A2(n_433),
.B(n_428),
.C(n_427),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_680),
.B(n_433),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_635),
.B(n_433),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_643),
.B(n_433),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_654),
.B(n_267),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_745),
.A2(n_310),
.B(n_311),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_745),
.A2(n_749),
.B(n_748),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_748),
.A2(n_433),
.B(n_428),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_657),
.A2(n_270),
.B(n_294),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_657),
.A2(n_433),
.B(n_428),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_643),
.B(n_433),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_689),
.B(n_427),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_671),
.B(n_11),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_689),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_702),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_766),
.B(n_13),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_702),
.B(n_427),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_749),
.A2(n_774),
.B(n_772),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_857),
.B(n_715),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_814),
.A2(n_778),
.B1(n_755),
.B2(n_776),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_880),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_876),
.B(n_715),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_881),
.A2(n_778),
.B(n_770),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_821),
.B(n_767),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_892),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_856),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_838),
.A2(n_777),
.B1(n_769),
.B2(n_773),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_780),
.A2(n_756),
.B1(n_760),
.B2(n_692),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_844),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_835),
.Y(n_976)
);

OAI22x1_ASAP7_75t_L g977 ( 
.A1(n_934),
.A2(n_754),
.B1(n_719),
.B2(n_714),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_790),
.B(n_774),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_809),
.B(n_754),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_829),
.B(n_714),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_798),
.B(n_759),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_800),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_891),
.A2(n_768),
.B(n_15),
.C(n_18),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_939),
.B(n_759),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_837),
.B(n_759),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_927),
.B(n_726),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_920),
.B(n_428),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_877),
.A2(n_304),
.B(n_194),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_934),
.B(n_14),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_832),
.B(n_426),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_782),
.B(n_726),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_828),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_810),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_794),
.A2(n_304),
.B(n_194),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_904),
.A2(n_726),
.B1(n_428),
.B2(n_427),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_822),
.B(n_15),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_848),
.B(n_22),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_850),
.A2(n_304),
.B(n_194),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_925),
.A2(n_304),
.B1(n_426),
.B2(n_427),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_925),
.A2(n_428),
.B(n_427),
.C(n_426),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_920),
.B(n_428),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_844),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_SL g1003 ( 
.A1(n_886),
.A2(n_726),
.B1(n_304),
.B2(n_427),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_882),
.B(n_726),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_883),
.A2(n_23),
.B(n_25),
.C(n_26),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_892),
.B(n_427),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_882),
.B(n_23),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_824),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_845),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_782),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_804),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_887),
.A2(n_428),
.B1(n_426),
.B2(n_36),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_896),
.A2(n_28),
.B(n_29),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_851),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_865),
.B(n_29),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_874),
.B(n_42),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_865),
.B(n_887),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_L g1018 ( 
.A1(n_884),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_896),
.A2(n_44),
.B(n_45),
.C(n_47),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_935),
.B(n_426),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_858),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_797),
.B(n_426),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_795),
.A2(n_426),
.B(n_93),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_797),
.B(n_426),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_915),
.B(n_426),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_817),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_796),
.A2(n_87),
.B(n_151),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_817),
.B(n_50),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_805),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_817),
.B(n_51),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_922),
.A2(n_95),
.B(n_150),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_852),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_852),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_847),
.A2(n_839),
.B(n_830),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_868),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_918),
.B(n_52),
.C(n_55),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_946),
.B(n_57),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_886),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_946),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_779),
.A2(n_64),
.B(n_73),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_817),
.B(n_78),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_805),
.A2(n_80),
.B1(n_82),
.B2(n_86),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_852),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_869),
.B(n_105),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_885),
.A2(n_107),
.B(n_113),
.C(n_120),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_909),
.B(n_122),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_828),
.B(n_153),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_923),
.B(n_131),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_898),
.A2(n_135),
.B(n_142),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_962),
.A2(n_146),
.B(n_901),
.C(n_914),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_910),
.B(n_933),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_910),
.B(n_843),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_852),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_873),
.A2(n_792),
.B(n_861),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_783),
.A2(n_803),
.B(n_816),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_818),
.B(n_813),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_959),
.A2(n_866),
.B1(n_855),
.B2(n_815),
.Y(n_1057)
);

INVx6_ASAP7_75t_L g1058 ( 
.A(n_903),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_870),
.B(n_902),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_908),
.B(n_931),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_937),
.B(n_903),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_849),
.A2(n_842),
.B1(n_938),
.B2(n_941),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_912),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_937),
.B(n_806),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_819),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_819),
.B(n_823),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_842),
.A2(n_823),
.B1(n_961),
.B2(n_960),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_789),
.A2(n_802),
.B(n_812),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_826),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_912),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_899),
.B(n_917),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_860),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_912),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_784),
.A2(n_924),
.B(n_811),
.C(n_807),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_929),
.A2(n_815),
.B(n_940),
.C(n_945),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_905),
.B(n_889),
.C(n_907),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_916),
.A2(n_853),
.B(n_831),
.C(n_836),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_793),
.A2(n_801),
.B(n_808),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_833),
.B(n_841),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_955),
.A2(n_930),
.B(n_953),
.C(n_964),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_893),
.Y(n_1081)
);

OA22x2_ASAP7_75t_L g1082 ( 
.A1(n_879),
.A2(n_951),
.B1(n_919),
.B2(n_961),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_919),
.B(n_960),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_791),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_878),
.A2(n_785),
.B(n_834),
.C(n_799),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_820),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_897),
.A2(n_862),
.B(n_863),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_864),
.B(n_894),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_872),
.A2(n_788),
.B(n_786),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_853),
.A2(n_943),
.B1(n_825),
.B2(n_840),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_921),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_827),
.A2(n_854),
.B(n_785),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_840),
.B(n_911),
.Y(n_1093)
);

CKINVDCx16_ASAP7_75t_R g1094 ( 
.A(n_875),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_911),
.B(n_952),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_799),
.Y(n_1096)
);

AND2x6_ASAP7_75t_L g1097 ( 
.A(n_916),
.B(n_943),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_834),
.A2(n_878),
.B(n_948),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_890),
.B(n_936),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_948),
.A2(n_787),
.B(n_846),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_932),
.A2(n_900),
.B1(n_888),
.B2(n_895),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_846),
.A2(n_859),
.B(n_867),
.Y(n_1102)
);

CKINVDCx16_ASAP7_75t_R g1103 ( 
.A(n_956),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_958),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_926),
.A2(n_928),
.B(n_947),
.C(n_944),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1087),
.A2(n_954),
.B(n_963),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1054),
.A2(n_859),
.B(n_949),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1010),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1092),
.A2(n_963),
.B(n_958),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_989),
.A2(n_949),
.B(n_950),
.C(n_957),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1055),
.A2(n_950),
.B(n_957),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1034),
.A2(n_781),
.B(n_906),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_999),
.A2(n_942),
.B(n_1000),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1039),
.B(n_942),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1017),
.B(n_972),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1089),
.A2(n_1078),
.B(n_1068),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_1010),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_982),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1008),
.B(n_970),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1074),
.A2(n_1050),
.B(n_1007),
.C(n_1015),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_977),
.A2(n_999),
.A3(n_1090),
.B(n_1075),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1100),
.A2(n_1098),
.B(n_998),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1090),
.A2(n_1080),
.A3(n_1057),
.B(n_1105),
.Y(n_1123)
);

AOI21x1_ASAP7_75t_L g1124 ( 
.A1(n_988),
.A2(n_994),
.B(n_1057),
.Y(n_1124)
);

OAI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_993),
.A2(n_1047),
.B1(n_1029),
.B2(n_1012),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1056),
.A2(n_969),
.B(n_1088),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1056),
.A2(n_1099),
.B(n_974),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1094),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1077),
.A2(n_1085),
.B(n_966),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1014),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1008),
.B(n_1071),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_966),
.A2(n_1101),
.B(n_974),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1023),
.A2(n_1049),
.B(n_1040),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1021),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1035),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1102),
.A2(n_1004),
.B(n_1020),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1019),
.A2(n_1029),
.B(n_1013),
.C(n_1036),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_976),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1010),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1042),
.A2(n_1027),
.B(n_1045),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_1063),
.B(n_1070),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_978),
.A2(n_1044),
.B1(n_996),
.B2(n_968),
.Y(n_1142)
);

NAND2x1_ASAP7_75t_L g1143 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1042),
.A2(n_1048),
.B(n_1046),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1072),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1091),
.B(n_979),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1031),
.A2(n_1104),
.B(n_1082),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1063),
.B(n_1070),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1059),
.B(n_1060),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1052),
.A2(n_1051),
.B(n_1022),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1024),
.A2(n_1093),
.B(n_980),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_984),
.B(n_997),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1062),
.A2(n_1103),
.B1(n_973),
.B2(n_1063),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1095),
.A2(n_1001),
.B(n_987),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_992),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1041),
.A2(n_981),
.B(n_1064),
.Y(n_1156)
);

INVx5_ASAP7_75t_L g1157 ( 
.A(n_1063),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1066),
.A2(n_1079),
.B(n_1083),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1043),
.A2(n_986),
.B(n_1096),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1070),
.A2(n_1038),
.B1(n_983),
.B2(n_1005),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1043),
.A2(n_1096),
.B(n_1086),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1047),
.Y(n_1162)
);

INVxp67_ASAP7_75t_SL g1163 ( 
.A(n_990),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1011),
.A2(n_1065),
.A3(n_1081),
.B(n_1069),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1067),
.A2(n_1018),
.B(n_1026),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_995),
.A2(n_1028),
.B(n_1030),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1025),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1070),
.B(n_975),
.Y(n_1168)
);

O2A1O1Ixp5_ASAP7_75t_SL g1169 ( 
.A1(n_1061),
.A2(n_985),
.B(n_1097),
.C(n_1076),
.Y(n_1169)
);

OAI22x1_ASAP7_75t_L g1170 ( 
.A1(n_1084),
.A2(n_1037),
.B1(n_1016),
.B2(n_1047),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_975),
.B(n_1002),
.Y(n_1171)
);

O2A1O1Ixp5_ASAP7_75t_L g1172 ( 
.A1(n_1006),
.A2(n_971),
.B(n_992),
.C(n_1097),
.Y(n_1172)
);

AO21x1_ASAP7_75t_L g1173 ( 
.A1(n_1006),
.A2(n_1097),
.B(n_971),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_975),
.B(n_1002),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1097),
.A2(n_1003),
.A3(n_1043),
.B(n_1053),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1043),
.Y(n_1176)
);

AOI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1032),
.A2(n_1033),
.B1(n_1053),
.B2(n_1073),
.Y(n_1177)
);

OAI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_967),
.A2(n_1002),
.B1(n_1073),
.B2(n_1058),
.Y(n_1178)
);

INVx5_ASAP7_75t_L g1179 ( 
.A(n_1073),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1032),
.A2(n_1033),
.B(n_1053),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_965),
.B(n_1033),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_991),
.B(n_491),
.Y(n_1182)
);

CKINVDCx9p33_ASAP7_75t_R g1183 ( 
.A(n_968),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1054),
.A2(n_877),
.B(n_871),
.Y(n_1184)
);

INVx8_ASAP7_75t_L g1185 ( 
.A(n_1063),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1054),
.A2(n_877),
.B(n_871),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_1074),
.A2(n_1050),
.B(n_814),
.C(n_1007),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1008),
.B(n_491),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1008),
.B(n_491),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_989),
.A2(n_1071),
.B(n_934),
.C(n_1044),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_989),
.A2(n_1015),
.B(n_999),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1054),
.A2(n_1087),
.B(n_1055),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_SL g1193 ( 
.A1(n_1074),
.A2(n_1050),
.B(n_814),
.C(n_1007),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_989),
.A2(n_1071),
.B(n_934),
.C(n_1044),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1094),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_992),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_982),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_1010),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_989),
.A2(n_934),
.B1(n_1013),
.B2(n_626),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1087),
.A2(n_913),
.B(n_1092),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_989),
.A2(n_1071),
.B(n_934),
.C(n_1044),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1009),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1087),
.A2(n_913),
.B(n_1092),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1008),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1054),
.A2(n_877),
.B(n_871),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1009),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1017),
.B(n_972),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_993),
.B(n_678),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1010),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_982),
.Y(n_1210)
);

AOI21xp33_ASAP7_75t_L g1211 ( 
.A1(n_989),
.A2(n_1015),
.B(n_999),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1087),
.A2(n_913),
.B(n_1092),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_977),
.A2(n_999),
.A3(n_1000),
.B(n_1090),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_999),
.A2(n_1000),
.B(n_805),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_993),
.B(n_611),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_SL g1216 ( 
.A(n_989),
.B(n_626),
.C(n_611),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_989),
.A2(n_1071),
.B(n_934),
.C(n_1044),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1094),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_989),
.A2(n_1071),
.B(n_934),
.C(n_1044),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_999),
.A2(n_1000),
.B(n_805),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_977),
.A2(n_999),
.A3(n_1000),
.B(n_1090),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_989),
.A2(n_1017),
.B1(n_1015),
.B2(n_1007),
.Y(n_1222)
);

AOI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_989),
.A2(n_1015),
.B(n_999),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1054),
.A2(n_877),
.B(n_871),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_989),
.A2(n_934),
.B1(n_1013),
.B2(n_626),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_SL g1226 ( 
.A(n_1094),
.B(n_611),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_982),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1087),
.A2(n_913),
.B(n_1092),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1054),
.A2(n_877),
.B(n_871),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1087),
.A2(n_913),
.B(n_1092),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1054),
.A2(n_1087),
.B(n_1055),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1017),
.A2(n_999),
.B(n_856),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_982),
.Y(n_1233)
);

AND2x2_ASAP7_75t_SL g1234 ( 
.A(n_989),
.B(n_920),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_993),
.B(n_611),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_999),
.A2(n_1000),
.B(n_805),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1009),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1017),
.B(n_972),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1054),
.A2(n_877),
.B(n_871),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_989),
.A2(n_934),
.B1(n_1013),
.B2(n_626),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1009),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_1094),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_989),
.A2(n_1071),
.B(n_934),
.C(n_1044),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_982),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_989),
.A2(n_457),
.B(n_463),
.C(n_1019),
.Y(n_1245)
);

CKINVDCx11_ASAP7_75t_R g1246 ( 
.A(n_1242),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1123),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1138),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1179),
.B(n_1168),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1208),
.B(n_1131),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1153),
.A2(n_1222),
.B1(n_1234),
.B2(n_1162),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1145),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1148),
.Y(n_1253)
);

INVx4_ASAP7_75t_SL g1254 ( 
.A(n_1175),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1199),
.A2(n_1240),
.B1(n_1225),
.B2(n_1142),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1119),
.B(n_1149),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1153),
.A2(n_1199),
.B1(n_1225),
.B2(n_1240),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1222),
.A2(n_1125),
.B1(n_1211),
.B2(n_1223),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1157),
.B(n_1179),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1211),
.A2(n_1223),
.B1(n_1191),
.B2(n_1170),
.Y(n_1260)
);

INVx8_ASAP7_75t_L g1261 ( 
.A(n_1185),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1130),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1142),
.A2(n_1132),
.B1(n_1207),
.B2(n_1238),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1134),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1118),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1132),
.A2(n_1160),
.B1(n_1220),
.B2(n_1214),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1115),
.A2(n_1207),
.B1(n_1238),
.B2(n_1214),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1160),
.A2(n_1236),
.B1(n_1220),
.B2(n_1113),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_1198),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1236),
.A2(n_1113),
.B1(n_1129),
.B2(n_1115),
.Y(n_1270)
);

AOI21xp33_ASAP7_75t_L g1271 ( 
.A1(n_1190),
.A2(n_1201),
.B(n_1194),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1128),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1217),
.B(n_1219),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1135),
.Y(n_1274)
);

CKINVDCx14_ASAP7_75t_R g1275 ( 
.A(n_1195),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1197),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1216),
.A2(n_1129),
.B1(n_1243),
.B2(n_1144),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1218),
.A2(n_1182),
.B1(n_1181),
.B2(n_1152),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1196),
.Y(n_1279)
);

BUFx2_ASAP7_75t_SL g1280 ( 
.A(n_1155),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1146),
.A2(n_1189),
.B1(n_1188),
.B2(n_1241),
.Y(n_1281)
);

NAND2x1p5_ASAP7_75t_L g1282 ( 
.A(n_1157),
.B(n_1179),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1202),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1206),
.A2(n_1237),
.B1(n_1167),
.B2(n_1204),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_1215),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1235),
.B(n_1171),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1114),
.A2(n_1140),
.B1(n_1163),
.B2(n_1127),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1183),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1155),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1174),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1245),
.A2(n_1137),
.B1(n_1232),
.B2(n_1114),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1185),
.A2(n_1114),
.B1(n_1166),
.B2(n_1157),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1117),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1198),
.Y(n_1294)
);

CKINVDCx6p67_ASAP7_75t_R g1295 ( 
.A(n_1198),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1178),
.B(n_1108),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1151),
.A2(n_1150),
.B1(n_1139),
.B2(n_1209),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1176),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1154),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1184),
.A2(n_1229),
.B(n_1224),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1185),
.A2(n_1121),
.B1(n_1177),
.B2(n_1126),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1117),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1139),
.A2(n_1209),
.B1(n_1186),
.B2(n_1239),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1226),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1110),
.A2(n_1205),
.B1(n_1161),
.B2(n_1156),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1210),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1168),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1227),
.A2(n_1244),
.B1(n_1233),
.B2(n_1173),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_R g1309 ( 
.A1(n_1120),
.A2(n_1187),
.B1(n_1193),
.B2(n_1123),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1164),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1158),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1121),
.B(n_1180),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1143),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1141),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1107),
.A2(n_1133),
.B1(n_1159),
.B2(n_1231),
.Y(n_1315)
);

CKINVDCx6p67_ASAP7_75t_R g1316 ( 
.A(n_1172),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1136),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1147),
.A2(n_1165),
.B1(n_1231),
.B2(n_1192),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1169),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1124),
.A2(n_1112),
.B(n_1221),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1192),
.A2(n_1109),
.B1(n_1111),
.B2(n_1213),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1122),
.A2(n_1106),
.B1(n_1221),
.B2(n_1213),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1175),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1175),
.Y(n_1324)
);

INVx6_ASAP7_75t_L g1325 ( 
.A(n_1116),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1213),
.A2(n_1221),
.B1(n_1200),
.B2(n_1203),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1212),
.A2(n_1194),
.B1(n_1201),
.B2(n_1190),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1228),
.A2(n_560),
.B1(n_989),
.B2(n_1222),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1230),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1148),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1222),
.A2(n_560),
.B1(n_989),
.B2(n_679),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1138),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1176),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1138),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1145),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1138),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1138),
.Y(n_1337)
);

INVx6_ASAP7_75t_L g1338 ( 
.A(n_1198),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1118),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1138),
.Y(n_1340)
);

BUFx2_ASAP7_75t_SL g1341 ( 
.A(n_1155),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1242),
.Y(n_1342)
);

BUFx8_ASAP7_75t_SL g1343 ( 
.A(n_1128),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1222),
.A2(n_560),
.B1(n_989),
.B2(n_679),
.Y(n_1344)
);

BUFx8_ASAP7_75t_L g1345 ( 
.A(n_1162),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1222),
.A2(n_560),
.B1(n_989),
.B2(n_679),
.Y(n_1346)
);

BUFx8_ASAP7_75t_L g1347 ( 
.A(n_1162),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1225),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1138),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1198),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1176),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1242),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1176),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1138),
.Y(n_1354)
);

BUFx8_ASAP7_75t_SL g1355 ( 
.A(n_1128),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1118),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1176),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1153),
.A2(n_560),
.B1(n_989),
.B2(n_934),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1176),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1138),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1199),
.A2(n_1240),
.B1(n_1225),
.B2(n_1142),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1138),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1222),
.A2(n_560),
.B1(n_989),
.B2(n_679),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1196),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1131),
.B(n_1119),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1138),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1148),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1145),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1247),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1256),
.B(n_1365),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1331),
.A2(n_1344),
.B1(n_1363),
.B2(n_1346),
.C(n_1361),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1271),
.A2(n_1273),
.B(n_1361),
.C(n_1255),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1290),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1247),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1310),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1312),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1343),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1311),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1255),
.A2(n_1348),
.B(n_1291),
.C(n_1327),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1317),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1248),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1262),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1254),
.B(n_1299),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1263),
.B(n_1267),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1329),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1300),
.A2(n_1315),
.B(n_1305),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1264),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1274),
.Y(n_1388)
);

NAND2xp33_ASAP7_75t_SL g1389 ( 
.A(n_1277),
.B(n_1288),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1283),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1332),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1246),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1325),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1325),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1334),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1323),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1263),
.B(n_1267),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1299),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1266),
.A2(n_1268),
.B1(n_1344),
.B2(n_1331),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1268),
.B(n_1266),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1318),
.A2(n_1321),
.B(n_1320),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1336),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1337),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1340),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1358),
.A2(n_1363),
.B1(n_1346),
.B2(n_1251),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1349),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1354),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1360),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1362),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1285),
.B(n_1286),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1366),
.Y(n_1411)
);

O2A1O1Ixp5_ASAP7_75t_L g1412 ( 
.A1(n_1287),
.A2(n_1297),
.B(n_1303),
.C(n_1326),
.Y(n_1412)
);

AO21x1_ASAP7_75t_L g1413 ( 
.A1(n_1287),
.A2(n_1326),
.B(n_1303),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1279),
.B(n_1272),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1342),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1318),
.A2(n_1321),
.B(n_1322),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1250),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1270),
.B(n_1260),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1316),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1324),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1308),
.A2(n_1258),
.B(n_1357),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1252),
.B(n_1335),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1270),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1257),
.B(n_1284),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1298),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1298),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1265),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1276),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1251),
.A2(n_1358),
.B1(n_1364),
.B2(n_1296),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1281),
.B(n_1368),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1253),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1306),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1281),
.B(n_1284),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1297),
.A2(n_1314),
.B(n_1356),
.Y(n_1434)
);

AOI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1249),
.A2(n_1309),
.B(n_1339),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1319),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1301),
.A2(n_1328),
.B(n_1292),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_SL g1438 ( 
.A1(n_1275),
.A2(n_1353),
.B(n_1359),
.C(n_1357),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1328),
.B(n_1333),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1333),
.A2(n_1351),
.B(n_1353),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1292),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1319),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1301),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1278),
.A2(n_1359),
.B(n_1259),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1319),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1261),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1261),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1373),
.B(n_1352),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1373),
.B(n_1383),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1379),
.A2(n_1313),
.B(n_1341),
.C(n_1280),
.Y(n_1450)
);

AO32x2_ASAP7_75t_L g1451 ( 
.A1(n_1396),
.A2(n_1294),
.A3(n_1304),
.B1(n_1307),
.B2(n_1293),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1399),
.A2(n_1347),
.B1(n_1345),
.B2(n_1269),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1399),
.A2(n_1400),
.B1(n_1429),
.B2(n_1418),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1419),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1417),
.B(n_1367),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1381),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1372),
.A2(n_1282),
.B(n_1294),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1295),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1402),
.B(n_1330),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1413),
.A2(n_1412),
.B(n_1386),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1400),
.A2(n_1347),
.B(n_1345),
.C(n_1289),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1419),
.B(n_1302),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1402),
.B(n_1355),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1371),
.A2(n_1338),
.B1(n_1350),
.B2(n_1302),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1440),
.Y(n_1466)
);

CKINVDCx6p67_ASAP7_75t_R g1467 ( 
.A(n_1377),
.Y(n_1467)
);

AOI22x1_ASAP7_75t_SL g1468 ( 
.A1(n_1392),
.A2(n_1338),
.B1(n_1350),
.B2(n_1415),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1423),
.A2(n_1350),
.B1(n_1424),
.B2(n_1405),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1398),
.B(n_1376),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1410),
.B(n_1422),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1389),
.B(n_1430),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1413),
.A2(n_1386),
.B(n_1398),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1414),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1425),
.B(n_1426),
.Y(n_1475)
);

NAND4xp25_ASAP7_75t_L g1476 ( 
.A(n_1384),
.B(n_1397),
.C(n_1438),
.D(n_1433),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1376),
.B(n_1384),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1431),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1425),
.B(n_1426),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1437),
.B(n_1421),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1401),
.A2(n_1416),
.B(n_1445),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1424),
.A2(n_1421),
.B(n_1443),
.C(n_1441),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1369),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1370),
.B(n_1444),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1445),
.A2(n_1442),
.B(n_1436),
.C(n_1439),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1436),
.A2(n_1442),
.B(n_1435),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1391),
.B(n_1404),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1395),
.B(n_1403),
.Y(n_1492)
);

AO32x2_ASAP7_75t_L g1493 ( 
.A1(n_1446),
.A2(n_1406),
.A3(n_1395),
.B1(n_1409),
.B2(n_1408),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1404),
.B(n_1406),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1493),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1470),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1493),
.B(n_1380),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1493),
.B(n_1380),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1453),
.A2(n_1439),
.B1(n_1407),
.B2(n_1434),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1470),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1477),
.B(n_1407),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1456),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1466),
.B(n_1393),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1454),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1374),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1478),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1486),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1454),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1486),
.B(n_1374),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1483),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1494),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1476),
.A2(n_1436),
.B1(n_1434),
.B2(n_1432),
.Y(n_1512)
);

NOR2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1476),
.B(n_1447),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1482),
.B(n_1484),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1449),
.B(n_1394),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1459),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1481),
.A2(n_1428),
.B1(n_1427),
.B2(n_1375),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1378),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1459),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1496),
.B(n_1487),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1496),
.B(n_1491),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1501),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1497),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1497),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1500),
.B(n_1487),
.Y(n_1527)
);

OAI321xp33_ASAP7_75t_L g1528 ( 
.A1(n_1499),
.A2(n_1481),
.A3(n_1485),
.B1(n_1472),
.B2(n_1461),
.C(n_1490),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1509),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1516),
.A2(n_1495),
.B(n_1520),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1498),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1499),
.A2(n_1472),
.B1(n_1469),
.B2(n_1452),
.Y(n_1534)
);

OAI211xp5_ASAP7_75t_L g1535 ( 
.A1(n_1499),
.A2(n_1461),
.B(n_1462),
.C(n_1450),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1507),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.B(n_1475),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1480),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1516),
.A2(n_1490),
.B(n_1458),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1467),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1507),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1502),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1502),
.Y(n_1543)
);

OAI33xp33_ASAP7_75t_L g1544 ( 
.A1(n_1501),
.A2(n_1458),
.A3(n_1464),
.B1(n_1455),
.B2(n_1488),
.B3(n_1460),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1502),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1521),
.B(n_1471),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1520),
.A2(n_1465),
.B1(n_1457),
.B2(n_1420),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1517),
.Y(n_1548)
);

OAI31xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1504),
.A2(n_1463),
.A3(n_1448),
.B(n_1451),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1506),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_R g1552 ( 
.A(n_1514),
.B(n_1468),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1498),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1518),
.B(n_1479),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1536),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1525),
.B(n_1514),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1532),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1525),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1542),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1542),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1550),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1518),
.Y(n_1566)
);

AND2x4_ASAP7_75t_SL g1567 ( 
.A(n_1554),
.B(n_1515),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1543),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1543),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1545),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1534),
.A2(n_1513),
.B1(n_1512),
.B2(n_1519),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1545),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1524),
.B(n_1511),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1533),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1522),
.B(n_1511),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1539),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1550),
.B(n_1506),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1548),
.B(n_1508),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1550),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1539),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1549),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1527),
.B(n_1511),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1562),
.Y(n_1585)
);

NAND2xp67_ASAP7_75t_SL g1586 ( 
.A(n_1583),
.B(n_1546),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1562),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1556),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1563),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1581),
.B(n_1549),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1579),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1567),
.B(n_1531),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1558),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1563),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1563),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1577),
.B(n_1541),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1556),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1556),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1565),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1568),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1559),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1568),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1568),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1579),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1569),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1546),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1577),
.B(n_1541),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1583),
.B(n_1554),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1567),
.B(n_1551),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1569),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1569),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1570),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1570),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1584),
.B(n_1523),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_L g1616 ( 
.A(n_1581),
.B(n_1513),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1570),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1551),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1560),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1523),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1573),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1575),
.B(n_1537),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1558),
.B(n_1537),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1567),
.B(n_1538),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1573),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1592),
.B(n_1580),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1609),
.B(n_1565),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1626),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1626),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1605),
.B(n_1580),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1609),
.B(n_1565),
.Y(n_1632)
);

NAND2x1_ASAP7_75t_L g1633 ( 
.A(n_1593),
.B(n_1565),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1622),
.B(n_1555),
.Y(n_1636)
);

OR2x6_ASAP7_75t_L g1637 ( 
.A(n_1588),
.B(n_1535),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1607),
.B(n_1557),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1585),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1586),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1594),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1607),
.B(n_1575),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1587),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1622),
.B(n_1574),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1587),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1589),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1625),
.B(n_1557),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1625),
.B(n_1557),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1624),
.B(n_1566),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1566),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1589),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1590),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1566),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1574),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1602),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1590),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1615),
.B(n_1620),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1593),
.B(n_1572),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1600),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1595),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1629),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1635),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1637),
.A2(n_1572),
.B1(n_1534),
.B2(n_1528),
.Y(n_1664)
);

CKINVDCx16_ASAP7_75t_R g1665 ( 
.A(n_1637),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1658),
.B(n_1620),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1637),
.A2(n_1616),
.B(n_1619),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1637),
.A2(n_1560),
.B1(n_1582),
.B2(n_1578),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1640),
.A2(n_1598),
.B(n_1588),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1627),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1628),
.B(n_1540),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1641),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1644),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1640),
.A2(n_1599),
.B(n_1598),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1629),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1602),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1659),
.A2(n_1544),
.B1(n_1547),
.B2(n_1552),
.Y(n_1678)
);

AOI31xp33_ASAP7_75t_L g1679 ( 
.A1(n_1631),
.A2(n_1586),
.A3(n_1593),
.B(n_1618),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_R g1680 ( 
.A(n_1628),
.B(n_1600),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1633),
.A2(n_1599),
.B(n_1578),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1632),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1632),
.B(n_1610),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1630),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1638),
.A2(n_1571),
.B(n_1582),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1630),
.Y(n_1686)
);

NOR4xp25_ASAP7_75t_L g1687 ( 
.A(n_1672),
.B(n_1660),
.C(n_1656),
.D(n_1657),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1665),
.B(n_1670),
.Y(n_1688)
);

AOI321xp33_ASAP7_75t_L g1689 ( 
.A1(n_1664),
.A2(n_1578),
.A3(n_1582),
.B1(n_1656),
.B2(n_1512),
.C(n_1647),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1675),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1675),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1662),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_SL g1693 ( 
.A(n_1676),
.B(n_1647),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1679),
.A2(n_1636),
.B(n_1655),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1682),
.B(n_1666),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1678),
.A2(n_1582),
.B(n_1578),
.C(n_1571),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1668),
.A2(n_1571),
.B1(n_1653),
.B2(n_1633),
.C(n_1661),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1671),
.B(n_1654),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1683),
.Y(n_1699)
);

OAI322xp33_ASAP7_75t_L g1700 ( 
.A1(n_1664),
.A2(n_1661),
.A3(n_1657),
.B1(n_1639),
.B2(n_1652),
.C1(n_1651),
.C2(n_1643),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1667),
.A2(n_1639),
.B(n_1634),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1680),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1683),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1677),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1663),
.B(n_1654),
.Y(n_1705)
);

AOI32xp33_ASAP7_75t_L g1706 ( 
.A1(n_1702),
.A2(n_1668),
.A3(n_1686),
.B1(n_1684),
.B2(n_1648),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1699),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1693),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1699),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1705),
.B(n_1673),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1703),
.B(n_1649),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1703),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1704),
.B(n_1648),
.Y(n_1713)
);

AO22x1_ASAP7_75t_L g1714 ( 
.A1(n_1698),
.A2(n_1685),
.B1(n_1680),
.B2(n_1649),
.Y(n_1714)
);

AOI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1700),
.A2(n_1687),
.B(n_1697),
.C(n_1694),
.Y(n_1715)
);

XNOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1688),
.B(n_1513),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_L g1717 ( 
.A(n_1716),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1715),
.A2(n_1696),
.B1(n_1704),
.B2(n_1674),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1710),
.B(n_1705),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1711),
.B(n_1691),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1711),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1706),
.B(n_1696),
.C(n_1689),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1714),
.A2(n_1669),
.B1(n_1695),
.B2(n_1691),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1713),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1707),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1722),
.A2(n_1701),
.B1(n_1712),
.B2(n_1709),
.C(n_1708),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1721),
.Y(n_1727)
);

NAND4xp75_ASAP7_75t_L g1728 ( 
.A(n_1718),
.B(n_1690),
.C(n_1692),
.D(n_1681),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_L g1729 ( 
.A(n_1725),
.B(n_1634),
.C(n_1652),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1723),
.A2(n_1693),
.B(n_1651),
.C(n_1646),
.Y(n_1730)
);

XNOR2x1_ASAP7_75t_L g1731 ( 
.A(n_1728),
.B(n_1724),
.Y(n_1731)
);

OAI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1726),
.A2(n_1730),
.B(n_1727),
.C(n_1719),
.Y(n_1732)
);

XNOR2xp5_ASAP7_75t_L g1733 ( 
.A(n_1729),
.B(n_1720),
.Y(n_1733)
);

AOI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1730),
.A2(n_1717),
.B(n_1646),
.C(n_1645),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1727),
.A2(n_1474),
.B1(n_1645),
.B2(n_1643),
.Y(n_1735)
);

OAI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1726),
.A2(n_1650),
.B(n_1621),
.C(n_1604),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1731),
.Y(n_1737)
);

OAI322xp33_ASAP7_75t_L g1738 ( 
.A1(n_1733),
.A2(n_1608),
.A3(n_1597),
.B1(n_1595),
.B2(n_1617),
.C1(n_1614),
.C2(n_1613),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1735),
.B(n_1650),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1732),
.B(n_1736),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1734),
.B(n_1618),
.Y(n_1741)
);

NAND4xp25_ASAP7_75t_L g1742 ( 
.A(n_1740),
.B(n_1593),
.C(n_1506),
.D(n_1597),
.Y(n_1742)
);

NAND4xp75_ASAP7_75t_L g1743 ( 
.A(n_1741),
.B(n_1737),
.C(n_1739),
.D(n_1738),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1737),
.B(n_1741),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1743),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1744),
.B1(n_1742),
.B2(n_1621),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

AOI21xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1746),
.A2(n_1745),
.B(n_1617),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1747),
.A2(n_1614),
.B(n_1613),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1748),
.A2(n_1608),
.B1(n_1611),
.B2(n_1612),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1749),
.A2(n_1612),
.B1(n_1611),
.B2(n_1606),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1750),
.A2(n_1606),
.B1(n_1604),
.B2(n_1603),
.Y(n_1752)
);

XNOR2x1_ASAP7_75t_L g1753 ( 
.A(n_1751),
.B(n_1752),
.Y(n_1753)
);

AOI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1603),
.B(n_1601),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1601),
.B1(n_1596),
.B2(n_1564),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1596),
.B1(n_1561),
.B2(n_1576),
.C(n_1573),
.Y(n_1756)
);

AOI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1564),
.B(n_1555),
.C(n_1576),
.Y(n_1757)
);


endmodule