module fake_netlist_6_225_n_386 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_386);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_386;

wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_350;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_122;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_352;
wire n_374;
wire n_366;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_277;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_364;
wire n_295;
wire n_385;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_0),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_37),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_19),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_4),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_14),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_50),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_41),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_68),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_70),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_20),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_29),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_21),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_39),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_53),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_46),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_9),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_52),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_44),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_32),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_96),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_72),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_35),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_7),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_30),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_31),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_77),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_33),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_58),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_34),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_66),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_132),
.B(n_0),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

OAI22x1_ASAP7_75t_R g183 ( 
.A1(n_169),
.A2(n_176),
.B1(n_136),
.B2(n_148),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_1),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_135),
.B(n_2),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_3),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_6),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_8),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_10),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_11),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_165),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_122),
.C(n_156),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_180),
.B(n_149),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_130),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_191),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_156),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_179),
.B(n_173),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_173),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_140),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_154),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_199),
.B1(n_157),
.B2(n_178),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_141),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_126),
.Y(n_234)
);

NOR2x2_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_183),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_142),
.B1(n_175),
.B2(n_174),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_218),
.B(n_225),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_222),
.B1(n_214),
.B2(n_211),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_143),
.B(n_144),
.C(n_171),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

NOR2x1p5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_129),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_150),
.B(n_152),
.C(n_153),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_158),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

NOR2x1p5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_131),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_159),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_160),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_133),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_164),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_226),
.B(n_167),
.Y(n_259)
);

BUFx6f_ASAP7_75t_SL g260 ( 
.A(n_226),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_208),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_211),
.B(n_161),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_166),
.B(n_172),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_177),
.B(n_168),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_241),
.B1(n_259),
.B2(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g268 ( 
.A(n_260),
.B(n_155),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_151),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_139),
.B(n_137),
.Y(n_270)
);

OR2x6_ASAP7_75t_SL g271 ( 
.A(n_235),
.B(n_15),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

AOI211xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_16),
.B(n_18),
.C(n_22),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_23),
.B(n_24),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_25),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_230),
.A2(n_42),
.B1(n_43),
.B2(n_47),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_48),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_49),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

OR2x6_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_54),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_56),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_57),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_59),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_60),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_233),
.A2(n_62),
.B(n_63),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_257),
.B(n_256),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_240),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_253),
.B(n_245),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_242),
.B(n_240),
.Y(n_293)
);

AO31x2_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_65),
.A3(n_67),
.B(n_69),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_71),
.B(n_74),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_265),
.Y(n_296)
);

AO31x2_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_76),
.A3(n_78),
.B(n_79),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_118),
.B(n_83),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_277),
.B(n_81),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_85),
.B(n_86),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_87),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_88),
.B(n_89),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_268),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_91),
.Y(n_305)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_94),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_95),
.B1(n_102),
.B2(n_103),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_289),
.B(n_275),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_280),
.B(n_288),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

AO21x2_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_278),
.B(n_270),
.Y(n_316)
);

AO31x2_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_274),
.A3(n_271),
.B(n_109),
.Y(n_317)
);

BUFx8_ASAP7_75t_SL g318 ( 
.A(n_301),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_304),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_273),
.C(n_107),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_104),
.B(n_110),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_308),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_306),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_306),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_298),
.B(n_295),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_320),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_324),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_317),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_317),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_317),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_317),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_306),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_308),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_327),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_338),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_341),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_333),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_337),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_328),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_345),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_353),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_345),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_345),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_352),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_351),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_364),
.A2(n_344),
.B(n_348),
.C(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_368),
.Y(n_369)
);

OAI221xp5_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_365),
.B1(n_362),
.B2(n_358),
.C(n_337),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_344),
.B1(n_361),
.B2(n_356),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_369),
.A2(n_344),
.B1(n_356),
.B2(n_358),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_294),
.Y(n_373)
);

OAI211xp5_ASAP7_75t_SL g374 ( 
.A1(n_372),
.A2(n_300),
.B(n_309),
.C(n_314),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_373),
.B(n_294),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

AND2x2_ASAP7_75t_SL g377 ( 
.A(n_376),
.B(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_377),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_297),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_114),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_374),
.B(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_115),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_293),
.B(n_331),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_383),
.A2(n_316),
.B(n_331),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_384),
.B1(n_332),
.B2(n_328),
.Y(n_386)
);


endmodule