module fake_jpeg_16934_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_20),
.B1(n_18),
.B2(n_24),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_24),
.B1(n_26),
.B2(n_13),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_20),
.B1(n_18),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_27),
.B2(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_25),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_18),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_30),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_48),
.B(n_40),
.C(n_4),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_16),
.B1(n_14),
.B2(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_58),
.B1(n_0),
.B2(n_2),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_25),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_15),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_25),
.B1(n_15),
.B2(n_3),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_0),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_0),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_85),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_46),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_84),
.C(n_67),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_10),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_84),
.B(n_2),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_10),
.Y(n_85)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_3),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_51),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_93),
.B(n_102),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_50),
.B(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_50),
.B1(n_51),
.B2(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_98),
.B1(n_83),
.B2(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_61),
.B1(n_80),
.B2(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_64),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_78),
.B1(n_88),
.B2(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_117),
.B1(n_122),
.B2(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_119),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_118),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_77),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_70),
.B1(n_40),
.B2(n_48),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_90),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_82),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_95),
.C(n_93),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.C(n_136),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_92),
.C(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_106),
.B1(n_118),
.B2(n_92),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_121),
.B(n_110),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_138),
.Y(n_142)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_98),
.C(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_124),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_99),
.C(n_107),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_147),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_117),
.A3(n_125),
.B1(n_109),
.B2(n_91),
.C1(n_113),
.C2(n_114),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_146),
.B(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_120),
.B1(n_107),
.B2(n_122),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_148),
.B1(n_9),
.B2(n_146),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_128),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_153),
.C(n_154),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_5),
.C(n_8),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_153),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_149),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_146),
.B(n_140),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_167),
.B(n_160),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_169),
.C(n_166),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_172),
.B(n_169),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_163),
.B1(n_164),
.B2(n_142),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_148),
.Y(n_176)
);


endmodule