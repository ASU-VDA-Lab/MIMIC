module fake_netlist_6_4799_n_866 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_866);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_866;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

BUFx2_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_50),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_60),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_45),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_185),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_82),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_99),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_121),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_85),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_54),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_58),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_1),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_24),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_107),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_41),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_33),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_73),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_38),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_96),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_117),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_119),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_13),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_112),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_128),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_184),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_131),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_20),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_18),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_48),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_95),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_129),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_89),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_70),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_37),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_81),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_0),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_98),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_190),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_152),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_146),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_67),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_147),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_35),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_0),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_195),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_2),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_2),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_238),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_231),
.B(n_3),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_227),
.B(n_26),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_3),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_27),
.Y(n_294)
);

BUFx8_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_254),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_197),
.B(n_4),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_250),
.B(n_4),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_198),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_199),
.B(n_28),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_202),
.B(n_5),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_5),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_215),
.B(n_259),
.Y(n_307)
);

BUFx8_ASAP7_75t_SL g308 ( 
.A(n_219),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_204),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_208),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g311 ( 
.A(n_196),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_220),
.B(n_6),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_222),
.B(n_229),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_232),
.B(n_29),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_200),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_201),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_203),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_219),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_240),
.B(n_6),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_249),
.B(n_7),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_251),
.B(n_30),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_307),
.B1(n_277),
.B2(n_293),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_215),
.B1(n_259),
.B2(n_266),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_7),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_258),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_207),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_301),
.A2(n_275),
.B1(n_273),
.B2(n_260),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_279),
.A2(n_266),
.B1(n_205),
.B2(n_276),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_209),
.Y(n_336)
);

AO22x2_ASAP7_75t_L g337 ( 
.A1(n_293),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_279),
.A2(n_272),
.B1(n_270),
.B2(n_269),
.Y(n_338)
);

AO22x2_ASAP7_75t_L g339 ( 
.A1(n_281),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_268),
.B1(n_267),
.B2(n_264),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_281),
.A2(n_255),
.B1(n_246),
.B2(n_245),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_282),
.A2(n_244),
.B1(n_243),
.B2(n_241),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_288),
.B(n_210),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_322),
.A2(n_223),
.B1(n_235),
.B2(n_234),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_211),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_217),
.B1(n_233),
.B2(n_228),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_297),
.B(n_212),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_288),
.A2(n_226),
.B1(n_225),
.B2(n_216),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_290),
.B(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_239),
.B1(n_214),
.B2(n_213),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_299),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_32),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_306),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_305),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g363 ( 
.A(n_289),
.B(n_14),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_313),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_296),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_300),
.B(n_317),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_289),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_34),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_289),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_286),
.B(n_310),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_287),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_284),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_308),
.B(n_25),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_314),
.B(n_36),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_303),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_43),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_304),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_287),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

XOR2x2_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_314),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_304),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_329),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_354),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_331),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_330),
.B(n_311),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_316),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_350),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_363),
.B(n_311),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_304),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_352),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_327),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_319),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_327),
.B(n_315),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_353),
.B(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_353),
.A2(n_345),
.B(n_356),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_338),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

NAND2x1p5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_315),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_R g417 ( 
.A(n_359),
.B(n_315),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_356),
.B(n_303),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_351),
.B(n_278),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_370),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_339),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_335),
.B(n_319),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_361),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

OR2x2_ASAP7_75t_SL g432 ( 
.A(n_361),
.B(n_278),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_326),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_365),
.B(n_326),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_346),
.B(n_319),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_376),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_358),
.B(n_285),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_330),
.B(n_319),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_354),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_330),
.B(n_319),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_395),
.B(n_326),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_320),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_285),
.Y(n_454)
);

AND2x2_ASAP7_75t_SL g455 ( 
.A(n_408),
.B(n_318),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_292),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_442),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_320),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_292),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_406),
.A2(n_294),
.B(n_323),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_391),
.B(n_292),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_320),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_440),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_382),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_324),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_324),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_419),
.B(n_433),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_397),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_437),
.A2(n_294),
.B(n_323),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_408),
.A2(n_294),
.B(n_323),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_445),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_435),
.B(n_324),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_435),
.B(n_324),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_318),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_396),
.B(n_318),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_398),
.B(n_438),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_413),
.B(n_320),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_446),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_388),
.B(n_320),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_387),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_439),
.B(n_318),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_400),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_323),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_422),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_404),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_410),
.B(n_323),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_426),
.A2(n_294),
.B(n_295),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_294),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_415),
.B(n_294),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_417),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_49),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_405),
.A2(n_295),
.B(n_52),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_295),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_389),
.B(n_51),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_425),
.B(n_53),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_431),
.B(n_55),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_455),
.B(n_389),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_454),
.B(n_423),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_514),
.B(n_404),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_455),
.B(n_429),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_488),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_434),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_451),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_455),
.B(n_448),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_448),
.B(n_429),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_454),
.B(n_384),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_471),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_436),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_471),
.B(n_436),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_477),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_467),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_467),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_427),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_474),
.B(n_441),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_477),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_467),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_457),
.B(n_384),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_469),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_469),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_474),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_399),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_496),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_469),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_484),
.B(n_447),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_465),
.B(n_428),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_484),
.B(n_447),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_495),
.B(n_432),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_496),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_470),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_456),
.B(n_401),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_488),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_486),
.B(n_409),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_482),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_514),
.B(n_430),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_486),
.B(n_412),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_417),
.Y(n_561)
);

NAND2x1p5_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_56),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_475),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_456),
.B(n_385),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_499),
.B(n_430),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_495),
.B(n_57),
.Y(n_567)
);

NAND2x1_ASAP7_75t_SL g568 ( 
.A(n_512),
.B(n_61),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_493),
.B(n_62),
.Y(n_569)
);

CKINVDCx11_ASAP7_75t_R g570 ( 
.A(n_499),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_465),
.B(n_63),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_487),
.B(n_64),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_537),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_557),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_537),
.Y(n_576)
);

CKINVDCx8_ASAP7_75t_R g577 ( 
.A(n_566),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_559),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

CKINVDCx8_ASAP7_75t_R g580 ( 
.A(n_522),
.Y(n_580)
);

BUFx12f_ASAP7_75t_L g581 ( 
.A(n_570),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_544),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_523),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_535),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_535),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_527),
.B(n_489),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_550),
.Y(n_587)
);

BUFx2_ASAP7_75t_R g588 ( 
.A(n_522),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_544),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_565),
.A2(n_489),
.B1(n_488),
.B2(n_493),
.Y(n_590)
);

INVx6_ASAP7_75t_SL g591 ( 
.A(n_569),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_526),
.B(n_461),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_537),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_569),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_524),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_535),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_524),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_529),
.B(n_461),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_528),
.B(n_507),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_570),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_520),
.A2(n_481),
.B1(n_515),
.B2(n_508),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_569),
.Y(n_606)
);

BUFx4f_ASAP7_75t_SL g607 ( 
.A(n_554),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_564),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_559),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_523),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_518),
.Y(n_612)
);

BUFx4f_ASAP7_75t_SL g613 ( 
.A(n_542),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_547),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

BUFx6f_ASAP7_75t_SL g616 ( 
.A(n_550),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_575),
.Y(n_617)
);

INVx6_ASAP7_75t_L g618 ( 
.A(n_581),
.Y(n_618)
);

CKINVDCx6p67_ASAP7_75t_R g619 ( 
.A(n_581),
.Y(n_619)
);

CKINVDCx11_ASAP7_75t_R g620 ( 
.A(n_603),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_590),
.A2(n_519),
.B1(n_558),
.B2(n_489),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_576),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_615),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_586),
.A2(n_539),
.B1(n_517),
.B2(n_542),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_587),
.A2(n_555),
.B1(n_525),
.B2(n_498),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_594),
.A2(n_555),
.B1(n_508),
.B2(n_515),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_603),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_574),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_583),
.A2(n_530),
.B1(n_560),
.B2(n_450),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_600),
.A2(n_560),
.B1(n_450),
.B2(n_561),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_610),
.A2(n_560),
.B1(n_450),
.B2(n_500),
.Y(n_632)
);

INVx6_ASAP7_75t_L g633 ( 
.A(n_611),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_612),
.A2(n_463),
.B1(n_472),
.B2(n_466),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_596),
.Y(n_635)
);

CKINVDCx11_ASAP7_75t_R g636 ( 
.A(n_577),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_596),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_578),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_611),
.Y(n_639)
);

CKINVDCx14_ASAP7_75t_R g640 ( 
.A(n_578),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_605),
.A2(n_516),
.B1(n_551),
.B2(n_547),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_599),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_604),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_604),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_598),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_L g649 ( 
.A1(n_608),
.A2(n_483),
.B1(n_463),
.B2(n_462),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_601),
.B(n_458),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_SL g651 ( 
.A1(n_594),
.A2(n_509),
.B1(n_481),
.B2(n_572),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_612),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_616),
.A2(n_483),
.B1(n_462),
.B2(n_463),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_592),
.A2(n_491),
.B1(n_459),
.B2(n_567),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_607),
.A2(n_466),
.B1(n_472),
.B2(n_483),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_605),
.A2(n_546),
.B(n_536),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_625),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_621),
.A2(n_594),
.B1(n_606),
.B2(n_616),
.Y(n_660)
);

BUFx4f_ASAP7_75t_SL g661 ( 
.A(n_619),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_626),
.B(n_602),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_627),
.A2(n_607),
.B1(n_472),
.B2(n_462),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_638),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_640),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_656),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_651),
.A2(n_606),
.B1(n_594),
.B2(n_580),
.Y(n_667)
);

AND2x4_ASAP7_75t_SL g668 ( 
.A(n_629),
.B(n_576),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_630),
.A2(n_466),
.B1(n_611),
.B2(n_606),
.Y(n_669)
);

BUFx8_ASAP7_75t_L g670 ( 
.A(n_624),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_649),
.A2(n_611),
.B1(n_606),
.B2(n_591),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_636),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_631),
.A2(n_591),
.B1(n_491),
.B2(n_605),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_623),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_654),
.A2(n_591),
.B1(n_613),
.B2(n_617),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_633),
.A2(n_562),
.B1(n_572),
.B2(n_580),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_635),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_652),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_642),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_644),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_637),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_646),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_620),
.Y(n_683)
);

BUFx12f_ASAP7_75t_L g684 ( 
.A(n_618),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_647),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_656),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_648),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_656),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_618),
.A2(n_562),
.B1(n_639),
.B2(n_633),
.Y(n_689)
);

BUFx12f_ASAP7_75t_L g690 ( 
.A(n_639),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_632),
.A2(n_459),
.B1(n_584),
.B2(n_585),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_657),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_622),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_SL g694 ( 
.A(n_629),
.B(n_568),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_655),
.A2(n_585),
.B1(n_597),
.B2(n_501),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_653),
.B(n_609),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_622),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_622),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_645),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_654),
.A2(n_597),
.B1(n_501),
.B2(n_502),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_SL g701 ( 
.A1(n_628),
.A2(n_613),
.B1(n_588),
.B2(n_614),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_634),
.A2(n_516),
.B1(n_614),
.B2(n_595),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_645),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_645),
.B(n_598),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_659),
.A2(n_595),
.B1(n_492),
.B2(n_502),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_667),
.A2(n_641),
.B1(n_543),
.B2(n_516),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_662),
.A2(n_660),
.B1(n_675),
.B2(n_673),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_696),
.A2(n_503),
.B1(n_658),
.B2(n_548),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_678),
.B(n_485),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_687),
.B(n_485),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_663),
.A2(n_503),
.B1(n_516),
.B2(n_556),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_692),
.B(n_576),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_671),
.B(n_700),
.C(n_669),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_665),
.A2(n_516),
.B1(n_480),
.B2(n_543),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_674),
.B(n_681),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_683),
.A2(n_573),
.B1(n_579),
.B2(n_593),
.Y(n_716)
);

AOI221xp5_ASAP7_75t_L g717 ( 
.A1(n_676),
.A2(n_479),
.B1(n_460),
.B2(n_510),
.C(n_504),
.Y(n_717)
);

OAI211xp5_ASAP7_75t_L g718 ( 
.A1(n_689),
.A2(n_479),
.B(n_504),
.C(n_480),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_681),
.B(n_480),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_701),
.A2(n_516),
.B1(n_643),
.B2(n_574),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_682),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_698),
.B(n_593),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_695),
.A2(n_579),
.B1(n_551),
.B2(n_643),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_672),
.A2(n_532),
.B1(n_540),
.B2(n_541),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_SL g725 ( 
.A1(n_683),
.A2(n_579),
.B1(n_589),
.B2(n_582),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_691),
.A2(n_589),
.B1(n_582),
.B2(n_496),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_670),
.A2(n_506),
.B1(n_497),
.B2(n_490),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_672),
.A2(n_545),
.B1(n_563),
.B2(n_533),
.Y(n_728)
);

OAI221xp5_ASAP7_75t_L g729 ( 
.A1(n_694),
.A2(n_452),
.B1(n_464),
.B2(n_496),
.C(n_475),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_664),
.B(n_534),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_670),
.A2(n_449),
.B1(n_453),
.B2(n_476),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_664),
.A2(n_549),
.B1(n_538),
.B2(n_552),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_670),
.A2(n_684),
.B1(n_694),
.B2(n_702),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_682),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_679),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_677),
.Y(n_736)
);

OAI222xp33_ASAP7_75t_L g737 ( 
.A1(n_680),
.A2(n_513),
.B1(n_571),
.B2(n_553),
.C1(n_506),
.C2(n_449),
.Y(n_737)
);

AOI222xp33_ASAP7_75t_L g738 ( 
.A1(n_661),
.A2(n_453),
.B1(n_476),
.B2(n_506),
.C1(n_553),
.C2(n_571),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_690),
.A2(n_511),
.B1(n_513),
.B2(n_506),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_684),
.A2(n_476),
.B1(n_513),
.B2(n_478),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_679),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_699),
.B(n_65),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_707),
.B(n_685),
.C(n_703),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_736),
.B(n_697),
.Y(n_744)
);

OA21x2_ASAP7_75t_L g745 ( 
.A1(n_708),
.A2(n_703),
.B(n_697),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_715),
.B(n_699),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_SL g747 ( 
.A1(n_707),
.A2(n_668),
.B(n_704),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_SL g748 ( 
.A(n_725),
.B(n_690),
.C(n_666),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_L g749 ( 
.A1(n_708),
.A2(n_704),
.B1(n_666),
.B2(n_688),
.C(n_686),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_L g750 ( 
.A1(n_716),
.A2(n_688),
.B1(n_686),
.B2(n_693),
.C(n_478),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_721),
.B(n_734),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_713),
.B(n_705),
.C(n_724),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_711),
.A2(n_688),
.B1(n_686),
.B2(n_704),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_712),
.B(n_693),
.Y(n_754)
);

OAI21xp33_ASAP7_75t_SL g755 ( 
.A1(n_733),
.A2(n_668),
.B(n_511),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_711),
.A2(n_720),
.B1(n_709),
.B2(n_724),
.Y(n_756)
);

OAI221xp5_ASAP7_75t_L g757 ( 
.A1(n_727),
.A2(n_478),
.B1(n_473),
.B2(n_511),
.C(n_74),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_735),
.B(n_68),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_722),
.B(n_69),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_718),
.B(n_511),
.C(n_473),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_741),
.B(n_71),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_742),
.B(n_75),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_730),
.B(n_76),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_710),
.B(n_77),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_719),
.B(n_78),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_728),
.B(n_473),
.C(n_80),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_728),
.B(n_473),
.C(n_83),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_79),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_754),
.B(n_714),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_752),
.B(n_717),
.C(n_714),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_743),
.B(n_729),
.C(n_739),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_751),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_747),
.B(n_723),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_749),
.B(n_738),
.C(n_731),
.Y(n_774)
);

OAI211xp5_ASAP7_75t_SL g775 ( 
.A1(n_748),
.A2(n_740),
.B(n_732),
.C(n_726),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_746),
.B(n_740),
.Y(n_776)
);

AO21x2_ASAP7_75t_L g777 ( 
.A1(n_760),
.A2(n_737),
.B(n_86),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_745),
.Y(n_779)
);

AO21x2_ASAP7_75t_L g780 ( 
.A1(n_758),
.A2(n_84),
.B(n_88),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_745),
.B(n_90),
.Y(n_781)
);

NOR2x1_ASAP7_75t_R g782 ( 
.A(n_762),
.B(n_92),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_759),
.B(n_93),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_778),
.B(n_756),
.Y(n_784)
);

AND4x2_ASAP7_75t_L g785 ( 
.A(n_773),
.B(n_755),
.C(n_750),
.D(n_756),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_772),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_779),
.B(n_761),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_769),
.B(n_753),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_769),
.B(n_753),
.Y(n_789)
);

NAND4xp75_ASAP7_75t_L g790 ( 
.A(n_781),
.B(n_768),
.C(n_763),
.D(n_764),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_781),
.Y(n_791)
);

AO22x2_ASAP7_75t_L g792 ( 
.A1(n_770),
.A2(n_767),
.B1(n_766),
.B2(n_765),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_782),
.B(n_757),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_773),
.B(n_94),
.Y(n_794)
);

AOI22x1_ASAP7_75t_SL g795 ( 
.A1(n_785),
.A2(n_774),
.B1(n_771),
.B2(n_775),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_784),
.B(n_776),
.Y(n_796)
);

XNOR2xp5_ASAP7_75t_L g797 ( 
.A(n_790),
.B(n_783),
.Y(n_797)
);

XOR2x2_ASAP7_75t_L g798 ( 
.A(n_793),
.B(n_788),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_786),
.B(n_791),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_795),
.A2(n_787),
.B1(n_789),
.B2(n_792),
.Y(n_800)
);

OA22x2_ASAP7_75t_L g801 ( 
.A1(n_797),
.A2(n_783),
.B1(n_792),
.B2(n_794),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_799),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_796),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_798),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_804),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_802),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_800),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_803),
.Y(n_808)
);

AND4x1_ASAP7_75t_L g809 ( 
.A(n_807),
.B(n_794),
.C(n_800),
.D(n_801),
.Y(n_809)
);

AOI31xp33_ASAP7_75t_L g810 ( 
.A1(n_807),
.A2(n_805),
.A3(n_806),
.B(n_808),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_807),
.A2(n_780),
.B1(n_777),
.B2(n_104),
.Y(n_811)
);

OAI31xp33_ASAP7_75t_L g812 ( 
.A1(n_807),
.A2(n_780),
.A3(n_777),
.B(n_105),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_812),
.A2(n_193),
.B1(n_103),
.B2(n_108),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_810),
.A2(n_101),
.B1(n_109),
.B2(n_110),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_SL g815 ( 
.A1(n_809),
.A2(n_111),
.B(n_113),
.C(n_114),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_811),
.Y(n_816)
);

INVxp33_ASAP7_75t_SL g817 ( 
.A(n_814),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_816),
.Y(n_818)
);

NOR4xp25_ASAP7_75t_L g819 ( 
.A(n_813),
.B(n_116),
.C(n_118),
.D(n_120),
.Y(n_819)
);

NOR2x1_ASAP7_75t_L g820 ( 
.A(n_815),
.B(n_124),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_814),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_816),
.B(n_125),
.Y(n_822)
);

NOR2x1_ASAP7_75t_L g823 ( 
.A(n_814),
.B(n_126),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_818),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_823),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_820),
.A2(n_127),
.B1(n_130),
.B2(n_132),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_822),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_821),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_817),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_819),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_818),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_828),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_829),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_824),
.B(n_135),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_825),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_831),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_827),
.Y(n_837)
);

AND4x1_ASAP7_75t_L g838 ( 
.A(n_826),
.B(n_136),
.C(n_137),
.D(n_140),
.Y(n_838)
);

AO22x2_ASAP7_75t_L g839 ( 
.A1(n_830),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_830),
.A2(n_144),
.B(n_148),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_836),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_835),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_833),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_832),
.B(n_150),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_837),
.Y(n_845)
);

OA22x2_ASAP7_75t_L g846 ( 
.A1(n_834),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_834),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_839),
.Y(n_848)
);

AO22x2_ASAP7_75t_L g849 ( 
.A1(n_848),
.A2(n_840),
.B1(n_838),
.B2(n_158),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_841),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_841),
.Y(n_851)
);

AO22x2_ASAP7_75t_L g852 ( 
.A1(n_842),
.A2(n_191),
.B1(n_156),
.B2(n_159),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_843),
.A2(n_155),
.B1(n_160),
.B2(n_161),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_846),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_850),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_851),
.Y(n_856)
);

OR2x2_ASAP7_75t_SL g857 ( 
.A(n_854),
.B(n_847),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_849),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_858),
.A2(n_845),
.B1(n_844),
.B2(n_852),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_855),
.A2(n_853),
.B1(n_165),
.B2(n_167),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_857),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_859),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_862),
.A2(n_861),
.B1(n_856),
.B2(n_860),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_863),
.Y(n_864)
);

AOI221xp5_ASAP7_75t_L g865 ( 
.A1(n_864),
.A2(n_170),
.B1(n_171),
.B2(n_175),
.C(n_176),
.Y(n_865)
);

AOI211xp5_ASAP7_75t_L g866 ( 
.A1(n_865),
.A2(n_179),
.B(n_180),
.C(n_182),
.Y(n_866)
);


endmodule