module real_aes_8554_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_691;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_0), .A2(n_129), .B1(n_506), .B2(n_509), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_1), .A2(n_64), .B1(n_416), .B2(n_520), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_2), .A2(n_43), .B1(n_260), .B2(n_665), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_3), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_4), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_5), .A2(n_213), .B1(n_471), .B2(n_472), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_6), .A2(n_85), .B1(n_380), .B2(n_504), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_7), .A2(n_29), .B1(n_378), .B2(n_380), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_8), .A2(n_100), .B1(n_260), .B2(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_9), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_10), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_11), .A2(n_39), .B1(n_474), .B2(n_519), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_12), .A2(n_101), .B1(n_456), .B2(n_490), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_13), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_14), .A2(n_220), .B1(n_261), .B2(n_504), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_15), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_16), .A2(n_179), .B1(n_416), .B2(n_419), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_17), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_18), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_19), .A2(n_119), .B1(n_530), .B2(n_577), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_20), .Y(n_648) );
AOI22x1_ASAP7_75t_L g236 ( .A1(n_21), .A2(n_237), .B1(n_342), .B2(n_343), .Y(n_236) );
INVx1_ASAP7_75t_L g342 ( .A(n_21), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_22), .A2(n_168), .B1(n_319), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_23), .A2(n_215), .B1(n_631), .B2(n_694), .Y(n_693) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_24), .A2(n_76), .B1(n_246), .B2(n_251), .Y(n_254) );
INVx1_ASAP7_75t_L g680 ( .A(n_24), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_25), .A2(n_56), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_26), .A2(n_194), .B1(n_260), .B2(n_665), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_27), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_28), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_30), .A2(n_209), .B1(n_380), .B2(n_412), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_31), .A2(n_109), .B1(n_432), .B2(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_32), .A2(n_41), .B1(n_278), .B2(n_508), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_33), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_34), .A2(n_159), .B1(n_370), .B2(n_372), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_35), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_36), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_37), .A2(n_83), .B1(n_372), .B2(n_509), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_38), .A2(n_131), .B1(n_261), .B2(n_639), .Y(n_638) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_40), .A2(n_77), .B1(n_246), .B2(n_247), .Y(n_256) );
INVx1_ASAP7_75t_L g681 ( .A(n_40), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g374 ( .A1(n_42), .A2(n_82), .B1(n_260), .B2(n_375), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_44), .Y(n_575) );
INVx1_ASAP7_75t_L g604 ( .A(n_45), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_46), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_47), .B(n_459), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_48), .A2(n_167), .B1(n_289), .B2(n_432), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_49), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_50), .A2(n_75), .B1(n_267), .B2(n_410), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_51), .A2(n_91), .B1(n_241), .B2(n_271), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_52), .A2(n_182), .B1(n_325), .B2(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_53), .A2(n_184), .B1(n_471), .B2(n_472), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_54), .A2(n_104), .B1(n_265), .B2(n_270), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_55), .A2(n_68), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_57), .A2(n_143), .B1(n_364), .B2(n_631), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_58), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_59), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_60), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_61), .A2(n_108), .B1(n_312), .B2(n_447), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_62), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_63), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_65), .A2(n_176), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_66), .A2(n_174), .B1(n_359), .B2(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_67), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_69), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_70), .A2(n_84), .B1(n_292), .B2(n_561), .Y(n_601) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_71), .A2(n_130), .B1(n_139), .B2(n_456), .C1(n_700), .C2(n_701), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_72), .A2(n_147), .B1(n_383), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_73), .A2(n_155), .B1(n_416), .B2(n_436), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_74), .A2(n_120), .B1(n_366), .B2(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_78), .A2(n_207), .B1(n_364), .B2(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_79), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g229 ( .A(n_80), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_81), .A2(n_158), .B1(n_561), .B2(n_562), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_86), .A2(n_157), .B1(n_288), .B2(n_292), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_87), .Y(n_385) );
INVx1_ASAP7_75t_L g226 ( .A(n_88), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_89), .A2(n_144), .B1(n_410), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_90), .A2(n_107), .B1(n_326), .B2(n_365), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_92), .A2(n_121), .B1(n_278), .B2(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_93), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_94), .A2(n_156), .B1(n_384), .B2(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_95), .A2(n_187), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_96), .A2(n_196), .B1(n_584), .B2(n_585), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_97), .A2(n_211), .B1(n_326), .B2(n_352), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_98), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_99), .B(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_102), .A2(n_105), .B1(n_372), .B2(n_688), .Y(n_687) );
OA22x2_ASAP7_75t_L g391 ( .A1(n_103), .A2(n_392), .B1(n_393), .B2(n_420), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_103), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_106), .A2(n_137), .B1(n_375), .B2(n_721), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g729 ( .A1(n_110), .A2(n_138), .B1(n_163), .B2(n_320), .C1(n_463), .C2(n_701), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_111), .B(n_356), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_112), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_113), .Y(n_438) );
XNOR2x2_ASAP7_75t_L g554 ( .A(n_114), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_115), .B(n_488), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_116), .A2(n_186), .B1(n_436), .B2(n_502), .Y(n_540) );
INVx2_ASAP7_75t_L g230 ( .A(n_117), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_118), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_122), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_123), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_124), .A2(n_197), .B1(n_456), .B2(n_581), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_125), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_126), .Y(n_494) );
AND2x6_ASAP7_75t_L g225 ( .A(n_127), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_127), .Y(n_674) );
AO22x2_ASAP7_75t_L g245 ( .A1(n_128), .A2(n_177), .B1(n_246), .B2(n_247), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_132), .A2(n_192), .B1(n_491), .B2(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_133), .B(n_585), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_134), .A2(n_204), .B1(n_289), .B2(n_416), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_135), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_136), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_140), .A2(n_165), .B1(n_412), .B2(n_413), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_141), .A2(n_216), .B1(n_410), .B2(n_419), .Y(n_727) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_142), .A2(n_223), .B(n_231), .C(n_682), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_145), .A2(n_152), .B1(n_366), .B2(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_146), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_148), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_149), .A2(n_221), .B1(n_265), .B2(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_150), .A2(n_170), .B1(n_490), .B2(n_491), .Y(n_489) );
AO22x2_ASAP7_75t_L g250 ( .A1(n_151), .A2(n_198), .B1(n_246), .B2(n_251), .Y(n_250) );
INVxp67_ASAP7_75t_L g713 ( .A(n_153), .Y(n_713) );
XOR2x2_ASAP7_75t_L g715 ( .A(n_153), .B(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_154), .A2(n_590), .B1(n_618), .B2(n_619), .Y(n_589) );
INVx1_ASAP7_75t_L g618 ( .A(n_154), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_160), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_161), .A2(n_188), .B1(n_383), .B2(n_384), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_162), .A2(n_178), .B1(n_352), .B2(n_447), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_164), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_166), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_169), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_171), .B(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_172), .A2(n_206), .B1(n_325), .B2(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_173), .B(n_359), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_175), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_177), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_180), .B(n_613), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_181), .Y(n_328) );
INVx1_ASAP7_75t_L g425 ( .A(n_183), .Y(n_425) );
INVx1_ASAP7_75t_L g666 ( .A(n_185), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_189), .Y(n_476) );
OA22x2_ASAP7_75t_L g521 ( .A1(n_190), .A2(n_522), .B1(n_523), .B2(n_546), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_190), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_191), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_193), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_195), .A2(n_203), .B1(n_688), .B2(n_697), .Y(n_728) );
INVx1_ASAP7_75t_L g677 ( .A(n_198), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_199), .Y(n_350) );
AOI211xp5_ASAP7_75t_L g482 ( .A1(n_200), .A2(n_444), .B(n_483), .C(n_493), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_201), .A2(n_219), .B1(n_359), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_202), .A2(n_205), .B1(n_260), .B2(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g246 ( .A(n_208), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_210), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_212), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_214), .A2(n_684), .B1(n_702), .B2(n_703), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_214), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_217), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_218), .Y(n_655) );
INVx2_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_226), .Y(n_673) );
OA21x2_ASAP7_75t_L g711 ( .A1(n_227), .A2(n_672), .B(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_552), .B1(n_667), .B2(n_668), .C(n_669), .Y(n_231) );
INVx1_ASAP7_75t_L g667 ( .A(n_232), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B1(n_387), .B2(n_551), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_236), .B1(n_344), .B2(n_386), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_SL g343 ( .A(n_237), .Y(n_343) );
AND2x2_ASAP7_75t_SL g237 ( .A(n_238), .B(n_296), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_275), .Y(n_238) );
OAI221xp5_ASAP7_75t_SL g239 ( .A1(n_240), .A2(n_257), .B1(n_258), .B2(n_263), .C(n_264), .Y(n_239) );
INVx2_ASAP7_75t_L g502 ( .A(n_240), .Y(n_502) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_241), .Y(n_559) );
BUFx3_ASAP7_75t_L g599 ( .A(n_241), .Y(n_599) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_242), .Y(n_383) );
INVx2_ASAP7_75t_L g417 ( .A(n_242), .Y(n_417) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
AND2x6_ASAP7_75t_L g267 ( .A(n_243), .B(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g278 ( .A(n_243), .B(n_279), .Y(n_278) );
AND2x6_ASAP7_75t_L g320 ( .A(n_243), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_249), .Y(n_243) );
AND2x2_ASAP7_75t_L g262 ( .A(n_244), .B(n_250), .Y(n_262) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_245), .B(n_250), .Y(n_274) );
AND2x2_ASAP7_75t_L g284 ( .A(n_245), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g316 ( .A(n_245), .B(n_254), .Y(n_316) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g251 ( .A(n_248), .Y(n_251) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
INVx1_ASAP7_75t_L g315 ( .A(n_250), .Y(n_315) );
AND2x4_ASAP7_75t_L g261 ( .A(n_252), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g272 ( .A(n_252), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_252), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g381 ( .A(n_252), .B(n_284), .Y(n_381) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
OR2x2_ASAP7_75t_L g269 ( .A(n_253), .B(n_256), .Y(n_269) );
AND2x2_ASAP7_75t_L g279 ( .A(n_253), .B(n_256), .Y(n_279) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g321 ( .A(n_254), .B(n_256), .Y(n_321) );
AND2x2_ASAP7_75t_L g314 ( .A(n_255), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g295 ( .A(n_256), .Y(n_295) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g475 ( .A(n_261), .Y(n_475) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_261), .Y(n_568) );
INVx1_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_262), .B(n_279), .Y(n_308) );
AND2x6_ASAP7_75t_L g357 ( .A(n_262), .B(n_279), .Y(n_357) );
AND2x4_ASAP7_75t_L g362 ( .A(n_262), .B(n_268), .Y(n_362) );
INVx4_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx5_ASAP7_75t_SL g504 ( .A(n_266), .Y(n_504) );
INVx1_ASAP7_75t_L g697 ( .A(n_266), .Y(n_697) );
INVx11_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx11_ASAP7_75t_L g379 ( .A(n_267), .Y(n_379) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g302 ( .A(n_269), .B(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_SL g384 ( .A(n_272), .Y(n_384) );
BUFx3_ASAP7_75t_L g419 ( .A(n_272), .Y(n_419) );
BUFx2_ASAP7_75t_L g436 ( .A(n_272), .Y(n_436) );
BUFx3_ASAP7_75t_L g520 ( .A(n_272), .Y(n_520) );
AND2x2_ASAP7_75t_L g432 ( .A(n_273), .B(n_334), .Y(n_432) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x6_ASAP7_75t_L g294 ( .A(n_274), .B(n_295), .Y(n_294) );
OAI221xp5_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_280), .B1(n_281), .B2(n_286), .C(n_287), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx6_ASAP7_75t_L g371 ( .A(n_278), .Y(n_371) );
BUFx3_ASAP7_75t_L g412 ( .A(n_278), .Y(n_412) );
BUFx3_ASAP7_75t_L g594 ( .A(n_278), .Y(n_594) );
AND2x2_ASAP7_75t_L g291 ( .A(n_279), .B(n_284), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_281), .A2(n_371), .B1(n_570), .B2(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g514 ( .A(n_282), .Y(n_514) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g341 ( .A(n_285), .Y(n_341) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_289), .Y(n_721) );
INVx5_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx3_ASAP7_75t_L g373 ( .A(n_290), .Y(n_373) );
INVx3_ASAP7_75t_L g472 ( .A(n_290), .Y(n_472) );
INVx4_ASAP7_75t_L g508 ( .A(n_290), .Y(n_508) );
INVx8_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx4f_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g375 ( .A(n_293), .Y(n_375) );
BUFx2_ASAP7_75t_L g562 ( .A(n_293), .Y(n_562) );
BUFx2_ASAP7_75t_L g665 ( .A(n_293), .Y(n_665) );
INVx6_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_294), .A2(n_338), .B1(n_405), .B2(n_406), .Y(n_404) );
INVx1_ASAP7_75t_SL g509 ( .A(n_294), .Y(n_509) );
INVx1_ASAP7_75t_SL g639 ( .A(n_294), .Y(n_639) );
INVx1_ASAP7_75t_L g367 ( .A(n_295), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_309), .C(n_329), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_304), .B2(n_305), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g397 ( .A(n_302), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_302), .A2(n_307), .B1(n_438), .B2(n_439), .C(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g606 ( .A(n_302), .Y(n_606) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g485 ( .A(n_307), .Y(n_485) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g400 ( .A(n_308), .Y(n_400) );
OAI222xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_317), .B1(n_318), .B2(n_322), .C1(n_323), .C2(n_328), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_310), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_310), .A2(n_609), .B1(n_610), .B2(n_611), .C(n_612), .Y(n_608) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g656 ( .A(n_311), .Y(n_656) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
BUFx2_ASAP7_75t_L g413 ( .A(n_313), .Y(n_413) );
BUFx4f_ASAP7_75t_SL g463 ( .A(n_313), .Y(n_463) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_313), .Y(n_694) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
AND2x4_ASAP7_75t_L g326 ( .A(n_316), .B(n_327), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_316), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g366 ( .A(n_316), .B(n_367), .Y(n_366) );
OAI222xp33_ASAP7_75t_L g525 ( .A1(n_318), .A2(n_526), .B1(n_527), .B2(n_528), .C1(n_529), .C2(n_532), .Y(n_525) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g454 ( .A(n_319), .Y(n_454) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
BUFx3_ASAP7_75t_L g444 ( .A(n_320), .Y(n_444) );
INVx2_ASAP7_75t_L g574 ( .A(n_320), .Y(n_574) );
INVx2_ASAP7_75t_SL g609 ( .A(n_320), .Y(n_609) );
INVx4_ASAP7_75t_L g651 ( .A(n_320), .Y(n_651) );
INVx1_ASAP7_75t_L g339 ( .A(n_321), .Y(n_339) );
AND2x4_ASAP7_75t_L g353 ( .A(n_321), .B(n_341), .Y(n_353) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g614 ( .A(n_325), .Y(n_614) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx12f_ASAP7_75t_L g447 ( .A(n_326), .Y(n_447) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_326), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_335), .B2(n_336), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_331), .A2(n_336), .B1(n_616), .B2(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_333), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_338), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g386 ( .A(n_344), .Y(n_386) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
XOR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_385), .Y(n_345) );
NAND3x1_ASAP7_75t_L g346 ( .A(n_347), .B(n_368), .C(n_376), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_354), .Y(n_347) );
OAI21xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_350), .B(n_351), .Y(n_348) );
BUFx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_353), .Y(n_441) );
BUFx2_ASAP7_75t_SL g456 ( .A(n_353), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .C(n_363), .Y(n_354) );
BUFx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx4f_ASAP7_75t_L g461 ( .A(n_357), .Y(n_461) );
INVx1_ASAP7_75t_SL g537 ( .A(n_357), .Y(n_537) );
BUFx2_ASAP7_75t_L g585 ( .A(n_357), .Y(n_585) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g459 ( .A(n_361), .Y(n_459) );
INVx2_ASAP7_75t_L g488 ( .A(n_361), .Y(n_488) );
INVx2_ASAP7_75t_L g584 ( .A(n_361), .Y(n_584) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g526 ( .A(n_364), .Y(n_526) );
INVx4_ASAP7_75t_L g578 ( .A(n_364), .Y(n_578) );
BUFx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g490 ( .A(n_366), .Y(n_490) );
INVx1_ASAP7_75t_L g582 ( .A(n_366), .Y(n_582) );
BUFx3_ASAP7_75t_L g631 ( .A(n_366), .Y(n_631) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_374), .Y(n_368) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g471 ( .A(n_371), .Y(n_471) );
INVx2_ASAP7_75t_L g688 ( .A(n_371), .Y(n_688) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_382), .Y(n_376) );
INVx4_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp33_ASAP7_75t_SL g401 ( .A1(n_379), .A2(n_402), .B(n_403), .Y(n_401) );
INVx4_ASAP7_75t_L g430 ( .A(n_379), .Y(n_430) );
INVx3_ASAP7_75t_L g600 ( .A(n_379), .Y(n_600) );
BUFx3_ASAP7_75t_L g545 ( .A(n_380), .Y(n_545) );
BUFx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
BUFx3_ASAP7_75t_L g467 ( .A(n_381), .Y(n_467) );
INVx1_ASAP7_75t_L g551 ( .A(n_387), .Y(n_551) );
XNOR2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_421), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g420 ( .A(n_393), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_407), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_401), .C(n_404), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_397), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_399), .A2(n_604), .B1(n_605), .B2(n_607), .Y(n_603) );
OA211x2_ASAP7_75t_L g690 ( .A1(n_399), .A2(n_691), .B(n_692), .C(n_693), .Y(n_690) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g649 ( .A(n_400), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_414), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
BUFx2_ASAP7_75t_L g595 ( .A(n_410), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g429 ( .A(n_417), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_478), .B1(n_549), .B2(n_550), .Y(n_421) );
INVx1_ASAP7_75t_L g549 ( .A(n_422), .Y(n_549) );
OAI22xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .B1(n_448), .B2(n_477), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
XNOR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NOR4xp75_ASAP7_75t_L g426 ( .A(n_427), .B(n_433), .C(n_437), .D(n_442), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_431), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_SL g492 ( .A(n_441), .Y(n_492) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_445), .B(n_446), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
BUFx4f_ASAP7_75t_SL g701 ( .A(n_447), .Y(n_701) );
INVx2_ASAP7_75t_SL g477 ( .A(n_448), .Y(n_477) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
XOR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_476), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_464), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_457), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_455), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .C(n_462), .Y(n_457) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
INVxp67_ASAP7_75t_L g512 ( .A(n_471), .Y(n_512) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_475), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_515) );
INVx1_ASAP7_75t_L g550 ( .A(n_478), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_521), .B1(n_547), .B2(n_548), .Y(n_478) );
INVx2_ASAP7_75t_L g548 ( .A(n_479), .Y(n_548) );
XNOR2x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_499), .Y(n_481) );
OAI211xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B(n_486), .C(n_489), .Y(n_483) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .C(n_515), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g565 ( .A(n_504), .Y(n_565) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_508), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_510) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g547 ( .A(n_521), .Y(n_547) );
INVx1_ASAP7_75t_SL g546 ( .A(n_523), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_538), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_533), .Y(n_524) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_SL g724 ( .A(n_537), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g668 ( .A(n_552), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_643), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_586), .B1(n_587), .B2(n_642), .Y(n_553) );
INVx2_ASAP7_75t_L g642 ( .A(n_554), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_556), .B(n_572), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_563), .C(n_569), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_563) );
INVx4_ASAP7_75t_L g719 ( .A(n_567), .Y(n_719) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_579), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_575), .B(n_576), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_574), .A2(n_625), .B(n_626), .Y(n_624) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_620), .B1(n_621), .B2(n_641), .Y(n_587) );
INVx2_ASAP7_75t_L g641 ( .A(n_588), .Y(n_641) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g619 ( .A(n_590), .Y(n_619) );
AND2x2_ASAP7_75t_SL g590 ( .A(n_591), .B(n_602), .Y(n_590) );
NOR2xp33_ASAP7_75t_SL g591 ( .A(n_592), .B(n_597), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_608), .C(n_615), .Y(n_602) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
XOR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .Y(n_621) );
NAND2x1_ASAP7_75t_SL g622 ( .A(n_623), .B(n_632), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .C(n_630), .Y(n_627) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_636), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_666), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_658), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_650), .C(n_654), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_653), .Y(n_650) );
INVx4_ASAP7_75t_L g700 ( .A(n_651), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
OR2x2_ASAP7_75t_SL g732 ( .A(n_671), .B(n_676), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_672), .Y(n_705) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_673), .B(n_708), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g708 ( .A(n_674), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_704), .A3(n_706), .B1(n_709), .B2(n_713), .C1(n_714), .C2(n_730), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_684), .Y(n_703) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND4xp75_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .C(n_695), .D(n_699), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_710), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND4xp75_ASAP7_75t_L g716 ( .A(n_717), .B(n_722), .C(n_726), .D(n_729), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
AND2x2_ASAP7_75t_SL g722 ( .A(n_723), .B(n_725), .Y(n_722) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
endmodule