module fake_jpeg_4842_n_96 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_27),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_16),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_43)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_6),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_15),
.C(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_53),
.Y(n_65)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_21),
.C(n_12),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_36),
.C(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_49),
.B1(n_45),
.B2(n_40),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_17),
.B(n_20),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_46),
.B(n_52),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_17),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_11),
.B1(n_44),
.B2(n_45),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_64),
.B1(n_62),
.B2(n_57),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_50),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_34),
.C(n_49),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_76),
.C(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_52),
.B(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_71),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_75),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_51),
.C(n_42),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_69),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_59),
.C(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_83),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_76),
.B(n_66),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_88),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_69),
.B1(n_73),
.B2(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_81),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_91),
.B1(n_77),
.B2(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_37),
.Y(n_94)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_63),
.C(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_63),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);


endmodule