module fake_jpeg_29807_n_33 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_2),
.A2(n_5),
.B1(n_12),
.B2(n_6),
.Y(n_14)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_3),
.B1(n_6),
.B2(n_13),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_9),
.B(n_10),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_22),
.B(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_1),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_17),
.C(n_4),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_17),
.C(n_4),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_3),
.C(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_24),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_25),
.B(n_31),
.Y(n_33)
);


endmodule