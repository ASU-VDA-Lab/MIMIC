module fake_jpeg_27454_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_68),
.Y(n_72)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_48),
.Y(n_71)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_58),
.B1(n_52),
.B2(n_49),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_53),
.B1(n_32),
.B2(n_24),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_97),
.Y(n_107)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_90),
.B1(n_98),
.B2(n_66),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_92),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_31),
.B1(n_32),
.B2(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_77),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_38),
.B1(n_31),
.B2(n_40),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_89),
.B1(n_76),
.B2(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_40),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_105),
.B1(n_116),
.B2(n_22),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_38),
.B1(n_56),
.B2(n_66),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_78),
.B1(n_75),
.B2(n_69),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_31),
.B(n_66),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_113),
.B(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_29),
.B1(n_27),
.B2(n_17),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_56),
.B1(n_67),
.B2(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_47),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_47),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_56),
.B1(n_53),
.B2(n_59),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_67),
.C(n_47),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_46),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_67),
.B1(n_46),
.B2(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_93),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_1),
.B(n_2),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_130),
.B1(n_142),
.B2(n_147),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_75),
.B1(n_78),
.B2(n_98),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_21),
.C(n_19),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_138),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_62),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_143),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_152),
.B1(n_23),
.B2(n_17),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_102),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_155),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_61),
.B(n_80),
.C(n_93),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_88),
.B(n_81),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_69),
.B1(n_22),
.B2(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_150),
.B1(n_25),
.B2(n_30),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_115),
.B(n_103),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_18),
.B1(n_91),
.B2(n_35),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_154),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_25),
.B1(n_17),
.B2(n_30),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_25),
.B1(n_30),
.B2(n_35),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_46),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_120),
.B1(n_112),
.B2(n_125),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_159),
.B1(n_161),
.B2(n_169),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_157),
.A2(n_171),
.B(n_179),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_115),
.B(n_109),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_158),
.A2(n_147),
.B(n_150),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_119),
.B1(n_100),
.B2(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_108),
.B1(n_110),
.B2(n_116),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_181),
.B1(n_185),
.B2(n_151),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_168),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_43),
.C(n_23),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_11),
.C(n_16),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_110),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_167),
.B(n_177),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_118),
.C(n_81),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_146),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_154),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_91),
.B1(n_35),
.B2(n_88),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_36),
.B1(n_34),
.B2(n_28),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_36),
.B1(n_34),
.B2(n_28),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_188),
.B1(n_128),
.B2(n_141),
.Y(n_216)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_149),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_36),
.B1(n_34),
.B2(n_28),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_189),
.B(n_173),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_216),
.B1(n_157),
.B2(n_158),
.Y(n_221)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_198),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_127),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_196),
.B(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_200),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_144),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_144),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_203),
.B(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_139),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_132),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_179),
.B(n_175),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_188),
.B1(n_186),
.B2(n_166),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_156),
.A2(n_131),
.B1(n_149),
.B2(n_114),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_187),
.B1(n_173),
.B2(n_182),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_210),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_242),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_236),
.B1(n_216),
.B2(n_200),
.Y(n_258)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_233),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_179),
.B(n_178),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_231),
.B(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_204),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_167),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_193),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_177),
.C(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_245),
.C(n_192),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_36),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_26),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_21),
.C(n_26),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_215),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_182),
.C(n_114),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_252),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_217),
.B1(n_206),
.B2(n_201),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_248),
.A2(n_251),
.B1(n_255),
.B2(n_233),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_257),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_193),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_198),
.B1(n_194),
.B2(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_265),
.B1(n_222),
.B2(n_225),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_114),
.C(n_21),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_34),
.C(n_26),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_26),
.C(n_16),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_267),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_236),
.B1(n_227),
.B2(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_275),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_244),
.B(n_241),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_278),
.B(n_284),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_231),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_281),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_252),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_220),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_261),
.C(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_276),
.B(n_249),
.C(n_237),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_296),
.B1(n_291),
.B2(n_298),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_269),
.C(n_271),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_230),
.B1(n_228),
.B2(n_265),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_296),
.B1(n_277),
.B2(n_285),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_230),
.B1(n_224),
.B2(n_239),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_298),
.B1(n_4),
.B2(n_5),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_223),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_5),
.B(n_6),
.Y(n_313)
);

OAI221xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_243),
.B1(n_240),
.B2(n_261),
.C(n_263),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_295),
.B(n_299),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_254),
.B(n_259),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_9),
.B(n_14),
.C(n_12),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_274),
.C(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_304),
.C(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_274),
.C(n_281),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_5),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_16),
.B(n_12),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_12),
.C(n_11),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_7),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_9),
.B(n_6),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_292),
.B1(n_299),
.B2(n_288),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_8),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_317),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_307),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_310),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_7),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_321),
.B(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_316),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_301),
.C(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_315),
.C(n_323),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_309),
.B(n_303),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_333),
.C(n_328),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_332),
.B1(n_325),
.B2(n_330),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_322),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_326),
.C(n_7),
.Y(n_338)
);

OAI21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_7),
.B(n_8),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_8),
.B(n_253),
.Y(n_340)
);


endmodule