module fake_jpeg_2451_n_617 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_617);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_617;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_63),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_64),
.Y(n_220)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_66),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_67),
.B(n_70),
.Y(n_147)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_71),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_11),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_77),
.Y(n_163)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_76),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_10),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_78),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_79),
.B(n_89),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_12),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_80),
.B(n_124),
.Y(n_167)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_83),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_41),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_84),
.B(n_19),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_87),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_96),
.B(n_102),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_55),
.Y(n_100)
);

CKINVDCx9p33_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_101),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_28),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_40),
.A2(n_9),
.B(n_18),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_57),
.B(n_48),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_26),
.B(n_9),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_112),
.B(n_125),
.Y(n_218)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_120),
.B(n_121),
.Y(n_203)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_56),
.A2(n_13),
.B(n_18),
.Y(n_123)
);

HAxp5_ASAP7_75t_SL g209 ( 
.A(n_123),
.B(n_0),
.CON(n_209),
.SN(n_209)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_28),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_31),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

CKINVDCx10_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_36),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_33),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_56),
.C(n_49),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_130),
.B(n_159),
.C(n_201),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_137),
.A2(n_171),
.B(n_196),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_46),
.B1(n_53),
.B2(n_43),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_148),
.A2(n_153),
.B1(n_161),
.B2(n_166),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_61),
.A2(n_46),
.B1(n_53),
.B2(n_43),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_149),
.A2(n_157),
.B1(n_191),
.B2(n_214),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_76),
.A2(n_49),
.B1(n_50),
.B2(n_37),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_72),
.A2(n_50),
.B1(n_52),
.B2(n_57),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_118),
.B(n_57),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_158),
.B(n_179),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_62),
.B(n_91),
.C(n_103),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_73),
.A2(n_78),
.B1(n_83),
.B2(n_110),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_52),
.B1(n_48),
.B2(n_45),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_48),
.B1(n_45),
.B2(n_44),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_170),
.A2(n_200),
.B1(n_2),
.B2(n_207),
.Y(n_236)
);

OR2x2_ASAP7_75t_SL g171 ( 
.A(n_63),
.B(n_45),
.Y(n_171)
);

CKINVDCx12_ASAP7_75t_R g172 ( 
.A(n_64),
.Y(n_172)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_172),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_173),
.Y(n_294)
);

BUFx16f_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_177),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_180),
.B(n_181),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_44),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_44),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_187),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_85),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_184),
.A2(n_186),
.B1(n_145),
.B2(n_160),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_99),
.A2(n_37),
.B1(n_33),
.B2(n_52),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_59),
.B(n_37),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_97),
.B(n_33),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_189),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_97),
.B(n_0),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_190),
.B(n_210),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_81),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_58),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_66),
.A2(n_6),
.B1(n_16),
.B2(n_15),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_223),
.B1(n_95),
.B2(n_1),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_127),
.A2(n_6),
.B1(n_16),
.B2(n_15),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_2),
.B1(n_130),
.B2(n_135),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_209),
.A2(n_176),
.B(n_140),
.C(n_194),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_59),
.B(n_4),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_194),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_117),
.B(n_4),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_122),
.B(n_3),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_94),
.A2(n_3),
.B1(n_13),
.B2(n_14),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_126),
.B(n_3),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_178),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_226),
.B(n_237),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_227),
.A2(n_236),
.B1(n_247),
.B2(n_253),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_64),
.B1(n_3),
.B2(n_19),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_228),
.A2(n_254),
.B1(n_275),
.B2(n_283),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_0),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_229),
.B(n_231),
.Y(n_311)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_230),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_0),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_1),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_233),
.B(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_234),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_171),
.A2(n_2),
.B(n_196),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_235),
.A2(n_279),
.B(n_244),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_155),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_238),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_239),
.A2(n_293),
.B1(n_295),
.B2(n_298),
.Y(n_308)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_241),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_143),
.Y(n_242)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_242),
.Y(n_342)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_243),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_244),
.B(n_250),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_167),
.A2(n_2),
.B(n_163),
.C(n_215),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_246),
.A2(n_281),
.B(n_235),
.C(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_251),
.B(n_261),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_252),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_216),
.B1(n_222),
.B2(n_174),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_154),
.A2(n_147),
.B1(n_159),
.B2(n_164),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_189),
.B(n_152),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_131),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_258),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_267),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_263),
.B(n_274),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_197),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_164),
.B(n_168),
.C(n_131),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_265),
.B(n_287),
.C(n_285),
.Y(n_329)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_266),
.B(n_269),
.Y(n_353)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_133),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_134),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_268),
.B(n_277),
.Y(n_348)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_168),
.B(n_165),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_271),
.B(n_300),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_134),
.B(n_186),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_288),
.Y(n_315)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_273),
.B(n_276),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_151),
.A2(n_162),
.B1(n_185),
.B2(n_206),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_138),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g330 ( 
.A(n_278),
.Y(n_330)
);

NAND2x1_ASAP7_75t_L g279 ( 
.A(n_209),
.B(n_142),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_141),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_280),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_176),
.A2(n_165),
.B(n_138),
.C(n_184),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_199),
.A2(n_219),
.B1(n_206),
.B2(n_143),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_284),
.B(n_241),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_151),
.B(n_162),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_285),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_199),
.A2(n_219),
.B1(n_185),
.B2(n_144),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_286),
.A2(n_299),
.B1(n_292),
.B2(n_249),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_212),
.B(n_142),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_182),
.B(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_182),
.B(n_205),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_285),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_290),
.Y(n_335)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_144),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_292),
.Y(n_358)
);

OA22x2_ASAP7_75t_L g293 ( 
.A1(n_141),
.A2(n_193),
.B1(n_139),
.B2(n_169),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_214),
.A2(n_135),
.B1(n_139),
.B2(n_169),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_297),
.A2(n_264),
.B1(n_237),
.B2(n_296),
.Y(n_357)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_193),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_198),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_299),
.A2(n_305),
.B1(n_132),
.B2(n_146),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_140),
.B(n_194),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_150),
.B(n_204),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_301),
.B(n_304),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_150),
.B(n_204),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_132),
.A2(n_204),
.B1(n_150),
.B2(n_156),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_247),
.A2(n_198),
.B1(n_156),
.B2(n_146),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_317),
.B1(n_321),
.B2(n_326),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_297),
.A2(n_272),
.B1(n_291),
.B2(n_259),
.Y(n_317)
);

BUFx4f_ASAP7_75t_SL g386 ( 
.A(n_320),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_291),
.A2(n_132),
.B1(n_274),
.B2(n_257),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_274),
.A2(n_233),
.B1(n_231),
.B2(n_229),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_327),
.B(n_328),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_258),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_263),
.B(n_260),
.CI(n_279),
.CON(n_331),
.SN(n_331)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_331),
.B(n_345),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_225),
.A2(n_253),
.B1(n_294),
.B2(n_227),
.Y(n_334)
);

OA22x2_ASAP7_75t_L g403 ( 
.A1(n_334),
.A2(n_321),
.B1(n_327),
.B2(n_331),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_232),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_337),
.C(n_351),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_246),
.B(n_248),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_303),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_293),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_270),
.B(n_289),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_288),
.A2(n_281),
.B1(n_273),
.B2(n_282),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_349),
.A2(n_243),
.B1(n_255),
.B2(n_256),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_265),
.B(n_267),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_350),
.B(n_266),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_268),
.B(n_262),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_360),
.B1(n_252),
.B2(n_269),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_356),
.A2(n_284),
.B(n_277),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_357),
.A2(n_293),
.B1(n_230),
.B2(n_250),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_280),
.A2(n_234),
.B1(n_238),
.B2(n_298),
.Y(n_360)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_365),
.B(n_394),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_366),
.A2(n_378),
.B(n_404),
.Y(n_430)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

INVx6_ASAP7_75t_SL g370 ( 
.A(n_330),
.Y(n_370)
);

INVx13_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_319),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_373),
.B(n_374),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_319),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_376),
.B(n_382),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_377),
.A2(n_330),
.B1(n_338),
.B2(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_339),
.Y(n_379)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_293),
.B(n_302),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_380),
.A2(n_384),
.B(n_385),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_381),
.B(n_388),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_240),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_383),
.A2(n_391),
.B1(n_397),
.B2(n_403),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_328),
.A2(n_302),
.B(n_245),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_328),
.A2(n_276),
.B(n_242),
.Y(n_385)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_337),
.B(n_345),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_309),
.A2(n_317),
.B1(n_315),
.B2(n_333),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_409),
.B1(n_346),
.B2(n_343),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_334),
.A2(n_309),
.B1(n_315),
.B2(n_335),
.Y(n_391)
);

OA21x2_ASAP7_75t_L g392 ( 
.A1(n_349),
.A2(n_335),
.B(n_314),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_392),
.A2(n_398),
.B(n_380),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_393),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_336),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_311),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_396),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_311),
.B(n_351),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_329),
.B1(n_333),
.B2(n_308),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_344),
.A2(n_347),
.B(n_341),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_326),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_402),
.Y(n_440)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_339),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_407),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_340),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_338),
.B(n_340),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_313),
.A2(n_316),
.B1(n_331),
.B2(n_361),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_405),
.A2(n_406),
.B1(n_394),
.B2(n_396),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_331),
.A2(n_313),
.B1(n_361),
.B2(n_316),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_330),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_352),
.A2(n_344),
.B1(n_359),
.B2(n_325),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_371),
.B1(n_400),
.B2(n_399),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_412),
.A2(n_416),
.B1(n_426),
.B2(n_438),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_371),
.A2(n_306),
.B1(n_348),
.B2(n_307),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_420),
.A2(n_432),
.B1(n_385),
.B2(n_398),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_400),
.A2(n_348),
.B(n_355),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_424),
.A2(n_439),
.B(n_366),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_425),
.B(n_441),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_306),
.B1(n_307),
.B2(n_353),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_319),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_441),
.C(n_427),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_429),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_381),
.B(n_319),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_434),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_343),
.B1(n_355),
.B2(n_358),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_310),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_370),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_362),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_395),
.A2(n_343),
.B1(n_358),
.B2(n_323),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_376),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_346),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_369),
.B(n_363),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_443),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_382),
.B(n_312),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_404),
.Y(n_444)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_446),
.A2(n_392),
.B1(n_377),
.B2(n_379),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_447),
.A2(n_386),
.B(n_318),
.Y(n_475)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_450),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_467),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_452),
.B(n_482),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_438),
.Y(n_453)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_453),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_405),
.C(n_368),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_454),
.B(n_460),
.C(n_481),
.Y(n_488)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_456),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_412),
.B(n_368),
.CI(n_375),
.CON(n_457),
.SN(n_457)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_457),
.B(n_466),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_458),
.A2(n_463),
.B(n_467),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_423),
.A2(n_439),
.B1(n_447),
.B2(n_444),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_459),
.A2(n_468),
.B1(n_469),
.B2(n_417),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_375),
.Y(n_460)
);

AOI322xp5_ASAP7_75t_L g461 ( 
.A1(n_440),
.A2(n_388),
.A3(n_397),
.B1(n_403),
.B2(n_373),
.C1(n_374),
.C2(n_408),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_433),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_439),
.A2(n_407),
.B(n_392),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_464),
.A2(n_473),
.B1(n_476),
.B2(n_479),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_354),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_447),
.A2(n_403),
.B(n_386),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_423),
.A2(n_403),
.B1(n_392),
.B2(n_383),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_420),
.A2(n_403),
.B1(n_372),
.B2(n_367),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_354),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_470),
.B(n_422),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_418),
.A2(n_401),
.B(n_387),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_471),
.A2(n_475),
.B(n_421),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_322),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_478),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_446),
.A2(n_386),
.B1(n_387),
.B2(n_364),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_364),
.Y(n_474)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_426),
.A2(n_386),
.B1(n_390),
.B2(n_362),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_318),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_416),
.A2(n_362),
.B1(n_390),
.B2(n_432),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_422),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_428),
.Y(n_481)
);

MAJx2_ASAP7_75t_L g482 ( 
.A(n_428),
.B(n_413),
.C(n_415),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_419),
.Y(n_484)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_484),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_463),
.A2(n_418),
.B(n_424),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_486),
.A2(n_499),
.B(n_508),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_490),
.A2(n_493),
.B1(n_495),
.B2(n_496),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_468),
.A2(n_435),
.B1(n_414),
.B2(n_432),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_451),
.A2(n_435),
.B1(n_414),
.B2(n_417),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_469),
.A2(n_415),
.B1(n_430),
.B2(n_431),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_459),
.A2(n_430),
.B1(n_413),
.B2(n_420),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_497),
.A2(n_498),
.B1(n_511),
.B2(n_479),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_462),
.A2(n_429),
.B1(n_443),
.B2(n_424),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_458),
.A2(n_436),
.B(n_442),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_509),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_502),
.B(n_503),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_449),
.B(n_465),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_433),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_512),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_449),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_454),
.B(n_437),
.C(n_411),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_452),
.C(n_481),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_437),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_510),
.A2(n_514),
.B(n_508),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_462),
.A2(n_445),
.B1(n_411),
.B2(n_421),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_456),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_475),
.A2(n_421),
.B(n_411),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_515),
.B(n_524),
.C(n_536),
.Y(n_542)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_486),
.B(n_482),
.CI(n_457),
.CON(n_516),
.SN(n_516)
);

MAJx2_ASAP7_75t_L g549 ( 
.A(n_516),
.B(n_526),
.C(n_528),
.Y(n_549)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_517),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_500),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_522),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_523),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_488),
.C(n_483),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_464),
.B1(n_471),
.B2(n_477),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_525),
.A2(n_531),
.B1(n_534),
.B2(n_538),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_472),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_488),
.B(n_483),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_490),
.A2(n_448),
.B1(n_476),
.B2(n_473),
.Y(n_529)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_529),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_480),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_532),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_487),
.A2(n_478),
.B1(n_456),
.B2(n_457),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_445),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_533),
.A2(n_527),
.B(n_485),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_493),
.A2(n_510),
.B1(n_498),
.B2(n_495),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_494),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_535),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_491),
.B(n_499),
.C(n_497),
.Y(n_536)
);

FAx1_ASAP7_75t_SL g538 ( 
.A(n_494),
.B(n_485),
.CI(n_496),
.CON(n_538),
.SN(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_502),
.Y(n_539)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_510),
.A2(n_500),
.B1(n_513),
.B2(n_512),
.Y(n_540)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_544),
.B(n_533),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_515),
.B(n_492),
.C(n_513),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_546),
.B(n_548),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_492),
.C(n_511),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_527),
.A2(n_514),
.B(n_505),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_554),
.A2(n_538),
.B(n_516),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_484),
.Y(n_556)
);

MAJx2_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_557),
.C(n_526),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_519),
.B(n_489),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_532),
.B(n_489),
.C(n_504),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_558),
.B(n_560),
.Y(n_570)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_521),
.Y(n_559)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_559),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_504),
.C(n_528),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_561),
.B(n_564),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_558),
.Y(n_563)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_563),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_544),
.A2(n_554),
.B(n_552),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_550),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_531),
.C(n_520),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_566),
.B(n_548),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_542),
.B(n_534),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_567),
.B(n_569),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_559),
.A2(n_521),
.B(n_537),
.C(n_540),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_530),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_574),
.Y(n_582)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_551),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_572),
.B(n_547),
.Y(n_579)
);

OAI322xp33_ASAP7_75t_L g573 ( 
.A1(n_553),
.A2(n_516),
.A3(n_538),
.B1(n_518),
.B2(n_525),
.C1(n_522),
.C2(n_517),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_576),
.C(n_560),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_529),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_577),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_551),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_543),
.A2(n_552),
.B1(n_547),
.B2(n_545),
.Y(n_577)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_579),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_561),
.A2(n_542),
.B(n_543),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_580),
.A2(n_583),
.B(n_591),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_581),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_584),
.B(n_587),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_570),
.B(n_556),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_585),
.B(n_590),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_571),
.B(n_557),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_564),
.A2(n_549),
.B1(n_555),
.B2(n_568),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_567),
.B(n_555),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_588),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_600),
.Y(n_603)
);

NAND4xp25_ASAP7_75t_SL g597 ( 
.A(n_589),
.B(n_574),
.C(n_569),
.D(n_563),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_601),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_582),
.B(n_566),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_598),
.B(n_590),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_578),
.B(n_562),
.C(n_577),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_582),
.B(n_575),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_578),
.C(n_586),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_602),
.B(n_595),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_599),
.A2(n_589),
.B(n_586),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_605),
.A2(n_606),
.B(n_596),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_593),
.A2(n_568),
.B(n_572),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_607),
.Y(n_612)
);

AOI31xp67_ASAP7_75t_L g608 ( 
.A1(n_594),
.A2(n_549),
.A3(n_587),
.B(n_565),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_608),
.B(n_600),
.C(n_597),
.Y(n_610)
);

AOI21xp33_ASAP7_75t_L g614 ( 
.A1(n_609),
.A2(n_604),
.B(n_603),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_610),
.B(n_611),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_614),
.A2(n_612),
.B1(n_602),
.B2(n_607),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_613),
.B(n_592),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_584),
.Y(n_617)
);


endmodule