module fake_jpeg_6315_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_46),
.Y(n_51)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_20),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_16),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_20),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_56),
.B(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_15),
.B1(n_29),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_21),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_33),
.A2(n_22),
.B1(n_18),
.B2(n_17),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_83),
.B1(n_3),
.B2(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_28),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_18),
.B1(n_28),
.B2(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_80),
.Y(n_108)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_25),
.B1(n_21),
.B2(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_21),
.B1(n_25),
.B2(n_5),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_2),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_3),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_104),
.B1(n_81),
.B2(n_52),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_113),
.Y(n_130)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_105),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_13),
.C(n_7),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_8),
.C(n_9),
.Y(n_139)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_11),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_61),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_82),
.B1(n_75),
.B2(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_67),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_121),
.Y(n_156)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_83),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_138),
.B(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_90),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_59),
.B1(n_63),
.B2(n_55),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_138),
.B1(n_106),
.B2(n_111),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_54),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_54),
.C(n_79),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_132),
.C(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_131),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_136),
.Y(n_147)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_102),
.B1(n_121),
.B2(n_119),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_59),
.B1(n_68),
.B2(n_51),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_68),
.B1(n_67),
.B2(n_79),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_92),
.B(n_11),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_153),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_151),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_159),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_115),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_161),
.B1(n_165),
.B2(n_131),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_158),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_107),
.Y(n_159)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_72),
.B1(n_60),
.B2(n_53),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_118),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_97),
.B(n_95),
.Y(n_164)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_72),
.B1(n_53),
.B2(n_110),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_139),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_141),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_184),
.B(n_150),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_126),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_120),
.C(n_90),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_124),
.C(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_189),
.B(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_162),
.B1(n_157),
.B2(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_200),
.B1(n_176),
.B2(n_155),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_150),
.B(n_167),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_199),
.B1(n_146),
.B2(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

OAI22x1_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_161),
.B1(n_151),
.B2(n_166),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_169),
.B1(n_175),
.B2(n_161),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_192),
.B1(n_200),
.B2(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_173),
.C(n_183),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_203),
.C(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_173),
.C(n_172),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_186),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_159),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_218),
.C(n_209),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_216),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_160),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_191),
.C(n_164),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_224),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_211),
.B(n_218),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_144),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_187),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_224),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_208),
.B(n_214),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

OAI31xp33_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_234),
.A3(n_230),
.B(n_193),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_235),
.Y(n_236)
);


endmodule