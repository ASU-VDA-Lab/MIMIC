module fake_jpeg_27249_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_28),
.B1(n_34),
.B2(n_36),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_48),
.B1(n_46),
.B2(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_24),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_79),
.B1(n_89),
.B2(n_24),
.Y(n_118)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_77),
.B(n_39),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_48),
.B1(n_34),
.B2(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_27),
.A3(n_29),
.B1(n_20),
.B2(n_32),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_19),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_94),
.Y(n_103)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_34),
.B1(n_36),
.B2(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_27),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_26),
.Y(n_109)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_104),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_39),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_102),
.A2(n_105),
.B1(n_117),
.B2(n_125),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_39),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_69),
.B1(n_56),
.B2(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_86),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_64),
.B1(n_69),
.B2(n_43),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_43),
.B1(n_41),
.B2(n_24),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_25),
.B1(n_41),
.B2(n_21),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_92),
.B1(n_93),
.B2(n_75),
.Y(n_137)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_103),
.B1(n_121),
.B2(n_109),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_81),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_146),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g147 ( 
.A(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_153),
.B1(n_155),
.B2(n_76),
.Y(n_179)
);

BUFx24_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_39),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_110),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_72),
.B1(n_91),
.B2(n_74),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_123),
.B(n_122),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_159),
.B(n_171),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_119),
.B(n_103),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_118),
.B1(n_117),
.B2(n_104),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_179),
.B1(n_183),
.B2(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_31),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_121),
.C(n_111),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_181),
.C(n_147),
.Y(n_191)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_111),
.B(n_119),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_170),
.B1(n_176),
.B2(n_154),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_156),
.B1(n_131),
.B2(n_132),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_144),
.B(n_145),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_128),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_178),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_136),
.B1(n_135),
.B2(n_142),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_23),
.C(n_93),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_155),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_110),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_147),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_129),
.A2(n_127),
.B1(n_108),
.B2(n_70),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_127),
.B(n_19),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_21),
.B(n_26),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_162),
.Y(n_241)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_193),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_171),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_209),
.B1(n_218),
.B2(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_194),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_150),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_199),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_19),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_216),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_161),
.B1(n_175),
.B2(n_172),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_150),
.C(n_149),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_178),
.C(n_181),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_130),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_26),
.B(n_8),
.Y(n_206)
);

AOI32xp33_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_15),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_138),
.Y(n_207)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_13),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_175),
.A2(n_33),
.B(n_17),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_209),
.B(n_205),
.Y(n_244)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_167),
.B(n_138),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_210),
.B(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_214),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_226),
.C(n_231),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_230),
.B1(n_237),
.B2(n_211),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_166),
.C(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_203),
.B1(n_196),
.B2(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_210),
.C(n_189),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_157),
.C(n_182),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_240),
.C(n_31),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_160),
.B1(n_172),
.B2(n_176),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_171),
.B1(n_162),
.B2(n_17),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_190),
.B1(n_208),
.B2(n_204),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_255),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_245),
.B1(n_223),
.B2(n_225),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_220),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_149),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_195),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_231),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_149),
.B1(n_31),
.B2(n_33),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_25),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_244),
.B(n_9),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_12),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_280),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_240),
.C(n_226),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_265),
.C(n_263),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_222),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_232),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_237),
.B1(n_258),
.B2(n_230),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_223),
.B(n_238),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_256),
.B(n_235),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_296),
.C(n_280),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_246),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_290),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_250),
.B1(n_252),
.B2(n_248),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_288),
.B1(n_268),
.B2(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_260),
.C(n_255),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_251),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_241),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_257),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_272),
.B1(n_274),
.B2(n_10),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_23),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_6),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_302),
.B(n_304),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_309),
.B1(n_291),
.B2(n_286),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_277),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_272),
.C(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_23),
.C(n_8),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_301),
.B1(n_12),
.B2(n_11),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_300),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_304),
.B1(n_302),
.B2(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_324),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_0),
.B(n_1),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_310),
.B(n_1),
.Y(n_325)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_0),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_327),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_330),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_322),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_316),
.C(n_321),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_333),
.B(n_334),
.C(n_335),
.D(n_329),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_319),
.B(n_2),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_5),
.B(n_2),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_1),
.C(n_3),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_5),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_3),
.C(n_4),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_5),
.B(n_3),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_3),
.B(n_4),
.Y(n_342)
);


endmodule