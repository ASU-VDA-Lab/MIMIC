module fake_ariane_508_n_730 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_730);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_730;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_672;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_40),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_74),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_87),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_12),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_80),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_44),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_8),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_25),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_41),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_18),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_47),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_42),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_118),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_46),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_26),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_79),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_52),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_12),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_56),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_6),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_136),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_13),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_49),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_71),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_141),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_59),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_94),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_58),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_33),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_137),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_2),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_0),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_3),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_4),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_4),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_5),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

OAI21x1_ASAP7_75t_L g230 ( 
.A1(n_162),
.A2(n_86),
.B(n_146),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_5),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_191),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_165),
.B(n_7),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_156),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_167),
.B(n_9),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_151),
.B(n_9),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_155),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_171),
.A2(n_91),
.B(n_145),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_151),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_177),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_225),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_161),
.B1(n_179),
.B2(n_177),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_172),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_178),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_179),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_149),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g272 ( 
.A(n_214),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_180),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_241),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_212),
.B(n_185),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

AND3x2_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_200),
.C(n_196),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_153),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_241),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

BUFx6f_ASAP7_75t_SL g291 ( 
.A(n_225),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_204),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_228),
.B(n_157),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_242),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_213),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_231),
.B(n_176),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_249),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_221),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_271),
.B(n_221),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

AND2x6_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_215),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_251),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_240),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_240),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_216),
.B1(n_210),
.B2(n_238),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_260),
.A2(n_253),
.B1(n_210),
.B2(n_247),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_251),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_288),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_227),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_L g325 ( 
.A(n_273),
.B(n_160),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_227),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_244),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_246),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_264),
.B(n_229),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_243),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_250),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_264),
.B(n_250),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_259),
.A2(n_254),
.B(n_230),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_255),
.B(n_247),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_248),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_235),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g340 ( 
.A1(n_292),
.A2(n_253),
.B(n_245),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_262),
.A2(n_277),
.B1(n_259),
.B2(n_272),
.Y(n_344)
);

BUFx6f_ASAP7_75t_SL g345 ( 
.A(n_272),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_280),
.B(n_163),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_282),
.B(n_239),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_L g349 ( 
.A(n_273),
.B(n_173),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_276),
.B(n_10),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_273),
.A2(n_195),
.B1(n_182),
.B2(n_206),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_288),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_291),
.B(n_183),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_267),
.B(n_224),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_267),
.B(n_234),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_257),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_270),
.B(n_186),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_SL g361 ( 
.A(n_258),
.B(n_194),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_263),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_270),
.B(n_263),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_265),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_311),
.A2(n_312),
.B1(n_305),
.B2(n_317),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_197),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_199),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_306),
.A2(n_275),
.B(n_301),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_335),
.A2(n_275),
.B(n_301),
.Y(n_370)
);

BUFx12f_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_310),
.A2(n_274),
.B(n_295),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_265),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_269),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_318),
.A2(n_304),
.B(n_295),
.C(n_287),
.Y(n_375)
);

BUFx4f_ASAP7_75t_L g376 ( 
.A(n_322),
.Y(n_376)
);

AO21x1_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_304),
.B(n_286),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_202),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_313),
.A2(n_283),
.B1(n_274),
.B2(n_269),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_283),
.B(n_15),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_316),
.B(n_11),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_352),
.A2(n_15),
.B1(n_16),
.B2(n_258),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_320),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_16),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_338),
.A2(n_234),
.B1(n_20),
.B2(n_21),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_319),
.A2(n_234),
.B(n_22),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_324),
.A2(n_19),
.B(n_23),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_24),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_391)
);

AOI22x1_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_326),
.A2(n_34),
.B(n_35),
.Y(n_393)
);

BUFx12f_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_363),
.A2(n_37),
.B(n_38),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_323),
.B(n_39),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_323),
.B(n_322),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_43),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_L g399 ( 
.A(n_323),
.B(n_45),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_336),
.A2(n_48),
.B(n_50),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_51),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_323),
.B(n_53),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_325),
.A2(n_54),
.B(n_57),
.Y(n_405)
);

AOI21xp33_ASAP7_75t_L g406 ( 
.A1(n_359),
.A2(n_349),
.B(n_314),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_61),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_353),
.A2(n_62),
.B(n_63),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_346),
.A2(n_64),
.B(n_65),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_323),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_360),
.A2(n_72),
.B(n_73),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_357),
.A2(n_75),
.B(n_76),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_358),
.A2(n_77),
.B(n_78),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_343),
.B(n_148),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_362),
.A2(n_81),
.B(n_84),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_355),
.A2(n_85),
.B(n_88),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_364),
.A2(n_93),
.B(n_95),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_347),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_315),
.A2(n_102),
.B(n_103),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_309),
.B(n_356),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_315),
.B(n_356),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_315),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_345),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_345),
.B(n_110),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_361),
.A2(n_112),
.B(n_114),
.Y(n_427)
);

BUFx12f_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_385),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_368),
.Y(n_430)
);

INVx3_ASAP7_75t_SL g431 ( 
.A(n_384),
.Y(n_431)
);

O2A1O1Ixp5_ASAP7_75t_L g432 ( 
.A1(n_367),
.A2(n_366),
.B(n_377),
.C(n_400),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_120),
.C(n_121),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_376),
.B(n_122),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_123),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_372),
.A2(n_125),
.B(n_127),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_381),
.A2(n_128),
.B(n_130),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_131),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_398),
.A2(n_134),
.B(n_135),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_379),
.A2(n_139),
.B(n_140),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_376),
.B(n_422),
.Y(n_444)
);

AO21x2_ASAP7_75t_L g445 ( 
.A1(n_411),
.A2(n_142),
.B(n_143),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_394),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_419),
.A2(n_416),
.B(n_413),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_375),
.A2(n_405),
.B(n_397),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_369),
.A2(n_407),
.B(n_415),
.Y(n_449)
);

NAND2x1p5_ASAP7_75t_L g450 ( 
.A(n_388),
.B(n_426),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_416),
.A2(n_408),
.B(n_393),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_414),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_404),
.Y(n_454)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_419),
.A2(n_412),
.B(n_399),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_406),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_423),
.A2(n_424),
.B(n_403),
.Y(n_457)
);

OA22x2_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_383),
.B1(n_420),
.B2(n_410),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_389),
.A2(n_396),
.B(n_395),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_392),
.A2(n_409),
.B(n_427),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_387),
.A2(n_380),
.B(n_418),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_386),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_421),
.A2(n_335),
.B(n_365),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_366),
.B(n_365),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_365),
.B(n_312),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_365),
.A2(n_317),
.B1(n_318),
.B2(n_385),
.Y(n_470)
);

AO31x2_ASAP7_75t_L g471 ( 
.A1(n_377),
.A2(n_335),
.A3(n_391),
.B(n_370),
.Y(n_471)
);

BUFx12f_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_370),
.A2(n_307),
.B(n_367),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_368),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_366),
.B(n_365),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_368),
.B(n_342),
.Y(n_477)
);

OAI33xp33_ASAP7_75t_L g478 ( 
.A1(n_365),
.A2(n_318),
.A3(n_261),
.B1(n_344),
.B2(n_311),
.B3(n_378),
.Y(n_478)
);

AO21x2_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_451),
.B(n_463),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_449),
.B(n_448),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_435),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_460),
.A2(n_451),
.B(n_459),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_432),
.A2(n_474),
.B(n_438),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_444),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_441),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_478),
.A2(n_469),
.B1(n_458),
.B2(n_440),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_475),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_461),
.A2(n_437),
.B(n_457),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_436),
.A2(n_429),
.B1(n_447),
.B2(n_469),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_456),
.A2(n_468),
.B1(n_467),
.B2(n_462),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_454),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_430),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_L g495 ( 
.A1(n_462),
.A2(n_433),
.B1(n_452),
.B2(n_439),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_462),
.A2(n_450),
.B1(n_433),
.B2(n_473),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_443),
.A2(n_434),
.B(n_442),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_466),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g499 ( 
.A1(n_471),
.A2(n_445),
.B(n_429),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_471),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_471),
.A2(n_428),
.B(n_472),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_431),
.B(n_446),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_464),
.A2(n_476),
.B(n_432),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_463),
.A2(n_449),
.B(n_448),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_463),
.A2(n_451),
.B(n_432),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_465),
.Y(n_508)
);

AO21x2_ASAP7_75t_L g509 ( 
.A1(n_455),
.A2(n_451),
.B(n_463),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_458),
.A2(n_214),
.B1(n_318),
.B2(n_272),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_470),
.B(n_444),
.Y(n_511)
);

NOR2x1_ASAP7_75t_R g512 ( 
.A(n_428),
.B(n_276),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_435),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_318),
.B1(n_478),
.B2(n_261),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_475),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

NOR2x1_ASAP7_75t_SL g518 ( 
.A(n_473),
.B(n_469),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_463),
.A2(n_449),
.B(n_448),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_435),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_500),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_511),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_498),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_485),
.A2(n_511),
.B1(n_481),
.B2(n_510),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_514),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_498),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_503),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_515),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_486),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_515),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_502),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_518),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_479),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_482),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_514),
.B(n_488),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_480),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_508),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_509),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_516),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_507),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_488),
.B(n_494),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_507),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_520),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_513),
.B(n_517),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_492),
.B(n_493),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_507),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_492),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_522),
.B(n_499),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_521),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_540),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_501),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_526),
.B(n_501),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_531),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_519),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_526),
.B(n_484),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_531),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_512),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_528),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_528),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_532),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_536),
.B(n_506),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_529),
.B(n_484),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_496),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_540),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_529),
.B(n_484),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_542),
.B(n_506),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_524),
.B(n_497),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_552),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_544),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_542),
.B(n_483),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_524),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_490),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_532),
.B(n_495),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_546),
.B(n_490),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_553),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_537),
.B(n_547),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_537),
.B(n_495),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_562),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_558),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_577),
.B(n_551),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_560),
.B(n_546),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_576),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_579),
.B(n_548),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_579),
.B(n_554),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_548),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_575),
.B(n_548),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_565),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_560),
.B(n_546),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_548),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_576),
.B(n_546),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_578),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_576),
.B(n_546),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_559),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_564),
.B(n_554),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_570),
.B(n_550),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_556),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_556),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_557),
.B(n_546),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_567),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_568),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_578),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_589),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_547),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_559),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_561),
.B(n_543),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_573),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_586),
.B(n_534),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_591),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_617),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_619),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_587),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_571),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_592),
.B(n_587),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_603),
.B(n_614),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_612),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_613),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_608),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_603),
.B(n_582),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_582),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_609),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_610),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_572),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_605),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_596),
.B(n_561),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_605),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_571),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_597),
.B(n_598),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_606),
.B(n_585),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_596),
.B(n_563),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_590),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_597),
.B(n_574),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_599),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_598),
.B(n_574),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_618),
.B(n_588),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_635),
.B(n_534),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_628),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_641),
.B(n_606),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_629),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_630),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_627),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_636),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_618),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_642),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_638),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_637),
.B(n_607),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_625),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_643),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_640),
.B(n_594),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_645),
.Y(n_662)
);

XOR2x2_ASAP7_75t_L g663 ( 
.A(n_635),
.B(n_566),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_622),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_621),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_642),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_647),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_623),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_654),
.Y(n_669)
);

AOI222xp33_ASAP7_75t_L g670 ( 
.A1(n_656),
.A2(n_626),
.B1(n_624),
.B2(n_611),
.C1(n_604),
.C2(n_602),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_661),
.B(n_625),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_652),
.Y(n_672)
);

OAI222xp33_ASAP7_75t_L g673 ( 
.A1(n_656),
.A2(n_525),
.B1(n_604),
.B2(n_602),
.C1(n_632),
.C2(n_611),
.Y(n_673)
);

OAI21xp33_ASAP7_75t_L g674 ( 
.A1(n_666),
.A2(n_631),
.B(n_647),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_646),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_658),
.B(n_639),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_657),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_664),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_665),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_675),
.A2(n_659),
.B1(n_648),
.B2(n_650),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_672),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_674),
.B(n_650),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_669),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_676),
.B(n_653),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_678),
.B(n_652),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_677),
.B(n_668),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_683),
.Y(n_687)
);

AOI211xp5_ASAP7_75t_SL g688 ( 
.A1(n_680),
.A2(n_673),
.B(n_675),
.C(n_649),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_681),
.B(n_661),
.Y(n_689)
);

OAI221xp5_ASAP7_75t_L g690 ( 
.A1(n_682),
.A2(n_670),
.B1(n_663),
.B2(n_651),
.C(n_662),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_685),
.B(n_673),
.C(n_660),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_684),
.A2(n_604),
.B(n_602),
.C(n_593),
.Y(n_692)
);

OAI211xp5_ASAP7_75t_SL g693 ( 
.A1(n_688),
.A2(n_686),
.B(n_667),
.C(n_633),
.Y(n_693)
);

NAND4xp75_ASAP7_75t_L g694 ( 
.A(n_689),
.B(n_583),
.C(n_634),
.D(n_527),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_687),
.B(n_671),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_690),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_693),
.B(n_691),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_696),
.A2(n_692),
.B1(n_600),
.B2(n_593),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_697),
.B(n_694),
.C(n_695),
.Y(n_699)
);

NOR2x1_ASAP7_75t_L g700 ( 
.A(n_698),
.B(n_533),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_697),
.B(n_655),
.Y(n_701)
);

NOR2x1_ASAP7_75t_L g702 ( 
.A(n_701),
.B(n_533),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_699),
.B(n_679),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_700),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_701),
.Y(n_705)
);

XNOR2xp5_ASAP7_75t_L g706 ( 
.A(n_701),
.B(n_535),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_703),
.A2(n_539),
.B(n_541),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_705),
.A2(n_527),
.B(n_541),
.C(n_535),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_704),
.B(n_615),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_615),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_702),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_646),
.Y(n_712)
);

XOR2x2_ASAP7_75t_L g713 ( 
.A(n_712),
.B(n_593),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_710),
.A2(n_539),
.B1(n_583),
.B2(n_600),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_709),
.A2(n_539),
.B(n_541),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_711),
.A2(n_533),
.B1(n_615),
.B2(n_530),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_707),
.A2(n_607),
.B1(n_615),
.B2(n_608),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_713),
.Y(n_718)
);

OA21x2_ASAP7_75t_L g719 ( 
.A1(n_715),
.A2(n_708),
.B(n_539),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_717),
.A2(n_716),
.B1(n_714),
.B2(n_615),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_716),
.Y(n_721)
);

AO21x1_ASAP7_75t_L g722 ( 
.A1(n_721),
.A2(n_639),
.B(n_644),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_718),
.A2(n_530),
.B(n_538),
.C(n_594),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_720),
.B(n_644),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_SL g725 ( 
.A1(n_719),
.A2(n_580),
.B(n_600),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_724),
.Y(n_726)
);

AOI21xp33_ASAP7_75t_SL g727 ( 
.A1(n_723),
.A2(n_722),
.B(n_725),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_726),
.A2(n_727),
.B(n_530),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_728),
.B(n_601),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_729),
.A2(n_538),
.B(n_581),
.Y(n_730)
);


endmodule