module fake_aes_1581_n_25 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
AOI21x1_ASAP7_75t_L g13 ( .A1(n_1), .A2(n_5), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_16), .B(n_0), .Y(n_17) );
INVx1_ASAP7_75t_SL g18 ( .A(n_15), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_14), .B1(n_18), .B2(n_13), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AOI222xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_14), .B1(n_19), .B2(n_3), .C1(n_4), .C2(n_2), .Y(n_22) );
NAND2xp5_ASAP7_75t_SL g23 ( .A(n_22), .B(n_19), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_13), .B1(n_2), .B2(n_3), .Y(n_24) );
AOI322xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_0), .A3(n_4), .B1(n_6), .B2(n_7), .C1(n_11), .C2(n_12), .Y(n_25) );
endmodule