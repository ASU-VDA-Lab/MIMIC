module fake_jpeg_3046_n_502 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_76),
.Y(n_110)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_29),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_74),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_18),
.B(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_33),
.Y(n_82)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_19),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_97),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_96),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_2),
.Y(n_97)
);

NAND2x1_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_77),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_28),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_96),
.B1(n_93),
.B2(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_103),
.A2(n_132),
.B1(n_60),
.B2(n_94),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_23),
.C(n_25),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_40),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_106),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_29),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_112),
.B(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_32),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_55),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_21),
.B1(n_41),
.B2(n_43),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g197 ( 
.A1(n_125),
.A2(n_147),
.B1(n_45),
.B2(n_43),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_32),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_156),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_82),
.A2(n_27),
.B1(n_40),
.B2(n_19),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_58),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_142),
.B1(n_66),
.B2(n_65),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_39),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_59),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g147 ( 
.A1(n_92),
.A2(n_46),
.B1(n_38),
.B2(n_34),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_83),
.B(n_39),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_55),
.B(n_40),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_86),
.B(n_46),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_38),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_68),
.B(n_40),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_161),
.B(n_197),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_162),
.Y(n_249)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_117),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_167),
.B(n_185),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_168),
.A2(n_170),
.B1(n_176),
.B2(n_181),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_169),
.B(n_180),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_102),
.A2(n_38),
.B1(n_46),
.B2(n_40),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_172),
.A2(n_175),
.B1(n_191),
.B2(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_80),
.B1(n_71),
.B2(n_70),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_179),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_63),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_118),
.A2(n_62),
.B1(n_64),
.B2(n_21),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

CKINVDCx6p67_ASAP7_75t_R g184 ( 
.A(n_111),
.Y(n_184)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_189),
.B(n_192),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_45),
.B1(n_37),
.B2(n_42),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_190),
.A2(n_206),
.B1(n_141),
.B2(n_136),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_108),
.A2(n_41),
.B1(n_42),
.B2(n_37),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_110),
.B(n_68),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_122),
.B(n_94),
.CI(n_73),
.CON(n_193),
.SN(n_193)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_137),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_129),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_201),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_132),
.A2(n_41),
.B(n_57),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_103),
.A2(n_37),
.B1(n_78),
.B2(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_123),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_98),
.B(n_3),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_217),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_31),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_133),
.A2(n_154),
.B1(n_116),
.B2(n_155),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_216),
.B1(n_127),
.B2(n_135),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_113),
.B(n_3),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_212),
.Y(n_258)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_130),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_155),
.A2(n_31),
.B1(n_5),
.B2(n_6),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_127),
.B1(n_141),
.B2(n_136),
.Y(n_228)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_116),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_174),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_227),
.C(n_244),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_228),
.A2(n_243),
.B1(n_252),
.B2(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_109),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_232),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_124),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_SL g315 ( 
.A1(n_234),
.A2(n_240),
.B(n_7),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_169),
.B(n_135),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_251),
.C(n_180),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_266),
.B1(n_180),
.B2(n_199),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_182),
.C(n_194),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_163),
.A2(n_146),
.B1(n_119),
.B2(n_137),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_169),
.B(n_119),
.C(n_146),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_171),
.A2(n_144),
.B1(n_143),
.B2(n_140),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_160),
.B(n_152),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_193),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_188),
.Y(n_256)
);

INVx4_ASAP7_75t_SL g308 ( 
.A(n_256),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_173),
.A2(n_144),
.B1(n_143),
.B2(n_140),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_165),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_260),
.B(n_225),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_178),
.B(n_152),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_185),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_210),
.A2(n_152),
.B1(n_144),
.B2(n_143),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_271),
.B(n_258),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_226),
.A2(n_161),
.B1(n_193),
.B2(n_206),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_282),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_195),
.B(n_167),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_276),
.A2(n_300),
.B(n_312),
.Y(n_342)
);

OA22x2_ASAP7_75t_L g321 ( 
.A1(n_277),
.A2(n_243),
.B1(n_252),
.B2(n_257),
.Y(n_321)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_223),
.Y(n_281)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_226),
.A2(n_175),
.B1(n_197),
.B2(n_164),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_299),
.B1(n_264),
.B2(n_253),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_298),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_285),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_221),
.B(n_202),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_288),
.Y(n_341)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_164),
.B(n_204),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_306),
.C(n_314),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_231),
.A2(n_235),
.B1(n_220),
.B2(n_221),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_177),
.C(n_196),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_296),
.C(n_303),
.Y(n_340)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_232),
.B(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_293),
.B(n_258),
.Y(n_352)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_231),
.B(n_197),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_302),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_183),
.C(n_179),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_198),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_235),
.A2(n_212),
.B1(n_201),
.B2(n_159),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_249),
.A2(n_213),
.B(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_242),
.A2(n_215),
.B1(n_200),
.B2(n_208),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_236),
.B(n_205),
.C(n_217),
.Y(n_303)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_233),
.A2(n_205),
.B1(n_187),
.B2(n_166),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_310),
.B(n_258),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_186),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_241),
.A2(n_140),
.B1(n_126),
.B2(n_186),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_309),
.A2(n_317),
.B1(n_244),
.B2(n_227),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g310 ( 
.A1(n_233),
.A2(n_126),
.B1(n_186),
.B2(n_7),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_242),
.A2(n_5),
.B(n_6),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

BUFx4f_ASAP7_75t_SL g353 ( 
.A(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_242),
.B(n_126),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_262),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_236),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_321),
.A2(n_310),
.B(n_305),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_251),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_354),
.C(n_308),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_283),
.A2(n_237),
.B1(n_249),
.B2(n_248),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_333),
.B1(n_337),
.B2(n_343),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_332),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_335),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_307),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_295),
.A2(n_276),
.B1(n_282),
.B2(n_277),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_256),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_339),
.B(n_357),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_275),
.A2(n_218),
.B1(n_266),
.B2(n_222),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_275),
.A2(n_304),
.B1(n_306),
.B2(n_314),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_352),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_300),
.A2(n_238),
.B(n_224),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_346),
.A2(n_348),
.B(n_310),
.Y(n_377)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_304),
.B(n_262),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_347),
.Y(n_360)
);

XNOR2x2_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_245),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_291),
.Y(n_358)
);

XNOR2x2_ASAP7_75t_SL g356 ( 
.A(n_312),
.B(n_271),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_268),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_219),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_386),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_347),
.Y(n_361)
);

INVx11_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_330),
.A2(n_337),
.B1(n_320),
.B2(n_333),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_372),
.B1(n_348),
.B2(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_382),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_303),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_373),
.C(n_379),
.Y(n_412)
);

OA22x2_ASAP7_75t_L g367 ( 
.A1(n_348),
.A2(n_310),
.B1(n_305),
.B2(n_272),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

OAI32xp33_ASAP7_75t_L g371 ( 
.A1(n_326),
.A2(n_313),
.A3(n_294),
.B1(n_297),
.B2(n_302),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_347),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_376),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_317),
.B(n_274),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_319),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_378),
.B(n_383),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_342),
.A2(n_240),
.B(n_305),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_325),
.A2(n_230),
.B(n_218),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_355),
.A2(n_281),
.B1(n_223),
.B2(n_259),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_385),
.A2(n_387),
.B1(n_391),
.B2(n_324),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_355),
.A2(n_259),
.B1(n_292),
.B2(n_269),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_346),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_345),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_268),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_390),
.C(n_373),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_250),
.C(n_269),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_341),
.A2(n_250),
.B1(n_230),
.B2(n_11),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_393),
.Y(n_421)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_369),
.A2(n_341),
.B1(n_334),
.B2(n_326),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_396),
.A2(n_403),
.B1(n_388),
.B2(n_361),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_398),
.A2(n_360),
.B1(n_366),
.B2(n_377),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_356),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_409),
.Y(n_429)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_369),
.A2(n_325),
.B1(n_356),
.B2(n_321),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_405),
.A2(n_408),
.B1(n_413),
.B2(n_417),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_372),
.A2(n_343),
.B1(n_349),
.B2(n_353),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_365),
.B(n_344),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_372),
.A2(n_353),
.B1(n_344),
.B2(n_336),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_331),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_416),
.C(n_324),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_374),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_359),
.B(n_331),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_362),
.A2(n_353),
.B1(n_336),
.B2(n_327),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_427),
.B1(n_442),
.B2(n_413),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_389),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_426),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_395),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_431),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_419),
.A2(n_375),
.B(n_368),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_440),
.B(n_405),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_386),
.C(n_358),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_439),
.C(n_441),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_390),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_433),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_374),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_383),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_371),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_396),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_410),
.A2(n_376),
.B1(n_366),
.B2(n_382),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_435),
.A2(n_437),
.B1(n_432),
.B2(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_410),
.A2(n_368),
.B1(n_367),
.B2(n_381),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_391),
.Y(n_438)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_385),
.C(n_380),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_406),
.A2(n_367),
.B(n_370),
.C(n_321),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_387),
.C(n_327),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_327),
.B1(n_321),
.B2(n_335),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_443),
.A2(n_451),
.B1(n_418),
.B2(n_407),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_454),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_408),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_460),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_429),
.B(n_401),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

AOI211xp5_ASAP7_75t_L g448 ( 
.A1(n_437),
.A2(n_406),
.B(n_399),
.C(n_393),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_448),
.B(n_394),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_441),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_425),
.Y(n_473)
);

INVx11_ASAP7_75t_L g451 ( 
.A(n_440),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_399),
.C(n_392),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_439),
.C(n_433),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_430),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_458),
.B1(n_461),
.B2(n_427),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_435),
.A2(n_442),
.B1(n_421),
.B2(n_420),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_351),
.Y(n_460)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_461),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_466),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_351),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_467),
.A2(n_444),
.B1(n_457),
.B2(n_459),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_456),
.A2(n_429),
.B(n_426),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_468),
.A2(n_469),
.B(n_464),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_458),
.A2(n_418),
.B(n_407),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_471),
.A2(n_472),
.B1(n_464),
.B2(n_475),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_474),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_328),
.Y(n_474)
);

AO22x1_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_394),
.B1(n_411),
.B2(n_328),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_453),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_476),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_450),
.C(n_455),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_9),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g486 ( 
.A1(n_478),
.A2(n_470),
.B1(n_468),
.B2(n_462),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_473),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_483),
.Y(n_492)
);

AOI31xp67_ASAP7_75t_L g487 ( 
.A1(n_481),
.A2(n_484),
.A3(n_470),
.B(n_446),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_450),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_482),
.A2(n_10),
.B(n_11),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_459),
.B(n_455),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_486),
.A2(n_490),
.B(n_14),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_487),
.A2(n_477),
.B1(n_13),
.B2(n_14),
.Y(n_494)
);

AOI322xp5_ASAP7_75t_L g488 ( 
.A1(n_476),
.A2(n_469),
.A3(n_462),
.B1(n_475),
.B2(n_463),
.C1(n_13),
.C2(n_14),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_485),
.C(n_479),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_489),
.B(n_12),
.Y(n_495)
);

AO21x1_ASAP7_75t_SL g498 ( 
.A1(n_493),
.A2(n_494),
.B(n_496),
.Y(n_498)
);

NOR3xp33_ASAP7_75t_SL g497 ( 
.A(n_495),
.B(n_488),
.C(n_491),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_492),
.C(n_15),
.Y(n_499)
);

AOI322xp5_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_15),
.A3(n_16),
.B1(n_498),
.B2(n_245),
.C1(n_474),
.C2(n_272),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_15),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_15),
.Y(n_502)
);


endmodule