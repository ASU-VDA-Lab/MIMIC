module fake_netlist_5_1014_n_966 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_966);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_966;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_443;
wire n_293;
wire n_372;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_856;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_964;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_928;
wire n_858;
wire n_829;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_781;
wire n_834;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_857;
wire n_795;
wire n_695;
wire n_832;
wire n_707;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_914;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_960;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g190 ( 
.A(n_79),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_109),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_67),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_96),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_27),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_9),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_89),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_39),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_73),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_131),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_62),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_144),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_56),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_187),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_40),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_69),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_64),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_151),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_95),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_45),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

INVxp33_ASAP7_75t_R g231 ( 
.A(n_59),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_99),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_20),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_5),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_42),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_139),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_49),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_43),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_178),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_19),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_75),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_93),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_84),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_68),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_105),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_26),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_148),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_54),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_98),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_17),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_32),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_111),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_133),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_0),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_191),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_222),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_195),
.B(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_195),
.B(n_0),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_243),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_193),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_226),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_194),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_197),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_1),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_201),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_203),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_204),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_230),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_249),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_206),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_216),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_207),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_241),
.B(n_217),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_249),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_217),
.B(n_1),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_255),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_190),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_237),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_208),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_192),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_199),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_205),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_210),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_255),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_264),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_211),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_212),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_209),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_302),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_239),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_200),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_237),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_258),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_278),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_214),
.Y(n_342)
);

BUFx8_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

AND3x2_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_215),
.C(n_213),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_287),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_318),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_285),
.B(n_225),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

BUFx8_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_268),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_294),
.B(n_300),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_289),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_292),
.B(n_218),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_227),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_271),
.B(n_264),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_271),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_272),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_272),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_322),
.A2(n_314),
.B1(n_304),
.B2(n_246),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_323),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_320),
.B(n_314),
.Y(n_377)
);

CKINVDCx8_ASAP7_75t_R g378 ( 
.A(n_367),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_240),
.Y(n_379)
);

BUFx6f_ASAP7_75t_SL g380 ( 
.A(n_355),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_219),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_245),
.B1(n_265),
.B2(n_263),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_328),
.B(n_244),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_220),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_319),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_248),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_L g393 ( 
.A1(n_365),
.A2(n_253),
.B1(n_259),
.B2(n_262),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_221),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_223),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_342),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_231),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_352),
.B(n_266),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_361),
.B(n_24),
.Y(n_405)
);

BUFx4f_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_224),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_328),
.B(n_228),
.Y(n_408)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_25),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_348),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_229),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_328),
.B(n_232),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_328),
.B(n_233),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_327),
.B(n_257),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_356),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_351),
.B(n_238),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_321),
.A2(n_252),
.B1(n_251),
.B2(n_247),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_330),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_331),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_339),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_339),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g434 ( 
.A(n_362),
.B(n_28),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_331),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_347),
.B(n_254),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_330),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_357),
.B(n_2),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_2),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_347),
.B(n_29),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_341),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_357),
.B(n_30),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_354),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_377),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_347),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_354),
.Y(n_451)
);

AO22x2_ASAP7_75t_L g452 ( 
.A1(n_375),
.A2(n_368),
.B1(n_366),
.B2(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

OAI221xp5_ASAP7_75t_L g454 ( 
.A1(n_382),
.A2(n_358),
.B1(n_353),
.B2(n_345),
.C(n_341),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_389),
.B(n_359),
.Y(n_455)
);

NAND2x1p5_ASAP7_75t_L g456 ( 
.A(n_385),
.B(n_354),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g459 ( 
.A1(n_375),
.A2(n_368),
.B1(n_366),
.B2(n_372),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_354),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_419),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_413),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_400),
.A2(n_363),
.B1(n_359),
.B2(n_364),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_437),
.A2(n_406),
.B1(n_399),
.B2(n_443),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_376),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g475 ( 
.A1(n_428),
.A2(n_370),
.B1(n_373),
.B2(n_374),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_380),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_381),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_324),
.Y(n_480)
);

AO22x2_ASAP7_75t_L g481 ( 
.A1(n_428),
.A2(n_370),
.B1(n_373),
.B2(n_374),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_413),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_425),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_425),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_367),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_446),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_440),
.A2(n_369),
.B1(n_371),
.B2(n_353),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_406),
.B(n_325),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_441),
.A2(n_332),
.B1(n_334),
.B2(n_340),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_420),
.A2(n_356),
.B1(n_343),
.B2(n_371),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_421),
.B(n_338),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_423),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_380),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_427),
.A2(n_369),
.B1(n_371),
.B2(n_334),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_431),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_423),
.B(n_332),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_407),
.B(n_371),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_407),
.B(n_341),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_387),
.Y(n_505)
);

AO22x2_ASAP7_75t_L g506 ( 
.A1(n_388),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_411),
.B(n_345),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_379),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_398),
.B(n_345),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_442),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_398),
.B(n_345),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_379),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_386),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_386),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_402),
.A2(n_340),
.B1(n_356),
.B2(n_343),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_344),
.Y(n_516)
);

OAI221xp5_ASAP7_75t_L g517 ( 
.A1(n_392),
.A2(n_340),
.B1(n_335),
.B2(n_337),
.C(n_329),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_392),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_387),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_430),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

AO22x2_ASAP7_75t_L g525 ( 
.A1(n_393),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_525)
);

NAND2x1p5_ASAP7_75t_L g526 ( 
.A(n_445),
.B(n_340),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_445),
.B(n_329),
.Y(n_528)
);

AO22x2_ASAP7_75t_L g529 ( 
.A1(n_397),
.A2(n_415),
.B1(n_416),
.B2(n_408),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_405),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_409),
.B(n_336),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_409),
.B(n_335),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_SL g534 ( 
.A(n_455),
.B(n_477),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_451),
.B(n_439),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_493),
.B(n_397),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_450),
.B(n_442),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_478),
.B(n_409),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_480),
.B(n_343),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_460),
.B(n_343),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_465),
.B(n_408),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_466),
.B(n_378),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_490),
.B(n_415),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_491),
.B(n_502),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_416),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_489),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_504),
.B(n_356),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_461),
.B(n_445),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_337),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_483),
.B(n_390),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_497),
.B(n_390),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_516),
.B(n_391),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_516),
.B(n_391),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_410),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_503),
.B(n_391),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_453),
.B(n_404),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_522),
.B(n_404),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_457),
.B(n_404),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_521),
.B(n_418),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_458),
.B(n_462),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_515),
.B(n_418),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_494),
.B(n_418),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_469),
.B(n_410),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_470),
.B(n_511),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_495),
.B(n_456),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_449),
.B(n_410),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_467),
.B(n_468),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_484),
.B(n_424),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_533),
.B(n_424),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_523),
.B(n_434),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_527),
.B(n_434),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_530),
.B(n_434),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_471),
.B(n_472),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_485),
.B(n_532),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_463),
.B(n_434),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_449),
.B(n_12),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_464),
.B(n_31),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_473),
.B(n_13),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_487),
.B(n_14),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_519),
.B(n_14),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_486),
.B(n_33),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_492),
.B(n_15),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_524),
.B(n_15),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_474),
.B(n_476),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_479),
.B(n_482),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_528),
.B(n_35),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_531),
.B(n_36),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_507),
.B(n_37),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_SL g589 ( 
.A(n_520),
.B(n_16),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_509),
.B(n_38),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_498),
.B(n_41),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_501),
.B(n_44),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_505),
.B(n_526),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_488),
.B(n_46),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_492),
.B(n_16),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_529),
.B(n_17),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_566),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_566),
.B(n_499),
.Y(n_598)
);

AO31x2_ASAP7_75t_L g599 ( 
.A1(n_596),
.A2(n_529),
.A3(n_475),
.B(n_481),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_546),
.B(n_488),
.Y(n_600)
);

AOI21xp33_ASAP7_75t_L g601 ( 
.A1(n_544),
.A2(n_452),
.B(n_459),
.Y(n_601)
);

OAI21x1_ASAP7_75t_L g602 ( 
.A1(n_563),
.A2(n_517),
.B(n_454),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_573),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_508),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_542),
.B(n_452),
.C(n_459),
.Y(n_605)
);

AOI31xp33_ASAP7_75t_L g606 ( 
.A1(n_547),
.A2(n_525),
.A3(n_506),
.B(n_481),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_560),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_545),
.A2(n_500),
.B(n_475),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_546),
.B(n_500),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_525),
.Y(n_610)
);

AO21x2_ASAP7_75t_L g611 ( 
.A1(n_564),
.A2(n_518),
.B(n_512),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_549),
.B(n_506),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_543),
.B(n_508),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_534),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_554),
.A2(n_117),
.B(n_188),
.Y(n_615)
);

AO31x2_ASAP7_75t_L g616 ( 
.A1(n_580),
.A2(n_518),
.A3(n_512),
.B(n_20),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_576),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_584),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_536),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_562),
.A2(n_116),
.B(n_184),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_567),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_594),
.B(n_47),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_565),
.A2(n_119),
.B1(n_183),
.B2(n_181),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_570),
.A2(n_114),
.B(n_180),
.Y(n_624)
);

BUFx2_ASAP7_75t_SL g625 ( 
.A(n_535),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_538),
.A2(n_112),
.B(n_176),
.Y(n_626)
);

AO31x2_ASAP7_75t_L g627 ( 
.A1(n_575),
.A2(n_595),
.A3(n_561),
.B(n_541),
.Y(n_627)
);

NAND2x1p5_ASAP7_75t_L g628 ( 
.A(n_552),
.B(n_48),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_537),
.B(n_18),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_574),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_553),
.B(n_21),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_571),
.A2(n_123),
.B(n_50),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_557),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_568),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_548),
.B(n_22),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_572),
.A2(n_124),
.B(n_51),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_550),
.B(n_22),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_578),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_539),
.B(n_52),
.Y(n_639)
);

OAI22x1_ASAP7_75t_L g640 ( 
.A1(n_540),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_555),
.Y(n_641)
);

AOI31xp67_ASAP7_75t_L g642 ( 
.A1(n_587),
.A2(n_58),
.A3(n_60),
.B(n_61),
.Y(n_642)
);

AOI21xp33_ASAP7_75t_L g643 ( 
.A1(n_551),
.A2(n_63),
.B(n_65),
.Y(n_643)
);

AOI221x1_ASAP7_75t_L g644 ( 
.A1(n_579),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.C(n_76),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_585),
.B(n_77),
.Y(n_645)
);

CKINVDCx14_ASAP7_75t_R g646 ( 
.A(n_583),
.Y(n_646)
);

OAI22x1_ASAP7_75t_L g647 ( 
.A1(n_556),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_558),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_569),
.A2(n_82),
.B(n_83),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_593),
.B(n_85),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_608),
.A2(n_590),
.B(n_588),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_622),
.A2(n_586),
.B1(n_577),
.B2(n_592),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_617),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_603),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g655 ( 
.A1(n_601),
.A2(n_589),
.B1(n_591),
.B2(n_581),
.C(n_559),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_186),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_607),
.Y(n_657)
);

AO21x2_ASAP7_75t_L g658 ( 
.A1(n_613),
.A2(n_86),
.B(n_87),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_618),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_615),
.A2(n_88),
.B(n_90),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_641),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_621),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_604),
.A2(n_94),
.B1(n_97),
.B2(n_100),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_614),
.Y(n_664)
);

AOI22x1_ASAP7_75t_L g665 ( 
.A1(n_640),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_630),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_624),
.A2(n_108),
.B(n_110),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_597),
.B(n_115),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_630),
.Y(n_669)
);

NAND2x1_ASAP7_75t_L g670 ( 
.A(n_648),
.B(n_126),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_604),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_605),
.B(n_173),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_602),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_627),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_648),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_620),
.A2(n_130),
.B(n_132),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_626),
.A2(n_136),
.B(n_137),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_597),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_619),
.B(n_138),
.C(n_141),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_600),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_638),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_681)
);

CKINVDCx16_ASAP7_75t_R g682 ( 
.A(n_600),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_612),
.B(n_146),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_610),
.B(n_147),
.Y(n_685)
);

OAI21x1_ASAP7_75t_SL g686 ( 
.A1(n_632),
.A2(n_150),
.B(n_152),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_637),
.A2(n_153),
.B(n_154),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_627),
.Y(n_688)
);

AOI21xp33_ASAP7_75t_L g689 ( 
.A1(n_629),
.A2(n_156),
.B(n_157),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_625),
.B(n_158),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_604),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_692)
);

OAI221xp5_ASAP7_75t_L g693 ( 
.A1(n_610),
.A2(n_163),
.B1(n_165),
.B2(n_167),
.C(n_168),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_627),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_599),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_634),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_636),
.A2(n_169),
.B(n_170),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_649),
.A2(n_172),
.B(n_623),
.Y(n_698)
);

CKINVDCx11_ASAP7_75t_R g699 ( 
.A(n_633),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_599),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_642),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_673),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_695),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_700),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_654),
.B(n_599),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_674),
.Y(n_707)
);

OA21x2_ASAP7_75t_L g708 ( 
.A1(n_674),
.A2(n_644),
.B(n_606),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_688),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_672),
.A2(n_604),
.B1(n_646),
.B2(n_639),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_688),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_684),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_694),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_694),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_673),
.Y(n_715)
);

BUFx12f_ASAP7_75t_L g716 ( 
.A(n_699),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_666),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_666),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_653),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_653),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_701),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_684),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_669),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_667),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_667),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_702),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_680),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_675),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_699),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_662),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_664),
.Y(n_731)
);

AO21x2_ASAP7_75t_L g732 ( 
.A1(n_651),
.A2(n_611),
.B(n_643),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_660),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_690),
.B(n_635),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_660),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_696),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_665),
.A2(n_650),
.B1(n_647),
.B2(n_598),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_661),
.A2(n_645),
.B1(n_650),
.B2(n_628),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_696),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_676),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_682),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_658),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_658),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_658),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_657),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_684),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_659),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_679),
.A2(n_616),
.B1(n_687),
.B2(n_656),
.Y(n_749)
);

AO21x2_ASAP7_75t_L g750 ( 
.A1(n_686),
.A2(n_616),
.B(n_698),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_670),
.Y(n_751)
);

AO21x2_ASAP7_75t_L g752 ( 
.A1(n_686),
.A2(n_616),
.B(n_698),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_676),
.A2(n_677),
.B(n_697),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_684),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_670),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_678),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_683),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_677),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_697),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_683),
.B(n_668),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_664),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_678),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_734),
.B(n_685),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_716),
.B(n_691),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_716),
.B(n_691),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_723),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_R g767 ( 
.A(n_729),
.B(n_691),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_742),
.B(n_668),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_757),
.B(n_691),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_760),
.B(n_668),
.Y(n_770)
);

BUFx10_ASAP7_75t_L g771 ( 
.A(n_754),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_761),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_R g773 ( 
.A(n_757),
.B(n_678),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_727),
.B(n_692),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_760),
.B(n_681),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_R g776 ( 
.A(n_708),
.B(n_706),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_720),
.Y(n_777)
);

OR2x4_ASAP7_75t_L g778 ( 
.A(n_723),
.B(n_693),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_719),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_R g780 ( 
.A(n_708),
.B(n_663),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_R g781 ( 
.A(n_731),
.B(n_671),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_R g782 ( 
.A(n_708),
.B(n_689),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_R g783 ( 
.A(n_708),
.B(n_652),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_726),
.B(n_655),
.Y(n_784)
);

XNOR2xp5_ASAP7_75t_L g785 ( 
.A(n_710),
.B(n_738),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_756),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_762),
.B(n_748),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_746),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_748),
.B(n_746),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_748),
.B(n_737),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_728),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_R g792 ( 
.A(n_747),
.B(n_722),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_735),
.B(n_737),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_R g794 ( 
.A(n_706),
.B(n_751),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_747),
.B(n_722),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_747),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_735),
.B(n_740),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_728),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_712),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_712),
.B(n_710),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_730),
.B(n_740),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_R g802 ( 
.A(n_730),
.B(n_755),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_739),
.B(n_718),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_R g804 ( 
.A(n_751),
.B(n_755),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_R g805 ( 
.A(n_741),
.B(n_736),
.Y(n_805)
);

XOR2x2_ASAP7_75t_SL g806 ( 
.A(n_749),
.B(n_745),
.Y(n_806)
);

XNOR2xp5_ASAP7_75t_L g807 ( 
.A(n_717),
.B(n_718),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_717),
.B(n_750),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_750),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_704),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_704),
.Y(n_811)
);

OAI221xp5_ASAP7_75t_SL g812 ( 
.A1(n_785),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.C(n_758),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_810),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_811),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_763),
.B(n_750),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_774),
.A2(n_752),
.B1(n_732),
.B2(n_759),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_773),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_766),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_808),
.B(n_705),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_787),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_802),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_791),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_798),
.B(n_705),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_789),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_788),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_801),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_771),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_752),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_790),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_809),
.B(n_744),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_797),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_793),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_803),
.B(n_743),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_803),
.B(n_800),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_786),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_807),
.B(n_743),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_806),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_784),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_783),
.B(n_782),
.C(n_767),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_775),
.A2(n_752),
.B1(n_732),
.B2(n_759),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_777),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_796),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_769),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_769),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_764),
.B(n_703),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_778),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_837),
.B(n_780),
.C(n_804),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_845),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_818),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_818),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_821),
.B(n_764),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_822),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_841),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_845),
.Y(n_854)
);

AOI221xp5_ASAP7_75t_L g855 ( 
.A1(n_837),
.A2(n_846),
.B1(n_815),
.B2(n_838),
.C(n_839),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_819),
.B(n_758),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_821),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_822),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_825),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_813),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_817),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_834),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_819),
.B(n_836),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_813),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_814),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_831),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_820),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_825),
.Y(n_868)
);

NAND4xp25_ASAP7_75t_L g869 ( 
.A(n_846),
.B(n_776),
.C(n_794),
.D(n_768),
.Y(n_869)
);

OAI31xp33_ASAP7_75t_L g870 ( 
.A1(n_812),
.A2(n_770),
.A3(n_772),
.B(n_781),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_836),
.B(n_765),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_863),
.B(n_843),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_865),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_849),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_828),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_861),
.B(n_863),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_867),
.B(n_844),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_862),
.B(n_844),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_850),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_857),
.B(n_827),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_859),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_852),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_865),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_858),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_855),
.B(n_840),
.C(n_816),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_862),
.B(n_844),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_860),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_848),
.B(n_854),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_864),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_880),
.B(n_853),
.Y(n_890)
);

AO221x2_ASAP7_75t_L g891 ( 
.A1(n_885),
.A2(n_847),
.B1(n_835),
.B2(n_853),
.C(n_870),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_876),
.B(n_875),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_878),
.A2(n_869),
.B1(n_851),
.B2(n_765),
.Y(n_893)
);

OAI221xp5_ASAP7_75t_L g894 ( 
.A1(n_880),
.A2(n_851),
.B1(n_827),
.B2(n_857),
.C(n_871),
.Y(n_894)
);

OAI221xp5_ASAP7_75t_L g895 ( 
.A1(n_874),
.A2(n_851),
.B1(n_857),
.B2(n_862),
.C(n_868),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_872),
.B(n_854),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_877),
.B(n_851),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_872),
.B(n_859),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_892),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_898),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_891),
.B(n_884),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_896),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_SL g903 ( 
.A1(n_891),
.A2(n_834),
.B(n_878),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_897),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_895),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_893),
.A2(n_775),
.B1(n_834),
.B2(n_842),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_890),
.B(n_878),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_899),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_903),
.A2(n_901),
.B1(n_906),
.B2(n_905),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_900),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_904),
.A2(n_894),
.B(n_881),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_907),
.B(n_902),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_909),
.B(n_888),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_908),
.B(n_906),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_912),
.B(n_882),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_910),
.Y(n_916)
);

INVx8_ASAP7_75t_L g917 ( 
.A(n_916),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_915),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_914),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_913),
.B(n_911),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_916),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_921),
.B(n_881),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_920),
.B(n_888),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_SL g924 ( 
.A(n_919),
.B(n_792),
.C(n_886),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_L g925 ( 
.A(n_918),
.B(n_917),
.C(n_799),
.Y(n_925)
);

NOR2x1_ASAP7_75t_L g926 ( 
.A(n_917),
.B(n_879),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_921),
.B(n_889),
.Y(n_927)
);

NAND2x1_ASAP7_75t_SL g928 ( 
.A(n_921),
.B(n_889),
.Y(n_928)
);

XNOR2xp5_ASAP7_75t_L g929 ( 
.A(n_924),
.B(n_795),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_926),
.A2(n_887),
.B(n_883),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_923),
.A2(n_887),
.B(n_883),
.C(n_873),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_927),
.Y(n_932)
);

AOI221xp5_ASAP7_75t_L g933 ( 
.A1(n_925),
.A2(n_873),
.B1(n_866),
.B2(n_826),
.C(n_832),
.Y(n_933)
);

OAI221xp5_ASAP7_75t_SL g934 ( 
.A1(n_928),
.A2(n_833),
.B1(n_866),
.B2(n_829),
.C(n_824),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_932),
.B(n_922),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_929),
.A2(n_856),
.B1(n_805),
.B2(n_823),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_933),
.Y(n_937)
);

XNOR2xp5_ASAP7_75t_L g938 ( 
.A(n_930),
.B(n_823),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_L g939 ( 
.A(n_934),
.B(n_829),
.C(n_824),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_SL g940 ( 
.A(n_937),
.B(n_931),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_935),
.B(n_856),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_936),
.B(n_833),
.C(n_830),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_SL g943 ( 
.A(n_938),
.B(n_831),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_R g944 ( 
.A(n_939),
.B(n_741),
.Y(n_944)
);

OAI321xp33_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_830),
.A3(n_707),
.B1(n_714),
.B2(n_711),
.C(n_713),
.Y(n_945)
);

NOR4xp25_ASAP7_75t_L g946 ( 
.A(n_940),
.B(n_733),
.C(n_736),
.D(n_741),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_943),
.A2(n_732),
.B1(n_741),
.B2(n_733),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_944),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_942),
.A2(n_733),
.B1(n_736),
.B2(n_725),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_948),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_947),
.Y(n_951)
);

NOR2x1p5_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_733),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_950),
.Y(n_953)
);

NAND2x1_ASAP7_75t_SL g954 ( 
.A(n_952),
.B(n_949),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_953),
.A2(n_951),
.B1(n_945),
.B2(n_736),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_954),
.A2(n_724),
.B1(n_725),
.B2(n_713),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_955),
.A2(n_725),
.B1(n_724),
.B2(n_753),
.Y(n_957)
);

NAND4xp25_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_725),
.C(n_724),
.D(n_715),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_955),
.A2(n_753),
.B(n_724),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_714),
.B1(n_707),
.B2(n_711),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_SL g961 ( 
.A1(n_959),
.A2(n_957),
.B1(n_709),
.B2(n_715),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_959),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_962),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_960),
.Y(n_964)
);

AOI221xp5_ASAP7_75t_L g965 ( 
.A1(n_963),
.A2(n_961),
.B1(n_715),
.B2(n_703),
.C(n_709),
.Y(n_965)
);

AOI211xp5_ASAP7_75t_L g966 ( 
.A1(n_965),
.A2(n_964),
.B(n_703),
.C(n_721),
.Y(n_966)
);


endmodule