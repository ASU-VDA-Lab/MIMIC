module fake_jpeg_13585_n_470 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_470);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_470;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_47),
.Y(n_144)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_48),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_52),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_32),
.Y(n_53)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_64),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_28),
.A2(n_15),
.B(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_63),
.B(n_70),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_15),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_66),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_11),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_11),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

BUFx12f_ASAP7_75t_SL g80 ( 
.A(n_36),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_87),
.B(n_90),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_93),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_37),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_39),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_37),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_117),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_103),
.B(n_106),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_41),
.B1(n_29),
.B2(n_18),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_104),
.A2(n_115),
.B1(n_129),
.B2(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_41),
.B1(n_18),
.B2(n_33),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_20),
.C(n_1),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_119),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_17),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_24),
.B1(n_39),
.B2(n_26),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_86),
.B1(n_84),
.B2(n_83),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_31),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_47),
.A2(n_24),
.B1(n_17),
.B2(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_49),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_51),
.B(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_31),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_1),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_60),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_3),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_55),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_72),
.B1(n_67),
.B2(n_77),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_57),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_0),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_163),
.Y(n_207)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_152),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_154),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_155),
.A2(n_171),
.B1(n_191),
.B2(n_101),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

BUFx16f_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_158),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_66),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_66),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_122),
.B1(n_101),
.B2(n_102),
.Y(n_217)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_176),
.Y(n_211)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_5),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_180),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_178)
);

AO21x2_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_121),
.B(n_108),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_141),
.B1(n_133),
.B2(n_132),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_179),
.A2(n_153),
.B(n_159),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_187),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_1),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_186),
.C(n_199),
.Y(n_208)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_197),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_100),
.B(n_2),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_95),
.B(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_136),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_195),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_110),
.B(n_4),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_5),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_103),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_106),
.Y(n_232)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_201),
.Y(n_240)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_149),
.B(n_140),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_205),
.A2(n_236),
.B1(n_239),
.B2(n_112),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_123),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_231),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_217),
.A2(n_228),
.B1(n_244),
.B2(n_204),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_164),
.A2(n_179),
.B(n_171),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_154),
.B(n_199),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_222),
.B(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_160),
.B(n_96),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_160),
.A2(n_114),
.B1(n_123),
.B2(n_138),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_114),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_153),
.B(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_249),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_191),
.B1(n_166),
.B2(n_154),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_245),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g243 ( 
.A1(n_162),
.A2(n_197),
.A3(n_151),
.B1(n_159),
.B2(n_94),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_162),
.A2(n_138),
.B1(n_122),
.B2(n_148),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_102),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_162),
.B(n_128),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_192),
.B(n_199),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_186),
.B(n_163),
.C(n_180),
.Y(n_256)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_212),
.Y(n_318)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_225),
.A2(n_170),
.B(n_175),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_260),
.A2(n_268),
.B(n_248),
.Y(n_332)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_173),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_263),
.B(n_270),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_178),
.B(n_193),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_265),
.A2(n_289),
.B(n_291),
.Y(n_300)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_266),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_209),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_269),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_225),
.A2(n_172),
.B(n_178),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_209),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_276),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_157),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_272),
.B(n_274),
.Y(n_331)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_210),
.B(n_169),
.Y(n_274)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_205),
.A2(n_178),
.B1(n_125),
.B2(n_148),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_293),
.B1(n_228),
.B2(n_232),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_216),
.B(n_196),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_287),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_217),
.A2(n_148),
.B1(n_125),
.B2(n_127),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_285),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_205),
.A2(n_127),
.B1(n_125),
.B2(n_165),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_205),
.A2(n_127),
.B1(n_201),
.B2(n_152),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_157),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_286),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_283),
.Y(n_299)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_205),
.A2(n_226),
.B1(n_213),
.B2(n_244),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_209),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_234),
.B(n_109),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_294),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_226),
.B(n_109),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_219),
.A2(n_195),
.B(n_119),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_246),
.B(n_240),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_183),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_213),
.A2(n_202),
.B1(n_184),
.B2(n_156),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_240),
.B1(n_247),
.B2(n_233),
.Y(n_325)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_207),
.B(n_116),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_218),
.Y(n_323)
);

NAND2x1p5_ASAP7_75t_R g297 ( 
.A(n_268),
.B(n_249),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_297),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_243),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_320),
.C(n_253),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_301),
.A2(n_304),
.B1(n_310),
.B2(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_235),
.B1(n_239),
.B2(n_208),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_305),
.B(n_318),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_285),
.A2(n_235),
.B1(n_231),
.B2(n_223),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_307),
.A2(n_313),
.B1(n_325),
.B2(n_267),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_278),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_326),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_208),
.B1(n_212),
.B2(n_206),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_281),
.A2(n_224),
.B1(n_220),
.B2(n_222),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_264),
.A2(n_211),
.B(n_206),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_322),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_242),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_323),
.B(n_270),
.Y(n_337)
);

AOI22x1_ASAP7_75t_L g324 ( 
.A1(n_264),
.A2(n_233),
.B1(n_215),
.B2(n_246),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_275),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_289),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_261),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_264),
.A2(n_247),
.B1(n_241),
.B2(n_248),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_260),
.A2(n_221),
.B(n_247),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_332),
.B(n_291),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_337),
.B(n_344),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_255),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_349),
.C(n_354),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_341),
.A2(n_345),
.B1(n_358),
.B2(n_360),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_342),
.B(n_297),
.Y(n_380)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_317),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_316),
.A2(n_290),
.B1(n_286),
.B2(n_269),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_307),
.B(n_288),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_346),
.B(n_348),
.Y(n_376)
);

XOR2x2_ASAP7_75t_SL g347 ( 
.A(n_298),
.B(n_256),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_318),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_312),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_315),
.Y(n_349)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_357),
.Y(n_366)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_263),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_331),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_364),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_254),
.C(n_261),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_362),
.C(n_329),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_301),
.A2(n_280),
.B1(n_265),
.B2(n_271),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_300),
.B(n_254),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_363),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_309),
.A2(n_291),
.B1(n_289),
.B2(n_262),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_361),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_303),
.B(n_274),
.C(n_287),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_304),
.A2(n_259),
.B1(n_292),
.B2(n_258),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_326),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_341),
.A2(n_310),
.B1(n_332),
.B2(n_308),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_369),
.A2(n_338),
.B1(n_357),
.B2(n_334),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_319),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_374),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_313),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_372),
.B(n_375),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_319),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_259),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_389),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_383),
.Y(n_407)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_330),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_327),
.C(n_300),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_386),
.C(n_362),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_322),
.C(n_324),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_309),
.B(n_324),
.Y(n_387)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_387),
.Y(n_393)
);

AOI21xp33_ASAP7_75t_L g388 ( 
.A1(n_339),
.A2(n_309),
.B(n_299),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_388),
.B(n_390),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_328),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_299),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_409),
.C(n_383),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_392),
.A2(n_403),
.B1(n_377),
.B2(n_365),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_335),
.Y(n_394)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_338),
.C(n_350),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_402),
.C(n_408),
.Y(n_415)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_350),
.C(n_345),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_382),
.A2(n_339),
.B1(n_358),
.B2(n_359),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_406),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_353),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_405),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_343),
.B(n_360),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_333),
.C(n_314),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_333),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_410),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_414),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_403),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_413)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_413),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_393),
.A2(n_385),
.B1(n_365),
.B2(n_369),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_389),
.C(n_380),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_427),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_386),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_395),
.C(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_424),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_392),
.A2(n_378),
.B1(n_384),
.B2(n_381),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_379),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_330),
.C(n_306),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_409),
.C(n_391),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_429),
.B(n_430),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_416),
.A2(n_405),
.B(n_398),
.C(n_406),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_431),
.A2(n_424),
.B1(n_423),
.B2(n_418),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_395),
.C(n_411),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_437),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_414),
.A2(n_401),
.B(n_411),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_434),
.A2(n_436),
.B(n_439),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_415),
.A2(n_276),
.B(n_294),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_306),
.C(n_273),
.Y(n_437)
);

AO21x1_ASAP7_75t_L g439 ( 
.A1(n_426),
.A2(n_321),
.B(n_284),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_425),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_427),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_443),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_438),
.A2(n_422),
.B1(n_419),
.B2(n_421),
.Y(n_444)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_444),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_431),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_447),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_412),
.C(n_417),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_451),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_284),
.B1(n_266),
.B2(n_241),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_SL g452 ( 
.A1(n_449),
.A2(n_439),
.B(n_433),
.C(n_435),
.Y(n_452)
);

AOI31xp67_ASAP7_75t_L g461 ( 
.A1(n_452),
.A2(n_442),
.A3(n_241),
.B(n_149),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_10),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_321),
.B(n_116),
.Y(n_458)
);

OAI221xp5_ASAP7_75t_L g459 ( 
.A1(n_458),
.A2(n_446),
.B1(n_443),
.B2(n_444),
.C(n_451),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_461),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_448),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_460),
.A2(n_462),
.B(n_455),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_463),
.B(n_464),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_460),
.A2(n_457),
.B(n_454),
.Y(n_464)
);

OAI311xp33_ASAP7_75t_L g467 ( 
.A1(n_465),
.A2(n_452),
.A3(n_7),
.B1(n_8),
.C1(n_9),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_6),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_466),
.B(n_7),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_7),
.Y(n_470)
);


endmodule