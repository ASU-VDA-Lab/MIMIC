module fake_ariane_2819_n_4410 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_478, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_17, n_225, n_235, n_464, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_4410);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_478;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_4410;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4030;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_3619;
wire n_589;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_4342;
wire n_691;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_610;
wire n_4403;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_690;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_4178;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_3765;
wire n_2006;
wire n_4090;
wire n_952;
wire n_864;
wire n_4058;
wire n_2446;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_4363;
wire n_524;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_634;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_2238;
wire n_1503;
wire n_764;
wire n_2529;
wire n_2374;
wire n_4103;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_568;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_520;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4106;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_500;
wire n_665;
wire n_754;
wire n_4260;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_829;
wire n_4148;
wire n_1062;
wire n_738;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_4038;
wire n_4132;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_953;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_2634;
wire n_3451;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_2663;
wire n_495;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_821;
wire n_561;
wire n_770;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_507;
wire n_901;
wire n_2782;
wire n_3879;
wire n_569;
wire n_4136;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_787;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_4176;
wire n_1207;
wire n_4124;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_3948;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4147;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2391;
wire n_2332;
wire n_3828;
wire n_3975;
wire n_3073;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_4018;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3613;
wire n_3325;
wire n_2885;
wire n_661;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_3003;
wire n_2874;
wire n_4117;
wire n_533;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3739;
wire n_1230;
wire n_1840;
wire n_612;
wire n_2739;
wire n_3728;
wire n_3962;
wire n_512;
wire n_1597;
wire n_4082;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_579;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_1021;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_570;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_2909;
wire n_1416;
wire n_3554;
wire n_490;
wire n_4276;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_575;
wire n_546;
wire n_3472;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_4109;
wire n_1716;
wire n_4108;
wire n_3777;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_4115;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_652;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_1179;
wire n_4311;
wire n_3284;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_2926;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_2791;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_4378;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_2398;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_513;
wire n_1292;
wire n_1972;
wire n_2015;
wire n_1178;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_669;
wire n_1491;
wire n_931;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_619;
wire n_4130;
wire n_967;
wire n_1083;
wire n_3937;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_746;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_615;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3629;
wire n_3666;
wire n_3372;
wire n_3891;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_3046;
wire n_2921;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_3257;
wire n_650;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3727;
wire n_3700;
wire n_712;
wire n_976;
wire n_3567;
wire n_909;
wire n_4003;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2795;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_799;
wire n_3884;
wire n_1147;
wire n_2829;
wire n_4367;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_965;
wire n_1914;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_646;
wire n_4254;
wire n_2507;
wire n_4219;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1234;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_3661;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_564;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_3971;
wire n_4315;
wire n_706;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_4207;
wire n_4201;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_3994;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_4049;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_4263;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3876;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4089;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_1198;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_4138;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_855;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_600;
wire n_1053;
wire n_1609;
wire n_3118;
wire n_4072;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_4323;
wire n_529;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_3922;
wire n_502;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_3599;
wire n_3618;
wire n_604;
wire n_677;
wire n_3705;
wire n_3022;
wire n_3983;
wire n_703;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_681;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_707;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_3788;
wire n_3939;
wire n_727;
wire n_699;
wire n_2075;
wire n_590;
wire n_1726;
wire n_3263;
wire n_3569;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3837;
wire n_3835;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_3819;
wire n_3761;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_4348;
wire n_688;
wire n_3139;
wire n_636;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_887;
wire n_729;
wire n_3403;
wire n_4261;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_627;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_957;
wire n_1402;
wire n_1242;
wire n_3957;
wire n_2774;
wire n_2754;
wire n_2707;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_877;
wire n_3995;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_527;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2949;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_3896;
wire n_4067;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_551;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1711;
wire n_1219;
wire n_4387;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_2594;
wire n_1239;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_560;
wire n_890;
wire n_4324;
wire n_842;
wire n_3626;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_4396;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_4114;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_837;
wire n_812;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_509;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3208;
wire n_3161;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4351;
wire n_3340;
wire n_4192;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_624;
wire n_3507;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_3864;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_4050;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_4306;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_602;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_805;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_695;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_4289;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2723;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_3925;
wire n_2928;
wire n_1118;
wire n_943;
wire n_678;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_961;
wire n_1807;
wire n_1046;
wire n_726;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_771;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3640;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_686;
wire n_4279;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_4330;
wire n_1130;
wire n_1450;
wire n_4152;
wire n_3718;
wire n_756;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_3017;
wire n_2320;
wire n_3140;
wire n_979;
wire n_2329;
wire n_2570;
wire n_2986;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2890;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2813;
wire n_515;
wire n_3381;
wire n_807;
wire n_3455;
wire n_3736;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_3605;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4404;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_4377;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_594;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4301;
wire n_3573;
wire n_2203;
wire n_2076;
wire n_2133;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_3291;
wire n_3654;
wire n_4188;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_4140;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_3982;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_4202;
wire n_2044;
wire n_928;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_3769;
wire n_4078;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_3055;
wire n_2854;
wire n_1291;
wire n_562;
wire n_4070;
wire n_2020;
wire n_748;
wire n_3987;
wire n_2310;
wire n_510;
wire n_4249;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_4139;
wire n_914;
wire n_689;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_2177;
wire n_1511;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_644;
wire n_3462;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_588;
wire n_3358;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4368;
wire n_3444;
wire n_4370;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_4091;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_667;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_4184;
wire n_846;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_2935;
wire n_4246;
wire n_715;
wire n_889;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1066;
wire n_1549;
wire n_4355;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_685;
wire n_911;
wire n_4061;
wire n_2658;
wire n_623;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_4155;
wire n_810;
wire n_3376;
wire n_4278;
wire n_1290;
wire n_1959;
wire n_3770;
wire n_3497;
wire n_617;
wire n_4375;
wire n_2396;
wire n_3243;
wire n_543;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_2692;
wire n_683;
wire n_601;
wire n_565;
wire n_3927;
wire n_628;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_743;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_3790;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_4241;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_639;
wire n_673;
wire n_3251;
wire n_3288;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_571;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3904;
wire n_3887;
wire n_593;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_526;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_3836;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_4366;
wire n_1157;
wire n_1584;
wire n_4384;
wire n_848;
wire n_1664;
wire n_3481;
wire n_629;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_4210;
wire n_532;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_540;
wire n_2624;
wire n_692;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_3926;
wire n_4209;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_4004;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_621;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_697;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_622;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3751;
wire n_4388;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_4110;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_4217;
wire n_530;
wire n_1785;
wire n_1262;
wire n_792;
wire n_4271;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_580;
wire n_3664;
wire n_1579;
wire n_494;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_3873;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_508;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_558;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_4053;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_581;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_4105;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_1630;
wire n_679;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_663;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_3897;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_3360;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_765;
wire n_2787;
wire n_4092;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_4057;
wire n_2770;
wire n_631;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_898;
wire n_857;
wire n_3042;
wire n_968;
wire n_1067;
wire n_4144;
wire n_4335;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_633;
wire n_900;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_761;
wire n_2212;
wire n_733;
wire n_3838;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_2897;
wire n_4339;
wire n_1322;
wire n_3273;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_4300;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_4064;
wire n_504;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_3970;
wire n_4371;
wire n_778;
wire n_2351;
wire n_1619;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_4080;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_3898;
wire n_2541;
wire n_694;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_4295;
wire n_3932;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_671;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_4087;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1409;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_4238;
wire n_904;
wire n_505;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_498;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_4397;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_539;
wire n_1150;
wire n_4266;
wire n_977;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_4373;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_4407;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_4165;
wire n_4154;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_4380;
wire n_4361;
wire n_3941;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4258;
wire n_2846;
wire n_4298;
wire n_3371;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_4250;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_881;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1477;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_4211;
wire n_3094;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_4408;
wire n_1983;
wire n_1273;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_4036;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_3918;
wire n_716;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_3244;
wire n_4383;
wire n_3499;
wire n_4391;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_4095;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_656;
wire n_492;
wire n_574;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3293;
wire n_3361;
wire n_4287;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3779;
wire n_3895;
wire n_3149;
wire n_537;
wire n_1063;
wire n_3934;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_4338;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_583;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_626;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_946;
wire n_3058;
wire n_757;
wire n_2047;
wire n_2792;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_3986;
wire n_2269;
wire n_1474;
wire n_2081;
wire n_937;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3894;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_4120;
wire n_4149;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2880;
wire n_2819;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4222;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_548;
wire n_3427;
wire n_2336;
wire n_523;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3430;
wire n_3483;
wire n_3249;
wire n_4046;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_390),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_148),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_260),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_295),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_147),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_304),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_370),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_42),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_452),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_476),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_424),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_175),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_22),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_325),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_371),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_402),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_262),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_412),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_209),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_306),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_114),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_44),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_386),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_143),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_248),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_250),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_420),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_286),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_387),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_189),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_187),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_69),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_82),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_288),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_152),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_149),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_221),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_264),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_408),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_462),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_467),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_57),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_161),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_466),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_248),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_132),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_174),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_487),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_448),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_320),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_252),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_255),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_21),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_329),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_307),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_36),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_230),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_2),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_344),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_2),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_64),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_40),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_124),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_245),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_295),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_11),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_339),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_249),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_103),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_67),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_472),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_52),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_97),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_212),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_300),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_436),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_63),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_377),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_47),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_82),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_433),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_211),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_45),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_89),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_303),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_367),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_33),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_128),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_58),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_355),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_24),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_481),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_357),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_187),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_260),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_403),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_74),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_324),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_368),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_236),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_226),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_482),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_300),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_484),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_421),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_362),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_156),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_410),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_348),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_324),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_196),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_16),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_451),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_431),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_68),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_325),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_326),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_454),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_332),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_209),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_303),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_291),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_192),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_486),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_369),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_373),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_393),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_284),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_168),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_129),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_61),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_81),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_396),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_257),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_327),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_374),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_201),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_309),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_99),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_239),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_228),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_428),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_8),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_77),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_56),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_157),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_249),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_13),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_246),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_228),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_214),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_115),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_1),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_139),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_123),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_4),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_185),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_381),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_345),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_477),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_163),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_455),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_392),
.Y(n_655)
);

BUFx5_ASAP7_75t_L g656 ( 
.A(n_153),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_22),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_51),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_102),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_63),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_268),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_470),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_322),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_69),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_269),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_430),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_335),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_14),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_24),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_270),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_138),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_222),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_14),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_323),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_88),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_247),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_425),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_326),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_85),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_398),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_42),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_315),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_31),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_213),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_465),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_111),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_52),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_206),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_169),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_351),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_144),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_39),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_351),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_328),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_203),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_190),
.Y(n_696)
);

CKINVDCx16_ASAP7_75t_R g697 ( 
.A(n_473),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_208),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_171),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_273),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_46),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_457),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_440),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_161),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_426),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_331),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_93),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_180),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_322),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_293),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_334),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_169),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_365),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_384),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_261),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_434),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_296),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_280),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_168),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_405),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_419),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_335),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_280),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_262),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_304),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_76),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_223),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_346),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_264),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_138),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_100),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_162),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_172),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_99),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_156),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_267),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_313),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_188),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_66),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_311),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_74),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_162),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_347),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_350),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_41),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_459),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_89),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_355),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_210),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_345),
.Y(n_750)
);

BUFx10_ASAP7_75t_L g751 ( 
.A(n_226),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_17),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_7),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_17),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_263),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_435),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_244),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_229),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_230),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_284),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_263),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_93),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_214),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_194),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_36),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_480),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_328),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_21),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_70),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_246),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_198),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_281),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_438),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_307),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_404),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_90),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_235),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_137),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_51),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_446),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_175),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_315),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_255),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_359),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_278),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_91),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_163),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_118),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_339),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_233),
.Y(n_790)
);

CKINVDCx11_ASAP7_75t_R g791 ( 
.A(n_221),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_35),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_330),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_483),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_274),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_445),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_185),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_314),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_439),
.Y(n_799)
);

CKINVDCx16_ASAP7_75t_R g800 ( 
.A(n_691),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_656),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_656),
.Y(n_802)
);

INVxp33_ASAP7_75t_SL g803 ( 
.A(n_568),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_791),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_641),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_656),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_656),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_641),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_656),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_656),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_548),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_656),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_656),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_656),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_497),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_658),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_497),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_501),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_501),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_505),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_505),
.Y(n_821)
);

INVxp33_ASAP7_75t_SL g822 ( 
.A(n_606),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_658),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_654),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_591),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_507),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_507),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_514),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_548),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_514),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_532),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_795),
.Y(n_832)
);

CKINVDCx16_ASAP7_75t_R g833 ( 
.A(n_691),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_591),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_532),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_535),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_535),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_731),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_562),
.Y(n_839)
);

INVxp33_ASAP7_75t_SL g840 ( 
.A(n_731),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_655),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_562),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_713),
.Y(n_843)
);

INVxp33_ASAP7_75t_L g844 ( 
.A(n_493),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_569),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_591),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_548),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_493),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_569),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_596),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_596),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_605),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_521),
.Y(n_853)
);

INVxp33_ASAP7_75t_L g854 ( 
.A(n_498),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_605),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_611),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_611),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_720),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_720),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_746),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_746),
.Y(n_861)
);

CKINVDCx16_ASAP7_75t_R g862 ( 
.A(n_509),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_756),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_491),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_756),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_526),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_526),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_615),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_548),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_509),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_714),
.Y(n_871)
);

INVxp33_ASAP7_75t_SL g872 ( 
.A(n_492),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_615),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_494),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_548),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_615),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_642),
.Y(n_877)
);

CKINVDCx14_ASAP7_75t_R g878 ( 
.A(n_652),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_642),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_548),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_495),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_528),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_526),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_620),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_608),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_558),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_608),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_608),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_502),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_642),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_644),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_644),
.Y(n_892)
);

INVxp33_ASAP7_75t_L g893 ( 
.A(n_498),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_652),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_670),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_670),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_670),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_707),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_707),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_586),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_707),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_712),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_712),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_712),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_727),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_508),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_644),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_516),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_664),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_727),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_664),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_664),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_620),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_690),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_620),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_727),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_620),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_620),
.Y(n_918)
);

INVxp33_ASAP7_75t_SL g919 ( 
.A(n_517),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_690),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_690),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_620),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_523),
.Y(n_923)
);

INVxp33_ASAP7_75t_SL g924 ( 
.A(n_524),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_640),
.Y(n_925)
);

INVxp33_ASAP7_75t_SL g926 ( 
.A(n_527),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_640),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_640),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_640),
.Y(n_929)
);

BUFx2_ASAP7_75t_SL g930 ( 
.A(n_652),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_640),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_697),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_640),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_614),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_529),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_669),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_669),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_669),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_646),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_536),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_537),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_669),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_669),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_669),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_672),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_542),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_653),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_672),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_672),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_543),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_843),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_811),
.Y(n_952)
);

INVx6_ASAP7_75t_L g953 ( 
.A(n_894),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_825),
.B(n_534),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_929),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_894),
.B(n_697),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_894),
.B(n_878),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_811),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_840),
.A2(n_657),
.B1(n_724),
.B2(n_665),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_929),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_942),
.Y(n_961)
);

BUFx12f_ASAP7_75t_L g962 ( 
.A(n_864),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_811),
.Y(n_963)
);

AND2x2_ASAP7_75t_SL g964 ( 
.A(n_862),
.B(n_504),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_801),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_918),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_918),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_844),
.B(n_749),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_834),
.B(n_534),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_918),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_801),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_802),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_846),
.B(n_578),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_929),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_929),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_929),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_894),
.B(n_572),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_829),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_930),
.B(n_572),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_800),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_833),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_802),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_806),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_809),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_806),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_809),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_894),
.B(n_714),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_807),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_930),
.B(n_625),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_894),
.B(n_685),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_950),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_807),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_879),
.B(n_578),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_829),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_890),
.B(n_581),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_881),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_847),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_847),
.Y(n_998)
);

OAI22x1_ASAP7_75t_R g999 ( 
.A1(n_804),
.A2(n_718),
.B1(n_737),
.B2(n_708),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_869),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_894),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_894),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_810),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_898),
.B(n_581),
.Y(n_1004)
);

INVx5_ASAP7_75t_L g1005 ( 
.A(n_869),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_871),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_871),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_889),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_901),
.B(n_490),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_810),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_SL g1011 ( 
.A(n_870),
.B(n_652),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_903),
.B(n_496),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_910),
.B(n_711),
.Y(n_1013)
);

BUFx8_ASAP7_75t_L g1014 ( 
.A(n_808),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_932),
.B(n_673),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_916),
.B(n_868),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_815),
.Y(n_1017)
);

CKINVDCx16_ASAP7_75t_R g1018 ( 
.A(n_824),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_803),
.A2(n_745),
.B1(n_761),
.B2(n_742),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_822),
.A2(n_783),
.B1(n_785),
.B2(n_769),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_841),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_875),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_875),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_880),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_906),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_805),
.A2(n_700),
.B1(n_704),
.B2(n_635),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_815),
.B(n_711),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_908),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_854),
.B(n_762),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_817),
.B(n_778),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_880),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_884),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_923),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_812),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_812),
.A2(n_522),
.B(n_504),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_813),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_884),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_813),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_814),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_817),
.B(n_818),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_814),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_823),
.A2(n_574),
.B1(n_594),
.B2(n_563),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_873),
.B(n_499),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_935),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_876),
.B(n_500),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_913),
.Y(n_1046)
);

AOI22x1_ASAP7_75t_SL g1047 ( 
.A1(n_853),
.A2(n_546),
.B1(n_551),
.B2(n_545),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_SL g1048 ( 
.A1(n_882),
.A2(n_555),
.B1(n_556),
.B2(n_552),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_922),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_940),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_922),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_925),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_808),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_838),
.A2(n_778),
.B1(n_557),
.B2(n_564),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_913),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_915),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_915),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_917),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_893),
.B(n_673),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_872),
.A2(n_600),
.B1(n_632),
.B2(n_566),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_874),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_941),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_917),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_946),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_925),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_927),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_948),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_848),
.B(n_673),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_877),
.B(n_895),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_948),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_927),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_949),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_928),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_896),
.B(n_506),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_928),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_949),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_979),
.B(n_919),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_952),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_980),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1069),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1069),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_L g1082 ( 
.A(n_962),
.B(n_818),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_1071),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_961),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1006),
.B(n_819),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1040),
.B(n_819),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_951),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_952),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_951),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_961),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_963),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_980),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_R g1093 ( 
.A(n_962),
.B(n_934),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_981),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1028),
.B(n_924),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1040),
.B(n_820),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_1028),
.B(n_926),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1071),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1050),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_958),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_978),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_963),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1050),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1021),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1040),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_958),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_954),
.B(n_897),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1006),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_966),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1006),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1021),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_978),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1007),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_954),
.B(n_899),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1007),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1018),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_1014),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1014),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_991),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_R g1121 ( 
.A(n_991),
.B(n_1008),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1071),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1008),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1007),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1049),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1049),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1051),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1051),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1033),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_1014),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_968),
.B(n_820),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1052),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_968),
.B(n_821),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1033),
.Y(n_1134)
);

XOR2xp5_ASAP7_75t_L g1135 ( 
.A(n_959),
.B(n_886),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1052),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_978),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_989),
.B(n_821),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1071),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1029),
.B(n_826),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1060),
.B(n_826),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1017),
.B(n_827),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1044),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1065),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1065),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_R g1146 ( 
.A(n_1044),
.B(n_947),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1062),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_978),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_978),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1071),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1066),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1066),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1062),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_966),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1017),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_967),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1064),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1017),
.Y(n_1158)
);

INVxp33_ASAP7_75t_L g1159 ( 
.A(n_999),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_965),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1064),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_956),
.B(n_827),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1053),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1053),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_954),
.B(n_902),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_997),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_997),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_967),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_970),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_969),
.B(n_904),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1053),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_970),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1016),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_996),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_965),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1025),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1073),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_997),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_971),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_957),
.B(n_828),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_971),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1029),
.B(n_1059),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1048),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1073),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_972),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_994),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_994),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_972),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1047),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_982),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1047),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_982),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_983),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1022),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_983),
.Y(n_1195)
);

XNOR2xp5_ASAP7_75t_L g1196 ( 
.A(n_1019),
.B(n_900),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_985),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1059),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1020),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_964),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_964),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_985),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1022),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1023),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_988),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1027),
.B(n_828),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1061),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1009),
.B(n_830),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1068),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1011),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1068),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_SL g1212 ( 
.A(n_1026),
.B(n_1054),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_988),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1023),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_997),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1072),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1027),
.B(n_830),
.Y(n_1217)
);

AND2x2_ASAP7_75t_SL g1218 ( 
.A(n_969),
.B(n_522),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_997),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1042),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_969),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_992),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1015),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1012),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_973),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1043),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_973),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_992),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_973),
.B(n_993),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1003),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1003),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1010),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_993),
.B(n_831),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_998),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_993),
.B(n_905),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1010),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1034),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_995),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_998),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1034),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1031),
.Y(n_1241)
);

INVx6_ASAP7_75t_L g1242 ( 
.A(n_984),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1036),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1036),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1045),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1031),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_995),
.B(n_831),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1038),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_995),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1074),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1027),
.B(n_835),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1004),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1038),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1039),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_990),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1039),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1004),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1004),
.B(n_835),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_998),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1032),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1041),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1013),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1041),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1035),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1035),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1032),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_987),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1013),
.Y(n_1268)
);

CKINVDCx16_ASAP7_75t_R g1269 ( 
.A(n_1013),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1037),
.Y(n_1270)
);

AND3x2_ASAP7_75t_L g1271 ( 
.A(n_1030),
.B(n_816),
.C(n_699),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1037),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1055),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1055),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1030),
.B(n_836),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1063),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_998),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1063),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_998),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1030),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_977),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1072),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1072),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1072),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_974),
.A2(n_837),
.B(n_836),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1072),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1002),
.B(n_837),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1001),
.B(n_839),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1076),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1075),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1075),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1075),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1076),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1075),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1075),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_R g1296 ( 
.A(n_1000),
.B(n_939),
.Y(n_1296)
);

CKINVDCx16_ASAP7_75t_R g1297 ( 
.A(n_1002),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1001),
.B(n_839),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1000),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1076),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1076),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1001),
.B(n_842),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1076),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1279),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1077),
.B(n_832),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1229),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1229),
.B(n_1218),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1229),
.B(n_842),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1134),
.B(n_845),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1218),
.Y(n_1310)
);

BUFx4f_ASAP7_75t_L g1311 ( 
.A(n_1287),
.Y(n_1311)
);

INVxp33_ASAP7_75t_L g1312 ( 
.A(n_1146),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1175),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_1287),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1285),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1155),
.B(n_849),
.C(n_845),
.Y(n_1316)
);

INVx5_ASAP7_75t_L g1317 ( 
.A(n_1242),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1279),
.Y(n_1318)
);

INVx8_ASAP7_75t_L g1319 ( 
.A(n_1206),
.Y(n_1319)
);

BUFx4f_ASAP7_75t_L g1320 ( 
.A(n_1287),
.Y(n_1320)
);

BUFx4f_ASAP7_75t_L g1321 ( 
.A(n_1206),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1173),
.B(n_953),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1179),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1224),
.B(n_953),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1299),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1285),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1186),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1265),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1265),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1249),
.B(n_849),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1186),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1187),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1185),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1297),
.B(n_673),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1269),
.B(n_850),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1294),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1188),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1094),
.Y(n_1339)
);

INVx8_ASAP7_75t_L g1340 ( 
.A(n_1206),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1238),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1190),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1192),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1299),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1187),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1194),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1160),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1193),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1094),
.B(n_850),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1264),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1181),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1238),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1194),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1252),
.B(n_726),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1195),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1131),
.B(n_953),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1197),
.Y(n_1357)
);

AO22x2_ASAP7_75t_L g1358 ( 
.A1(n_1135),
.A2(n_852),
.B1(n_855),
.B2(n_851),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1212),
.A2(n_852),
.B1(n_855),
.B2(n_851),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1252),
.B(n_726),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1210),
.B(n_953),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1082),
.B(n_1182),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1121),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1203),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1291),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1120),
.Y(n_1366)
);

AND2x6_ASAP7_75t_L g1367 ( 
.A(n_1086),
.B(n_856),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1131),
.B(n_856),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1133),
.B(n_857),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1202),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1133),
.B(n_857),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1101),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1291),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1182),
.B(n_726),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1203),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_SL g1376 ( 
.A(n_1099),
.B(n_726),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1221),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1204),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1140),
.B(n_858),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1181),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1221),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1225),
.A2(n_859),
.B1(n_860),
.B2(n_858),
.Y(n_1382)
);

BUFx4f_ASAP7_75t_L g1383 ( 
.A(n_1206),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1225),
.A2(n_860),
.B1(n_861),
.B2(n_859),
.Y(n_1384)
);

INVxp33_ASAP7_75t_SL g1385 ( 
.A(n_1087),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1205),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1213),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1220),
.A2(n_863),
.B1(n_865),
.B2(n_861),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1222),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1230),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1230),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1101),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1198),
.B(n_561),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1198),
.B(n_749),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1262),
.B(n_863),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1204),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1214),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1262),
.B(n_1268),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1268),
.A2(n_865),
.B1(n_762),
.B2(n_749),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1116),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1140),
.B(n_984),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1208),
.B(n_984),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1228),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1207),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1079),
.B(n_565),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1086),
.B(n_984),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1231),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1116),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1214),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1241),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1209),
.B(n_749),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1241),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1246),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1227),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1232),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1158),
.B(n_683),
.C(n_672),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1246),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1096),
.B(n_984),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1260),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1260),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1294),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1301),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1220),
.A2(n_762),
.B1(n_751),
.B2(n_672),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1209),
.A2(n_779),
.B1(n_659),
.B2(n_510),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1301),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1211),
.B(n_751),
.Y(n_1426)
);

INVx5_ASAP7_75t_L g1427 ( 
.A(n_1242),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1211),
.B(n_751),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1207),
.Y(n_1429)
);

INVxp33_ASAP7_75t_L g1430 ( 
.A(n_1135),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1266),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1255),
.B(n_751),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1255),
.B(n_762),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1266),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1120),
.B(n_571),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1123),
.B(n_573),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1096),
.B(n_866),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1236),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1257),
.B(n_1217),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1273),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_SL g1441 ( 
.A(n_1087),
.B(n_582),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1233),
.B(n_986),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1247),
.B(n_986),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1106),
.A2(n_672),
.B1(n_771),
.B2(n_683),
.Y(n_1444)
);

OAI21xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1141),
.A2(n_510),
.B(n_503),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1092),
.B(n_588),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1123),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1242),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1095),
.B(n_592),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1101),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1273),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1162),
.A2(n_1280),
.B1(n_1240),
.B2(n_1243),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1217),
.B(n_866),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1101),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1267),
.A2(n_598),
.B1(n_601),
.B2(n_597),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1292),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1237),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1180),
.B(n_986),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1078),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1244),
.A2(n_610),
.B1(n_613),
.B2(n_602),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1288),
.B(n_771),
.C(n_683),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1251),
.B(n_986),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1248),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1078),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1302),
.B(n_771),
.C(n_683),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1097),
.B(n_621),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1083),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1253),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1254),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1251),
.B(n_867),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1108),
.B(n_867),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1101),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1084),
.A2(n_683),
.B1(n_771),
.B2(n_659),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1256),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1261),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1263),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1138),
.B(n_986),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1088),
.Y(n_1478)
);

OAI21xp33_ASAP7_75t_L g1479 ( 
.A1(n_1142),
.A2(n_511),
.B(n_503),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1083),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1090),
.A2(n_771),
.B1(n_683),
.B2(n_779),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1088),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1129),
.A2(n_1143),
.B1(n_1153),
.B2(n_1147),
.Y(n_1483)
);

BUFx8_ASAP7_75t_SL g1484 ( 
.A(n_1099),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1083),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1129),
.B(n_622),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1267),
.B(n_624),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1100),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1100),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1107),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1107),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1098),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1110),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1089),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1108),
.B(n_511),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1110),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1154),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1089),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1108),
.B(n_512),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1115),
.A2(n_771),
.B1(n_513),
.B2(n_515),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1154),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1156),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1296),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_SL g1504 ( 
.A(n_1115),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1156),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1113),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1115),
.B(n_512),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1172),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1143),
.B(n_1147),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_L g1510 ( 
.A(n_1091),
.B(n_626),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1172),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1165),
.B(n_883),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1098),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1153),
.B(n_627),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1098),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1177),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1113),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1177),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1242),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1184),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1184),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1165),
.B(n_513),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1165),
.A2(n_636),
.B1(n_638),
.B2(n_631),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1170),
.B(n_515),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1157),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1125),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1200),
.B(n_637),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1170),
.B(n_883),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1170),
.B(n_519),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1122),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1118),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1126),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1157),
.B(n_639),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1161),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1127),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1113),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1200),
.B(n_1201),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1122),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1235),
.A2(n_519),
.B1(n_533),
.B2(n_525),
.Y(n_1539)
);

INVx5_ASAP7_75t_L g1540 ( 
.A(n_1113),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1201),
.B(n_1226),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1226),
.B(n_643),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1235),
.B(n_525),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1270),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1245),
.B(n_645),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1128),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1122),
.Y(n_1547)
);

CKINVDCx6p67_ASAP7_75t_R g1548 ( 
.A(n_1118),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1139),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1305),
.B(n_1235),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1339),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1459),
.Y(n_1552)
);

AO22x2_ASAP7_75t_L g1553 ( 
.A1(n_1358),
.A2(n_1196),
.B1(n_1199),
.B2(n_1159),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1484),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1339),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1309),
.B(n_1161),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1319),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1319),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1309),
.B(n_1174),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1459),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1459),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1313),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1313),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1482),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1319),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1323),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1311),
.B(n_1281),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1323),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1429),
.B(n_1104),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1333),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1377),
.B(n_1245),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1307),
.B(n_1080),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1377),
.B(n_1250),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1359),
.B(n_1258),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1333),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1319),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1338),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1319),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1321),
.B(n_1139),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1482),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1340),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1359),
.B(n_1281),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1340),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1307),
.B(n_1081),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1482),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1338),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1381),
.B(n_1250),
.Y(n_1587)
);

INVx5_ASAP7_75t_L g1588 ( 
.A(n_1340),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1340),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1306),
.B(n_1275),
.Y(n_1590)
);

BUFx10_ASAP7_75t_L g1591 ( 
.A(n_1494),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1306),
.B(n_1304),
.Y(n_1592)
);

BUFx4f_ASAP7_75t_L g1593 ( 
.A(n_1363),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1304),
.B(n_1318),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1342),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1342),
.Y(n_1596)
);

NAND3x1_ASAP7_75t_L g1597 ( 
.A(n_1388),
.B(n_538),
.C(n_533),
.Y(n_1597)
);

INVx5_ASAP7_75t_L g1598 ( 
.A(n_1340),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1343),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1343),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1328),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1311),
.A2(n_1111),
.B1(n_1114),
.B2(n_1109),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1311),
.B(n_1174),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1353),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1381),
.B(n_1341),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1341),
.B(n_1199),
.Y(n_1606)
);

BUFx10_ASAP7_75t_L g1607 ( 
.A(n_1498),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1348),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1314),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_1321),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1353),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1353),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1321),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1396),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1348),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1330),
.B(n_1085),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1363),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1352),
.B(n_1176),
.Y(n_1618)
);

AO22x2_ASAP7_75t_L g1619 ( 
.A1(n_1358),
.A2(n_1196),
.B1(n_1223),
.B2(n_1130),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1365),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1355),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1396),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1355),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1471),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1357),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1383),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1357),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1396),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1397),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1352),
.B(n_1176),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1542),
.B(n_1112),
.C(n_1104),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1370),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1314),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1370),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1385),
.A2(n_1112),
.B1(n_1130),
.B2(n_1119),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1358),
.A2(n_1136),
.B1(n_1144),
.B2(n_1132),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1386),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1397),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1397),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1304),
.B(n_1103),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1451),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1383),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1451),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1451),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1310),
.B(n_1362),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1318),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1310),
.B(n_1223),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1386),
.Y(n_1648)
);

BUFx4f_ASAP7_75t_L g1649 ( 
.A(n_1548),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1387),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1310),
.B(n_1124),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1447),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1328),
.Y(n_1653)
);

NAND2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1383),
.B(n_1139),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1330),
.B(n_1145),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1310),
.B(n_1102),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1367),
.A2(n_1103),
.B1(n_1117),
.B2(n_1151),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1387),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1525),
.B(n_1163),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1388),
.A2(n_541),
.B1(n_544),
.B2(n_538),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1308),
.B(n_1152),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1398),
.B(n_1105),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1389),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1389),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1328),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1516),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1545),
.A2(n_1119),
.B1(n_1191),
.B2(n_1189),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1365),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1525),
.B(n_1163),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1367),
.A2(n_1117),
.B1(n_1298),
.B2(n_1216),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1531),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1403),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1516),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1403),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1407),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1320),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1318),
.B(n_1164),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1398),
.B(n_1271),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1328),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1534),
.A2(n_1191),
.B1(n_1189),
.B2(n_1183),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1414),
.B(n_1150),
.Y(n_1681)
);

AND2x6_ASAP7_75t_L g1682 ( 
.A(n_1328),
.B(n_1282),
.Y(n_1682)
);

NAND3x1_ASAP7_75t_L g1683 ( 
.A(n_1455),
.B(n_544),
.C(n_541),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1439),
.B(n_1164),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1516),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1314),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1308),
.B(n_1168),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1395),
.B(n_1169),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1407),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1415),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1404),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1520),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1520),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1329),
.Y(n_1694)
);

INVx5_ASAP7_75t_L g1695 ( 
.A(n_1329),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1439),
.B(n_1171),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1520),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1415),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1521),
.Y(n_1699)
);

AND2x2_ASAP7_75t_SL g1700 ( 
.A(n_1320),
.B(n_547),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1404),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1325),
.B(n_1171),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1395),
.B(n_1272),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1329),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1438),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1329),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1521),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1438),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1457),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1349),
.B(n_1093),
.Y(n_1710)
);

INVx5_ASAP7_75t_L g1711 ( 
.A(n_1329),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1314),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1457),
.Y(n_1713)
);

AO22x2_ASAP7_75t_L g1714 ( 
.A1(n_1358),
.A2(n_1325),
.B1(n_1344),
.B2(n_1432),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1320),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1349),
.B(n_1335),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1521),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1437),
.B(n_1274),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1325),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1464),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1414),
.B(n_1150),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1463),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1344),
.B(n_1150),
.Y(n_1723)
);

AOI22x1_ASAP7_75t_L g1724 ( 
.A1(n_1463),
.A2(n_1295),
.B1(n_1216),
.B2(n_1290),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1468),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1504),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1372),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1344),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1372),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1366),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1372),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1468),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1471),
.Y(n_1733)
);

AO22x2_ASAP7_75t_L g1734 ( 
.A1(n_1433),
.A2(n_549),
.B1(n_550),
.B2(n_547),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1335),
.B(n_1183),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1469),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1365),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1464),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1478),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1421),
.B(n_1216),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1478),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1471),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1489),
.Y(n_1743)
);

NAND2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1421),
.B(n_1295),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1336),
.A2(n_1295),
.B1(n_1284),
.B2(n_1286),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1437),
.B(n_1368),
.Y(n_1746)
);

OA21x2_ASAP7_75t_L g1747 ( 
.A1(n_1315),
.A2(n_1289),
.B(n_1283),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1469),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1373),
.B(n_1527),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1421),
.B(n_1148),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1369),
.B(n_1276),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1474),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1471),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1471),
.B(n_1303),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1479),
.A2(n_1278),
.B1(n_550),
.B2(n_553),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1541),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1453),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1422),
.B(n_1149),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1367),
.A2(n_1300),
.B1(n_1293),
.B2(n_1290),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1474),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1504),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1489),
.Y(n_1762)
);

OAI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1453),
.A2(n_553),
.B1(n_554),
.B2(n_549),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1487),
.B(n_885),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1475),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1373),
.B(n_1282),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1504),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1367),
.A2(n_1303),
.B1(n_1137),
.B2(n_1148),
.Y(n_1768)
);

INVx8_ASAP7_75t_L g1769 ( 
.A(n_1367),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1373),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1453),
.B(n_1167),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1453),
.B(n_1167),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1453),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1422),
.B(n_1167),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1490),
.Y(n_1775)
);

INVx5_ASAP7_75t_L g1776 ( 
.A(n_1367),
.Y(n_1776)
);

NAND3x1_ASAP7_75t_L g1777 ( 
.A(n_1455),
.B(n_559),
.C(n_554),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_SL g1778 ( 
.A(n_1376),
.B(n_1466),
.C(n_1449),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1393),
.B(n_885),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1372),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1422),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1548),
.Y(n_1782)
);

AND2x2_ASAP7_75t_SL g1783 ( 
.A(n_1337),
.B(n_559),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1537),
.B(n_1113),
.Y(n_1784)
);

AO22x2_ASAP7_75t_L g1785 ( 
.A1(n_1475),
.A2(n_570),
.B1(n_575),
.B2(n_560),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1371),
.B(n_1137),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1367),
.A2(n_1148),
.B1(n_1149),
.B2(n_1137),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1379),
.A2(n_570),
.B1(n_575),
.B2(n_560),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1425),
.B(n_1277),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1476),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1479),
.A2(n_579),
.B1(n_580),
.B2(n_576),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1476),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1490),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1372),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1456),
.B(n_1137),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1526),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1491),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1394),
.B(n_1137),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1550),
.B(n_1512),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1660),
.A2(n_1763),
.B1(n_1746),
.B2(n_1655),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1749),
.B(n_1512),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1776),
.B(n_1425),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1749),
.B(n_1528),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1553),
.A2(n_1528),
.B1(n_1532),
.B2(n_1526),
.Y(n_1804)
);

NAND2x1p5_ASAP7_75t_L g1805 ( 
.A(n_1588),
.B(n_1425),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1776),
.B(n_1337),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1716),
.B(n_1470),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1776),
.B(n_1337),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1562),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1578),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1779),
.B(n_1470),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1786),
.A2(n_1337),
.B(n_1356),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1756),
.B(n_1556),
.Y(n_1813)
);

O2A1O1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1778),
.A2(n_1483),
.B(n_1509),
.C(n_1405),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1563),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1720),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1618),
.B(n_1503),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1566),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1571),
.A2(n_1446),
.B1(n_1441),
.B2(n_1312),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1764),
.B(n_1382),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1720),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1555),
.Y(n_1822)
);

NAND2x1_ASAP7_75t_L g1823 ( 
.A(n_1676),
.B(n_1408),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1568),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1738),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1776),
.B(n_1783),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1559),
.B(n_1523),
.Y(n_1827)
);

NOR2xp67_ASAP7_75t_L g1828 ( 
.A(n_1726),
.B(n_1503),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1738),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1553),
.A2(n_1535),
.B1(n_1546),
.B2(n_1532),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1570),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1784),
.A2(n_1350),
.B(n_1452),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1582),
.B(n_1384),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1739),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1700),
.B(n_1535),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1553),
.A2(n_1445),
.B1(n_1499),
.B2(n_1495),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1575),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1701),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1577),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1618),
.A2(n_1374),
.B(n_1436),
.C(n_1435),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1586),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1660),
.A2(n_1546),
.B1(n_1543),
.B2(n_1522),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1595),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1700),
.B(n_1507),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1571),
.A2(n_1486),
.B1(n_1533),
.B2(n_1514),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1784),
.A2(n_1350),
.B(n_1324),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1785),
.A2(n_1783),
.B1(n_1619),
.B2(n_1791),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1649),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1573),
.A2(n_1523),
.B1(n_1334),
.B2(n_1424),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1596),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1661),
.B(n_1524),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1616),
.B(n_1529),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1606),
.B(n_1426),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1572),
.B(n_1539),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1739),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_L g1856 ( 
.A(n_1769),
.B(n_1336),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1572),
.B(n_1361),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1572),
.B(n_1584),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1751),
.A2(n_1350),
.B(n_1322),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1599),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1578),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_SL g1862 ( 
.A(n_1554),
.B(n_1430),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1573),
.A2(n_1428),
.B1(n_1411),
.B2(n_1360),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1630),
.B(n_1336),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_SL g1865 ( 
.A(n_1640),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1741),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1671),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1600),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1695),
.B(n_1336),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1608),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1615),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1584),
.B(n_1347),
.Y(n_1872)
);

INVxp33_ASAP7_75t_L g1873 ( 
.A(n_1587),
.Y(n_1873)
);

AND2x6_ASAP7_75t_SL g1874 ( 
.A(n_1606),
.B(n_576),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1583),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1741),
.Y(n_1876)
);

BUFx3_ASAP7_75t_L g1877 ( 
.A(n_1649),
.Y(n_1877)
);

NAND2x1p5_ASAP7_75t_L g1878 ( 
.A(n_1588),
.B(n_1347),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1785),
.A2(n_1544),
.B1(n_1445),
.B2(n_1518),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1584),
.B(n_1347),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1587),
.A2(n_1354),
.B1(n_1380),
.B2(n_1351),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1565),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1630),
.A2(n_1380),
.B1(n_1390),
.B2(n_1351),
.Y(n_1883)
);

A2O1A1Ixp33_ASAP7_75t_SL g1884 ( 
.A1(n_1662),
.A2(n_1351),
.B(n_1380),
.C(n_1347),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1551),
.Y(n_1885)
);

NOR3xp33_ASAP7_75t_L g1886 ( 
.A(n_1631),
.B(n_1510),
.C(n_1460),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1635),
.A2(n_1423),
.B1(n_1399),
.B2(n_1500),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1569),
.B(n_1544),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1743),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1718),
.A2(n_1401),
.B(n_1406),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1574),
.B(n_1351),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1621),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1610),
.B(n_1400),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1695),
.B(n_1380),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1605),
.B(n_1662),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1623),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1605),
.B(n_1390),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1769),
.B(n_1390),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1688),
.B(n_1390),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1684),
.B(n_1391),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1583),
.Y(n_1901)
);

A2O1A1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1656),
.A2(n_1391),
.B(n_1316),
.C(n_1462),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1625),
.Y(n_1903)
);

NAND2xp33_ASAP7_75t_L g1904 ( 
.A(n_1769),
.B(n_1391),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1703),
.B(n_1391),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1627),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1632),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1593),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1634),
.B(n_1316),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1565),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1743),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1785),
.A2(n_1518),
.B1(n_1331),
.B2(n_1332),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1637),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1648),
.B(n_1400),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1667),
.A2(n_661),
.B1(n_667),
.B2(n_648),
.Y(n_1915)
);

AND3x1_ASAP7_75t_L g1916 ( 
.A(n_1659),
.B(n_580),
.C(n_579),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1650),
.B(n_1400),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1624),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1658),
.B(n_1488),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1565),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1663),
.B(n_1488),
.Y(n_1921)
);

A2O1A1Ixp33_ASAP7_75t_L g1922 ( 
.A1(n_1656),
.A2(n_1418),
.B(n_1480),
.C(n_1467),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1762),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1610),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_SL g1925 ( 
.A(n_1554),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1664),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1696),
.B(n_1467),
.Y(n_1927)
);

OAI21xp33_ASAP7_75t_L g1928 ( 
.A1(n_1652),
.A2(n_675),
.B(n_668),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1710),
.B(n_887),
.Y(n_1929)
);

O2A1O1Ixp5_ASAP7_75t_L g1930 ( 
.A1(n_1740),
.A2(n_1326),
.B(n_1315),
.C(n_1402),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1672),
.B(n_1493),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1565),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1674),
.B(n_1493),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1675),
.B(n_1496),
.Y(n_1934)
);

NAND2xp33_ASAP7_75t_L g1935 ( 
.A(n_1727),
.B(n_1729),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1689),
.B(n_1690),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1762),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1698),
.B(n_1496),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1695),
.B(n_1392),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1775),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_SL g1941 ( 
.A1(n_1798),
.A2(n_1480),
.B(n_1485),
.C(n_1467),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1695),
.B(n_1392),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_SL g1943 ( 
.A(n_1671),
.B(n_1540),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1775),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1711),
.B(n_1392),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1726),
.B(n_1408),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1619),
.A2(n_1331),
.B1(n_1332),
.B2(n_1327),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1711),
.B(n_1392),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1705),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1593),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1678),
.B(n_1467),
.Y(n_1951)
);

INVx4_ASAP7_75t_L g1952 ( 
.A(n_1588),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1678),
.B(n_1480),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1708),
.B(n_1709),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1713),
.B(n_1501),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1722),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1591),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1725),
.B(n_1501),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1669),
.A2(n_1408),
.B1(n_1485),
.B2(n_1480),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1732),
.B(n_1505),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1736),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1730),
.A2(n_1408),
.B1(n_1492),
.B2(n_1485),
.Y(n_1962)
);

OR2x6_ASAP7_75t_L g1963 ( 
.A(n_1767),
.B(n_1448),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1576),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1613),
.B(n_1485),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1793),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1748),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1750),
.A2(n_1458),
.B(n_1536),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1576),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1752),
.B(n_1505),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1617),
.A2(n_1547),
.B1(n_1513),
.B2(n_1515),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1711),
.B(n_1392),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1691),
.A2(n_1513),
.B1(n_1549),
.B2(n_1515),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1567),
.A2(n_1513),
.B1(n_1549),
.B2(n_1515),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1735),
.B(n_887),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1760),
.B(n_1508),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1793),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1765),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1790),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1711),
.B(n_1454),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1792),
.B(n_1508),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_L g1982 ( 
.A(n_1727),
.B(n_1454),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1796),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1636),
.B(n_1592),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1636),
.B(n_1492),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1592),
.B(n_1492),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1797),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1797),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1613),
.B(n_1492),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1592),
.B(n_1513),
.Y(n_1990)
);

AO22x1_ASAP7_75t_L g1991 ( 
.A1(n_1782),
.A2(n_682),
.B1(n_684),
.B2(n_678),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1687),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1591),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_L g1994 ( 
.A(n_1727),
.B(n_1454),
.Y(n_1994)
);

A2O1A1Ixp33_ASAP7_75t_SL g1995 ( 
.A1(n_1798),
.A2(n_1530),
.B(n_1538),
.C(n_1515),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1757),
.B(n_1530),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1603),
.B(n_585),
.C(n_584),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_SL g1998 ( 
.A1(n_1680),
.A2(n_689),
.B1(n_692),
.B2(n_688),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1552),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1773),
.B(n_1530),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1552),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1560),
.Y(n_2002)
);

NAND2xp33_ASAP7_75t_SL g2003 ( 
.A(n_1781),
.B(n_1530),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1560),
.Y(n_2004)
);

INVxp67_ASAP7_75t_L g2005 ( 
.A(n_1766),
.Y(n_2005)
);

INVx4_ASAP7_75t_L g2006 ( 
.A(n_1588),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1626),
.B(n_1538),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1591),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1590),
.B(n_1538),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1561),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1590),
.B(n_1538),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1952),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1873),
.B(n_1676),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1918),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1816),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1895),
.B(n_1624),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_SL g2017 ( 
.A(n_1813),
.B(n_1782),
.C(n_1603),
.Y(n_2017)
);

NOR2x1_ASAP7_75t_L g2018 ( 
.A(n_1848),
.B(n_1767),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_R g2019 ( 
.A(n_1925),
.B(n_1607),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1838),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1801),
.B(n_1781),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1858),
.B(n_1626),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1822),
.Y(n_2023)
);

BUFx12f_ASAP7_75t_L g2024 ( 
.A(n_1867),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_1822),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1803),
.B(n_1742),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1809),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1821),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1847),
.A2(n_1619),
.B1(n_1714),
.B2(n_1734),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1882),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1885),
.Y(n_2031)
);

AND2x4_ASAP7_75t_SL g2032 ( 
.A(n_1946),
.B(n_1607),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_R g2033 ( 
.A(n_1877),
.B(n_1607),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1815),
.Y(n_2034)
);

NOR2x1_ASAP7_75t_L g2035 ( 
.A(n_1828),
.B(n_1620),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1992),
.B(n_1733),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1818),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1800),
.B(n_1733),
.Y(n_2038)
);

AND2x6_ASAP7_75t_L g2039 ( 
.A(n_1984),
.B(n_1576),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1957),
.Y(n_2040)
);

NAND2x1p5_ASAP7_75t_L g2041 ( 
.A(n_1893),
.B(n_1598),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1946),
.B(n_1642),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1824),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1800),
.A2(n_1597),
.B1(n_1777),
.B2(n_1683),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1831),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2005),
.A2(n_1795),
.B(n_1721),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1837),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1825),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1993),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1827),
.B(n_1594),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_SL g2051 ( 
.A(n_1813),
.B(n_696),
.C(n_693),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_2008),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1839),
.Y(n_2053)
);

NOR3xp33_ASAP7_75t_SL g2054 ( 
.A(n_1927),
.B(n_701),
.C(n_698),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1885),
.Y(n_2055)
);

OAI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_1849),
.A2(n_1657),
.B1(n_1791),
.B2(n_1755),
.C(n_1742),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1853),
.B(n_1719),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1841),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2005),
.B(n_1651),
.Y(n_2059)
);

INVx3_ASAP7_75t_SL g2060 ( 
.A(n_1908),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1829),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1882),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1946),
.B(n_1642),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_SL g2064 ( 
.A(n_1927),
.B(n_709),
.C(n_706),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1843),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1950),
.B(n_1557),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1834),
.Y(n_2067)
);

INVx4_ASAP7_75t_L g2068 ( 
.A(n_1865),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1865),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1850),
.Y(n_2070)
);

AND2x4_ASAP7_75t_SL g2071 ( 
.A(n_1893),
.B(n_1761),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1799),
.B(n_1651),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1975),
.B(n_1594),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1847),
.A2(n_1714),
.B1(n_1734),
.B2(n_1763),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1852),
.B(n_1645),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_1952),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1860),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1855),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1833),
.B(n_1645),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1811),
.B(n_1567),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1874),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_1888),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_1807),
.B(n_1929),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_1918),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_SL g2085 ( 
.A1(n_1887),
.A2(n_1714),
.B1(n_1734),
.B2(n_1820),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1924),
.B(n_1557),
.Y(n_2086)
);

BUFx8_ASAP7_75t_L g2087 ( 
.A(n_1882),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1851),
.B(n_1561),
.Y(n_2088)
);

INVxp67_ASAP7_75t_SL g2089 ( 
.A(n_1982),
.Y(n_2089)
);

OR2x2_ASAP7_75t_SL g2090 ( 
.A(n_1844),
.B(n_1761),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1835),
.B(n_1564),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1924),
.B(n_1558),
.Y(n_2092)
);

BUFx2_ASAP7_75t_L g2093 ( 
.A(n_1882),
.Y(n_2093)
);

OAI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1853),
.A2(n_1788),
.B1(n_1753),
.B2(n_1728),
.Y(n_2094)
);

BUFx12f_ASAP7_75t_L g2095 ( 
.A(n_1910),
.Y(n_2095)
);

AND2x6_ASAP7_75t_L g2096 ( 
.A(n_1910),
.B(n_1576),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_R g2097 ( 
.A(n_1862),
.B(n_1620),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_1910),
.Y(n_2098)
);

NAND2xp33_ASAP7_75t_SL g2099 ( 
.A(n_1817),
.B(n_1715),
.Y(n_2099)
);

OR2x4_ASAP7_75t_L g2100 ( 
.A(n_1900),
.B(n_1681),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1857),
.B(n_1564),
.Y(n_2101)
);

BUFx2_ASAP7_75t_L g2102 ( 
.A(n_1910),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1920),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1830),
.B(n_1594),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1920),
.Y(n_2105)
);

INVx5_ASAP7_75t_L g2106 ( 
.A(n_1898),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1866),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1868),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1870),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1871),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1892),
.Y(n_2111)
);

BUFx10_ASAP7_75t_L g2112 ( 
.A(n_1951),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1876),
.Y(n_2113)
);

CKINVDCx14_ASAP7_75t_R g2114 ( 
.A(n_1915),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1998),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1896),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_1819),
.Y(n_2117)
);

OR2x6_ASAP7_75t_L g2118 ( 
.A(n_1826),
.B(n_1558),
.Y(n_2118)
);

XNOR2xp5_ASAP7_75t_L g2119 ( 
.A(n_1916),
.B(n_1677),
.Y(n_2119)
);

BUFx10_ASAP7_75t_L g2120 ( 
.A(n_1951),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1891),
.B(n_1580),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_1985),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1830),
.B(n_1677),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1903),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1889),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1953),
.B(n_1677),
.Y(n_2126)
);

AND3x1_ASAP7_75t_L g2127 ( 
.A(n_1928),
.B(n_1647),
.C(n_1646),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_1920),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1943),
.B(n_1668),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1906),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1899),
.B(n_1580),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1920),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1911),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1953),
.B(n_1702),
.Y(n_2134)
);

NOR2x1_ASAP7_75t_R g2135 ( 
.A(n_1826),
.B(n_1640),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1907),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_1991),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1900),
.A2(n_1597),
.B1(n_1777),
.B2(n_1683),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1923),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1842),
.A2(n_1755),
.B1(n_1788),
.B2(n_1759),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1905),
.B(n_1585),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1913),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1932),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1926),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1886),
.A2(n_1640),
.B1(n_1702),
.B2(n_1647),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1963),
.B(n_1589),
.Y(n_2146)
);

INVx4_ASAP7_75t_L g2147 ( 
.A(n_1932),
.Y(n_2147)
);

INVx4_ASAP7_75t_L g2148 ( 
.A(n_1932),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1842),
.A2(n_1668),
.B1(n_1770),
.B2(n_1737),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1932),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_2006),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_1854),
.B(n_1715),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1936),
.B(n_1585),
.Y(n_2153)
);

BUFx2_ASAP7_75t_L g2154 ( 
.A(n_1964),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_1996),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_2000),
.Y(n_2156)
);

AOI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_1832),
.A2(n_1326),
.B(n_1315),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1814),
.B(n_1737),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1965),
.B(n_1770),
.Y(n_2159)
);

OR2x6_ASAP7_75t_L g2160 ( 
.A(n_1805),
.B(n_1589),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_1964),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1949),
.Y(n_2162)
);

NOR3xp33_ASAP7_75t_SL g2163 ( 
.A(n_1864),
.B(n_715),
.C(n_710),
.Y(n_2163)
);

BUFx4f_ASAP7_75t_L g2164 ( 
.A(n_1964),
.Y(n_2164)
);

BUFx3_ASAP7_75t_L g2165 ( 
.A(n_1964),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1954),
.B(n_1604),
.Y(n_2166)
);

INVx2_ASAP7_75t_SL g2167 ( 
.A(n_1969),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1956),
.Y(n_2168)
);

BUFx3_ASAP7_75t_L g2169 ( 
.A(n_1969),
.Y(n_2169)
);

NAND2x1_ASAP7_75t_L g2170 ( 
.A(n_1898),
.B(n_1682),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2009),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1969),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1961),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1967),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_1969),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_1963),
.B(n_1598),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_1886),
.A2(n_1702),
.B1(n_1772),
.B2(n_1771),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2011),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1978),
.Y(n_2179)
);

NOR2x1_ASAP7_75t_L g2180 ( 
.A(n_1963),
.B(n_1723),
.Y(n_2180)
);

NAND2xp33_ASAP7_75t_SL g2181 ( 
.A(n_1872),
.B(n_1581),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_2006),
.Y(n_2182)
);

NOR2xp67_ASAP7_75t_L g2183 ( 
.A(n_1845),
.B(n_1598),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_1965),
.B(n_1771),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1937),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1804),
.B(n_1723),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1919),
.B(n_1604),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1921),
.B(n_1611),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_1986),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1940),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_1898),
.B(n_1598),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1979),
.Y(n_2192)
);

NOR3xp33_ASAP7_75t_SL g2193 ( 
.A(n_1840),
.B(n_719),
.C(n_717),
.Y(n_2193)
);

BUFx3_ASAP7_75t_L g2194 ( 
.A(n_1805),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1983),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1823),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_1880),
.B(n_1863),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1810),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1987),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1988),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1999),
.Y(n_2201)
);

INVx5_ASAP7_75t_L g2202 ( 
.A(n_1810),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_1804),
.B(n_1723),
.Y(n_2203)
);

NAND2x1p5_ASAP7_75t_L g2204 ( 
.A(n_1861),
.B(n_1581),
.Y(n_2204)
);

AND3x1_ASAP7_75t_SL g2205 ( 
.A(n_1836),
.B(n_585),
.C(n_584),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_1861),
.B(n_1581),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_1836),
.B(n_1590),
.Y(n_2207)
);

INVx1_ASAP7_75t_SL g2208 ( 
.A(n_1990),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_1914),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1944),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_1875),
.B(n_1581),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1966),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1881),
.B(n_1681),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1875),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_R g2215 ( 
.A(n_1935),
.B(n_1609),
.Y(n_2215)
);

NOR3xp33_ASAP7_75t_SL g2216 ( 
.A(n_1897),
.B(n_723),
.C(n_722),
.Y(n_2216)
);

NOR2x1_ASAP7_75t_L g2217 ( 
.A(n_1901),
.B(n_1609),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1977),
.Y(n_2218)
);

NOR2xp67_ASAP7_75t_L g2219 ( 
.A(n_1962),
.B(n_1670),
.Y(n_2219)
);

BUFx4f_ASAP7_75t_L g2220 ( 
.A(n_1901),
.Y(n_2220)
);

AND2x2_ASAP7_75t_SL g2221 ( 
.A(n_1947),
.B(n_1856),
.Y(n_2221)
);

BUFx12f_ASAP7_75t_L g2222 ( 
.A(n_1878),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2001),
.Y(n_2223)
);

NAND3xp33_ASAP7_75t_L g2224 ( 
.A(n_1997),
.B(n_1721),
.C(n_1766),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1878),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1939),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_1959),
.B(n_1771),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_L g2228 ( 
.A(n_1883),
.B(n_1772),
.Y(n_2228)
);

OAI21xp33_ASAP7_75t_L g2229 ( 
.A1(n_1997),
.A2(n_768),
.B(n_735),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2002),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1802),
.B(n_1772),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2004),
.Y(n_2232)
);

XNOR2xp5_ASAP7_75t_L g2233 ( 
.A(n_1947),
.B(n_1579),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2010),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1931),
.B(n_1611),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1933),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1934),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1939),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1938),
.Y(n_2239)
);

BUFx2_ASAP7_75t_SL g2240 ( 
.A(n_1942),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1879),
.B(n_1754),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1955),
.B(n_1612),
.Y(n_2242)
);

NAND2xp33_ASAP7_75t_R g2243 ( 
.A(n_1917),
.B(n_1774),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_1942),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_1802),
.B(n_1754),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_2042),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_2157),
.A2(n_1930),
.B(n_1846),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2224),
.A2(n_1902),
.B(n_1922),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2027),
.Y(n_2249)
);

OAI21x1_ASAP7_75t_L g2250 ( 
.A1(n_2157),
.A2(n_1930),
.B(n_1968),
.Y(n_2250)
);

OAI21x1_ASAP7_75t_L g2251 ( 
.A1(n_2121),
.A2(n_1859),
.B(n_1812),
.Y(n_2251)
);

OAI22x1_ASAP7_75t_L g2252 ( 
.A1(n_2044),
.A2(n_603),
.B1(n_607),
.B2(n_589),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2050),
.B(n_589),
.Y(n_2253)
);

OA22x2_ASAP7_75t_L g2254 ( 
.A1(n_2138),
.A2(n_1971),
.B1(n_1973),
.B2(n_1890),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2089),
.A2(n_1994),
.B(n_1904),
.Y(n_2255)
);

NAND2x1_ASAP7_75t_L g2256 ( 
.A(n_2012),
.B(n_1682),
.Y(n_2256)
);

AOI21xp5_ASAP7_75t_L g2257 ( 
.A1(n_2089),
.A2(n_2003),
.B(n_1808),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_2042),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2055),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2073),
.B(n_603),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_2096),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2057),
.B(n_607),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2072),
.A2(n_1808),
.B(n_1806),
.Y(n_2263)
);

OAI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2117),
.A2(n_2100),
.B1(n_2197),
.B2(n_2145),
.Y(n_2264)
);

AOI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2158),
.A2(n_1948),
.B(n_1945),
.Y(n_2265)
);

AOI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2072),
.A2(n_1806),
.B(n_1884),
.Y(n_2266)
);

AOI21x1_ASAP7_75t_L g2267 ( 
.A1(n_2183),
.A2(n_1948),
.B(n_1945),
.Y(n_2267)
);

OAI21x1_ASAP7_75t_L g2268 ( 
.A1(n_2121),
.A2(n_1724),
.B(n_1747),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_2222),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2083),
.B(n_1958),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2075),
.B(n_1960),
.Y(n_2271)
);

OAI22x1_ASAP7_75t_L g2272 ( 
.A1(n_2119),
.A2(n_623),
.B1(n_629),
.B2(n_612),
.Y(n_2272)
);

OAI21x1_ASAP7_75t_SL g2273 ( 
.A1(n_2046),
.A2(n_1909),
.B(n_1970),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2075),
.B(n_1976),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_SL g2275 ( 
.A1(n_2140),
.A2(n_1789),
.B(n_1774),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2034),
.Y(n_2276)
);

BUFx4f_ASAP7_75t_L g2277 ( 
.A(n_2060),
.Y(n_2277)
);

INVxp67_ASAP7_75t_SL g2278 ( 
.A(n_2243),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2082),
.B(n_1981),
.Y(n_2279)
);

NAND2x2_ASAP7_75t_L g2280 ( 
.A(n_2020),
.B(n_2103),
.Y(n_2280)
);

INVx6_ASAP7_75t_L g2281 ( 
.A(n_2087),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2131),
.A2(n_1747),
.B(n_1326),
.Y(n_2282)
);

OAI21x1_ASAP7_75t_L g2283 ( 
.A1(n_2131),
.A2(n_1747),
.B(n_1972),
.Y(n_2283)
);

OAI21x1_ASAP7_75t_L g2284 ( 
.A1(n_2141),
.A2(n_1980),
.B(n_1972),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2140),
.A2(n_1884),
.B(n_1941),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_2141),
.A2(n_1980),
.B(n_1758),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_2097),
.Y(n_2287)
);

OAI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2213),
.A2(n_1795),
.B(n_2007),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2112),
.B(n_1989),
.Y(n_2289)
);

AO31x2_ASAP7_75t_L g2290 ( 
.A1(n_2187),
.A2(n_1602),
.A3(n_1745),
.B(n_1614),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2037),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2031),
.B(n_612),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2213),
.A2(n_1995),
.B(n_1941),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2095),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2201),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2079),
.B(n_1879),
.Y(n_2296)
);

CKINVDCx11_ASAP7_75t_R g2297 ( 
.A(n_2024),
.Y(n_2297)
);

AOI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_2059),
.A2(n_1995),
.B(n_1894),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2197),
.A2(n_2007),
.B(n_1989),
.Y(n_2299)
);

OAI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2059),
.A2(n_1758),
.B(n_1750),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2079),
.B(n_2236),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2237),
.B(n_1912),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2016),
.B(n_1912),
.Y(n_2303)
);

AOI21xp33_ASAP7_75t_L g2304 ( 
.A1(n_2094),
.A2(n_1740),
.B(n_1774),
.Y(n_2304)
);

BUFx2_ASAP7_75t_L g2305 ( 
.A(n_2087),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2016),
.B(n_1754),
.Y(n_2306)
);

A2O1A1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2193),
.A2(n_1768),
.B(n_1787),
.C(n_1974),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_2126),
.B(n_1633),
.Y(n_2308)
);

OAI21x1_ASAP7_75t_L g2309 ( 
.A1(n_2170),
.A2(n_1894),
.B(n_1869),
.Y(n_2309)
);

OAI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2094),
.A2(n_2229),
.B(n_2193),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2199),
.Y(n_2311)
);

OAI21x1_ASAP7_75t_L g2312 ( 
.A1(n_2187),
.A2(n_1869),
.B(n_1614),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2025),
.B(n_2023),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_2134),
.A2(n_1789),
.B1(n_1633),
.B2(n_1712),
.Y(n_2314)
);

OAI21x1_ASAP7_75t_L g2315 ( 
.A1(n_2188),
.A2(n_1622),
.B(n_1612),
.Y(n_2315)
);

OAI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2056),
.A2(n_1789),
.B(n_1443),
.Y(n_2316)
);

OR2x6_ASAP7_75t_L g2317 ( 
.A(n_2118),
.B(n_1601),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_2188),
.A2(n_1628),
.B(n_1622),
.Y(n_2318)
);

NAND3xp33_ASAP7_75t_SL g2319 ( 
.A(n_2115),
.B(n_728),
.C(n_725),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2239),
.B(n_2023),
.Y(n_2320)
);

A2O1A1Ixp33_ASAP7_75t_L g2321 ( 
.A1(n_2056),
.A2(n_629),
.B(n_630),
.C(n_623),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2219),
.A2(n_1442),
.B(n_1744),
.Y(n_2322)
);

OAI21x1_ASAP7_75t_L g2323 ( 
.A1(n_2235),
.A2(n_1629),
.B(n_1628),
.Y(n_2323)
);

OAI21x1_ASAP7_75t_L g2324 ( 
.A1(n_2235),
.A2(n_1638),
.B(n_1629),
.Y(n_2324)
);

AO31x2_ASAP7_75t_L g2325 ( 
.A1(n_2242),
.A2(n_1639),
.A3(n_1641),
.B(n_1638),
.Y(n_2325)
);

AOI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2159),
.A2(n_2181),
.B(n_2184),
.Y(n_2326)
);

BUFx4_ASAP7_75t_SL g2327 ( 
.A(n_2040),
.Y(n_2327)
);

OAI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2152),
.A2(n_1744),
.B(n_1416),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2231),
.B(n_1601),
.Y(n_2329)
);

BUFx2_ASAP7_75t_L g2330 ( 
.A(n_2049),
.Y(n_2330)
);

NAND2x1p5_ASAP7_75t_L g2331 ( 
.A(n_2106),
.B(n_1601),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2014),
.B(n_1697),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_2242),
.A2(n_1641),
.B(n_1639),
.Y(n_2333)
);

OAI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2152),
.A2(n_1416),
.B(n_1461),
.Y(n_2334)
);

OAI21xp5_ASAP7_75t_L g2335 ( 
.A1(n_2080),
.A2(n_1465),
.B(n_1461),
.Y(n_2335)
);

OAI21x1_ASAP7_75t_L g2336 ( 
.A1(n_2153),
.A2(n_1644),
.B(n_1643),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2200),
.Y(n_2337)
);

OAI21x1_ASAP7_75t_L g2338 ( 
.A1(n_2153),
.A2(n_1644),
.B(n_1643),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_2063),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2014),
.B(n_888),
.Y(n_2340)
);

AOI21xp33_ASAP7_75t_L g2341 ( 
.A1(n_2085),
.A2(n_2074),
.B(n_2029),
.Y(n_2341)
);

OAI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2080),
.A2(n_1465),
.B(n_1686),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2043),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2088),
.A2(n_1653),
.B(n_1601),
.Y(n_2344)
);

AOI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_2088),
.A2(n_1665),
.B(n_1653),
.Y(n_2345)
);

O2A1O1Ixp33_ASAP7_75t_L g2346 ( 
.A1(n_2114),
.A2(n_633),
.B(n_647),
.C(n_630),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2045),
.Y(n_2347)
);

BUFx12f_ASAP7_75t_L g2348 ( 
.A(n_2069),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2166),
.A2(n_2129),
.B(n_2220),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2084),
.B(n_1673),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2047),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2084),
.B(n_1673),
.Y(n_2352)
);

NAND2x1p5_ASAP7_75t_L g2353 ( 
.A(n_2106),
.B(n_1653),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2230),
.Y(n_2354)
);

OAI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_2149),
.A2(n_1712),
.B(n_1686),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2112),
.B(n_1653),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2208),
.B(n_1666),
.Y(n_2357)
);

OAI21x1_ASAP7_75t_L g2358 ( 
.A1(n_2166),
.A2(n_1685),
.B(n_1666),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2155),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2026),
.B(n_1685),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2220),
.A2(n_1679),
.B(n_1665),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2015),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2123),
.B(n_633),
.Y(n_2363)
);

AOI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2100),
.A2(n_1679),
.B(n_1665),
.Y(n_2364)
);

OAI21x1_ASAP7_75t_L g2365 ( 
.A1(n_2091),
.A2(n_1693),
.B(n_1692),
.Y(n_2365)
);

OAI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2149),
.A2(n_1682),
.B(n_1477),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2120),
.B(n_1579),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2090),
.B(n_888),
.Y(n_2368)
);

OA21x2_ASAP7_75t_L g2369 ( 
.A1(n_2038),
.A2(n_1693),
.B(n_1692),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2051),
.B(n_647),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2026),
.B(n_1707),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_L g2372 ( 
.A(n_2013),
.B(n_651),
.C(n_649),
.Y(n_2372)
);

BUFx2_ASAP7_75t_L g2373 ( 
.A(n_2052),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2036),
.B(n_1707),
.Y(n_2374)
);

AOI21x1_ASAP7_75t_L g2375 ( 
.A1(n_2021),
.A2(n_1699),
.B(n_1697),
.Y(n_2375)
);

AOI211x1_ASAP7_75t_L g2376 ( 
.A1(n_2053),
.A2(n_651),
.B(n_660),
.C(n_649),
.Y(n_2376)
);

NAND2xp33_ASAP7_75t_L g2377 ( 
.A(n_2017),
.B(n_1682),
.Y(n_2377)
);

AOI21xp5_ASAP7_75t_L g2378 ( 
.A1(n_2221),
.A2(n_1679),
.B(n_1665),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2063),
.Y(n_2379)
);

OAI21x1_ASAP7_75t_L g2380 ( 
.A1(n_2091),
.A2(n_1717),
.B(n_1699),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2058),
.Y(n_2381)
);

INVx1_ASAP7_75t_SL g2382 ( 
.A(n_2019),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2036),
.B(n_1717),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2028),
.Y(n_2384)
);

AOI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2221),
.A2(n_1694),
.B(n_1679),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2106),
.Y(n_2386)
);

AO21x1_ASAP7_75t_L g2387 ( 
.A1(n_2038),
.A2(n_892),
.B(n_891),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2048),
.Y(n_2388)
);

INVx5_ASAP7_75t_L g2389 ( 
.A(n_2096),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2120),
.B(n_1694),
.Y(n_2390)
);

INVxp67_ASAP7_75t_SL g2391 ( 
.A(n_2155),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2202),
.A2(n_1704),
.B(n_1694),
.Y(n_2392)
);

AO21x2_ASAP7_75t_L g2393 ( 
.A1(n_2101),
.A2(n_1497),
.B(n_1491),
.Y(n_2393)
);

OAI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_2216),
.A2(n_1682),
.B(n_1549),
.Y(n_2394)
);

A2O1A1Ixp33_ASAP7_75t_L g2395 ( 
.A1(n_2085),
.A2(n_2228),
.B(n_2207),
.C(n_2074),
.Y(n_2395)
);

AOI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_2202),
.A2(n_1704),
.B(n_1694),
.Y(n_2396)
);

OAI22x1_ASAP7_75t_L g2397 ( 
.A1(n_2081),
.A2(n_663),
.B1(n_671),
.B2(n_660),
.Y(n_2397)
);

OAI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2216),
.A2(n_1549),
.B(n_1547),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2164),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_2164),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_2071),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_2177),
.B(n_1654),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2156),
.B(n_663),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2127),
.B(n_1704),
.Y(n_2404)
);

OAI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2054),
.A2(n_730),
.B(n_729),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_2203),
.B(n_891),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2061),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2156),
.B(n_671),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2106),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2065),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2178),
.B(n_674),
.Y(n_2411)
);

AO21x1_ASAP7_75t_L g2412 ( 
.A1(n_2227),
.A2(n_907),
.B(n_892),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2051),
.B(n_674),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2067),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2202),
.A2(n_1706),
.B(n_1704),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2202),
.A2(n_1706),
.B(n_1727),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2070),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2078),
.Y(n_2418)
);

NAND2x1p5_ASAP7_75t_L g2419 ( 
.A(n_2180),
.B(n_1706),
.Y(n_2419)
);

BUFx10_ASAP7_75t_L g2420 ( 
.A(n_2032),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2099),
.A2(n_1706),
.B(n_1729),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2017),
.B(n_1794),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2186),
.B(n_2104),
.Y(n_2423)
);

OAI21x1_ASAP7_75t_L g2424 ( 
.A1(n_2101),
.A2(n_1502),
.B(n_1497),
.Y(n_2424)
);

AO21x1_ASAP7_75t_L g2425 ( 
.A1(n_2231),
.A2(n_909),
.B(n_907),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2137),
.B(n_676),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2178),
.B(n_676),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2226),
.B(n_1729),
.Y(n_2428)
);

OAI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2054),
.A2(n_1654),
.B1(n_1547),
.B2(n_681),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2013),
.B(n_679),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2217),
.A2(n_1731),
.B(n_1729),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2209),
.A2(n_1780),
.B(n_1731),
.Y(n_2432)
);

AO21x1_ASAP7_75t_L g2433 ( 
.A1(n_2077),
.A2(n_911),
.B(n_909),
.Y(n_2433)
);

OAI21x1_ASAP7_75t_L g2434 ( 
.A1(n_2012),
.A2(n_2151),
.B(n_2076),
.Y(n_2434)
);

AOI222xp33_ASAP7_75t_SL g2435 ( 
.A1(n_2108),
.A2(n_687),
.B1(n_681),
.B2(n_694),
.C1(n_686),
.C2(n_679),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2109),
.Y(n_2436)
);

AND2x2_ASAP7_75t_SL g2437 ( 
.A(n_2029),
.B(n_1731),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2107),
.Y(n_2438)
);

OAI22x1_ASAP7_75t_L g2439 ( 
.A1(n_2233),
.A2(n_687),
.B1(n_694),
.B2(n_686),
.Y(n_2439)
);

OAI21x1_ASAP7_75t_L g2440 ( 
.A1(n_2076),
.A2(n_1511),
.B(n_1502),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2110),
.B(n_2111),
.Y(n_2441)
);

AOI221xp5_ASAP7_75t_SL g2442 ( 
.A1(n_2116),
.A2(n_743),
.B1(n_747),
.B2(n_732),
.C(n_695),
.Y(n_2442)
);

OR2x2_ASAP7_75t_L g2443 ( 
.A(n_2124),
.B(n_911),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2064),
.B(n_695),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2130),
.B(n_732),
.Y(n_2445)
);

OAI21x1_ASAP7_75t_L g2446 ( 
.A1(n_2151),
.A2(n_1511),
.B(n_1345),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2096),
.Y(n_2447)
);

AO31x2_ASAP7_75t_L g2448 ( 
.A1(n_2113),
.A2(n_1345),
.A3(n_1346),
.B(n_1327),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2182),
.A2(n_1364),
.B(n_1346),
.Y(n_2449)
);

AOI21x1_ASAP7_75t_L g2450 ( 
.A1(n_2209),
.A2(n_2244),
.B(n_2171),
.Y(n_2450)
);

NAND2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2176),
.B(n_1731),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2135),
.A2(n_1794),
.B(n_1780),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2160),
.A2(n_1794),
.B(n_1780),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_2033),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_2226),
.B(n_1780),
.Y(n_2455)
);

NOR2xp67_ASAP7_75t_L g2456 ( 
.A(n_2068),
.B(n_1794),
.Y(n_2456)
);

OA22x2_ASAP7_75t_L g2457 ( 
.A1(n_2022),
.A2(n_747),
.B1(n_748),
.B2(n_743),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2226),
.B(n_1454),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2160),
.A2(n_1540),
.B(n_1454),
.Y(n_2459)
);

AOI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2160),
.A2(n_1540),
.B(n_1472),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2064),
.A2(n_1547),
.B(n_1472),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2136),
.Y(n_2462)
);

BUFx2_ASAP7_75t_L g2463 ( 
.A(n_2068),
.Y(n_2463)
);

OAI21x1_ASAP7_75t_SL g2464 ( 
.A1(n_2147),
.A2(n_757),
.B(n_748),
.Y(n_2464)
);

OAI21x1_ASAP7_75t_L g2465 ( 
.A1(n_2182),
.A2(n_1375),
.B(n_1364),
.Y(n_2465)
);

OAI21x1_ASAP7_75t_L g2466 ( 
.A1(n_2204),
.A2(n_1378),
.B(n_1375),
.Y(n_2466)
);

OAI21x1_ASAP7_75t_L g2467 ( 
.A1(n_2204),
.A2(n_1409),
.B(n_1378),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2125),
.Y(n_2468)
);

OAI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2163),
.A2(n_1472),
.B(n_1450),
.Y(n_2469)
);

BUFx12f_ASAP7_75t_L g2470 ( 
.A(n_2030),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2142),
.B(n_757),
.Y(n_2471)
);

OAI21x1_ASAP7_75t_L g2472 ( 
.A1(n_2198),
.A2(n_1410),
.B(n_1409),
.Y(n_2472)
);

INVxp67_ASAP7_75t_SL g2473 ( 
.A(n_2189),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2144),
.B(n_2162),
.Y(n_2474)
);

AOI21x1_ASAP7_75t_L g2475 ( 
.A1(n_2244),
.A2(n_2171),
.B(n_2189),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2168),
.B(n_758),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2173),
.B(n_758),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2238),
.B(n_1450),
.Y(n_2478)
);

OR2x6_ASAP7_75t_L g2479 ( 
.A(n_2118),
.B(n_1450),
.Y(n_2479)
);

OAI21x1_ASAP7_75t_L g2480 ( 
.A1(n_2198),
.A2(n_1412),
.B(n_1410),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2174),
.B(n_764),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2179),
.Y(n_2482)
);

AOI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2191),
.A2(n_1540),
.B(n_1517),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2238),
.B(n_1506),
.Y(n_2484)
);

BUFx12f_ASAP7_75t_L g2485 ( 
.A(n_2030),
.Y(n_2485)
);

OA22x2_ASAP7_75t_L g2486 ( 
.A1(n_2022),
.A2(n_767),
.B1(n_776),
.B2(n_764),
.Y(n_2486)
);

AOI21xp33_ASAP7_75t_L g2487 ( 
.A1(n_2210),
.A2(n_1413),
.B(n_1412),
.Y(n_2487)
);

AOI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2191),
.A2(n_1540),
.B(n_1517),
.Y(n_2488)
);

INVx3_ASAP7_75t_L g2489 ( 
.A(n_2096),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2192),
.B(n_767),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2176),
.A2(n_1540),
.B(n_1517),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2133),
.Y(n_2492)
);

AOI21x1_ASAP7_75t_SL g2493 ( 
.A1(n_2206),
.A2(n_0),
.B(n_1),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2146),
.A2(n_1506),
.B(n_1448),
.Y(n_2494)
);

AOI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2146),
.A2(n_1506),
.B(n_1448),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2195),
.B(n_776),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2060),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2212),
.Y(n_2498)
);

OAI21x1_ASAP7_75t_L g2499 ( 
.A1(n_2234),
.A2(n_2041),
.B(n_2035),
.Y(n_2499)
);

AOI21x1_ASAP7_75t_SL g2500 ( 
.A1(n_2206),
.A2(n_0),
.B(n_3),
.Y(n_2500)
);

AOI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2118),
.A2(n_1519),
.B(n_1448),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2122),
.B(n_781),
.Y(n_2502)
);

AOI21x1_ASAP7_75t_L g2503 ( 
.A1(n_2093),
.A2(n_914),
.B(n_912),
.Y(n_2503)
);

AOI21x1_ASAP7_75t_L g2504 ( 
.A1(n_2102),
.A2(n_914),
.B(n_912),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2150),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2122),
.B(n_781),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2238),
.B(n_1148),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2223),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2245),
.A2(n_2214),
.B(n_2211),
.Y(n_2509)
);

AOI221xp5_ASAP7_75t_SL g2510 ( 
.A1(n_2214),
.A2(n_797),
.B1(n_787),
.B2(n_782),
.C(n_920),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2066),
.B(n_782),
.Y(n_2511)
);

OAI21x1_ASAP7_75t_L g2512 ( 
.A1(n_2234),
.A2(n_1417),
.B(n_1413),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_2215),
.B(n_2245),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2163),
.B(n_787),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2313),
.B(n_2241),
.Y(n_2515)
);

BUFx3_ASAP7_75t_L g2516 ( 
.A(n_2330),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2497),
.Y(n_2517)
);

BUFx6f_ASAP7_75t_L g2518 ( 
.A(n_2401),
.Y(n_2518)
);

AOI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2255),
.A2(n_2257),
.B(n_2299),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2473),
.B(n_2039),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2359),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_2288),
.A2(n_2062),
.B(n_2030),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_2401),
.Y(n_2523)
);

AOI22xp33_ASAP7_75t_L g2524 ( 
.A1(n_2341),
.A2(n_2205),
.B1(n_797),
.B2(n_2039),
.Y(n_2524)
);

BUFx12f_ASAP7_75t_L g2525 ( 
.A(n_2297),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2359),
.Y(n_2526)
);

OR2x2_ASAP7_75t_L g2527 ( 
.A(n_2391),
.B(n_2240),
.Y(n_2527)
);

NOR2xp67_ASAP7_75t_L g2528 ( 
.A(n_2389),
.B(n_2147),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2296),
.B(n_2039),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2253),
.B(n_2105),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2295),
.Y(n_2531)
);

AND2x4_ASAP7_75t_L g2532 ( 
.A(n_2389),
.B(n_2039),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2277),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2295),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2301),
.B(n_2039),
.Y(n_2535)
);

INVxp67_ASAP7_75t_SL g2536 ( 
.A(n_2369),
.Y(n_2536)
);

INVx1_ASAP7_75t_SL g2537 ( 
.A(n_2287),
.Y(n_2537)
);

INVx3_ASAP7_75t_SL g2538 ( 
.A(n_2454),
.Y(n_2538)
);

INVx4_ASAP7_75t_L g2539 ( 
.A(n_2281),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2423),
.B(n_2128),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2310),
.A2(n_2205),
.B1(n_2232),
.B2(n_2185),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2311),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2497),
.Y(n_2543)
);

A2O1A1Ixp33_ASAP7_75t_L g2544 ( 
.A1(n_2321),
.A2(n_2018),
.B(n_2066),
.C(n_2086),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2303),
.B(n_2320),
.Y(n_2545)
);

BUFx2_ASAP7_75t_L g2546 ( 
.A(n_2505),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2327),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2311),
.Y(n_2548)
);

NAND2x1p5_ASAP7_75t_L g2549 ( 
.A(n_2389),
.B(n_2194),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_2389),
.B(n_2161),
.Y(n_2550)
);

CKINVDCx16_ASAP7_75t_R g2551 ( 
.A(n_2348),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2271),
.B(n_2154),
.Y(n_2552)
);

BUFx6f_ASAP7_75t_L g2553 ( 
.A(n_2470),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2274),
.B(n_2062),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2363),
.B(n_2062),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2277),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_2450),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2264),
.A2(n_2190),
.B1(n_2218),
.B2(n_2139),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2327),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2337),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2470),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2485),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2348),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2261),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2261),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2373),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2337),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2249),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2349),
.B(n_2214),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2260),
.B(n_2262),
.Y(n_2570)
);

CKINVDCx8_ASAP7_75t_R g2571 ( 
.A(n_2454),
.Y(n_2571)
);

AOI222xp33_ASAP7_75t_L g2572 ( 
.A1(n_2395),
.A2(n_738),
.B1(n_734),
.B2(n_739),
.C1(n_736),
.C2(n_733),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_2479),
.B(n_2165),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2281),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2261),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2276),
.Y(n_2576)
);

AND2x4_ASAP7_75t_L g2577 ( 
.A(n_2479),
.B(n_2169),
.Y(n_2577)
);

O2A1O1Ixp33_ASAP7_75t_L g2578 ( 
.A1(n_2321),
.A2(n_921),
.B(n_920),
.C(n_2086),
.Y(n_2578)
);

BUFx4_ASAP7_75t_R g2579 ( 
.A(n_2420),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2291),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2360),
.B(n_2098),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2371),
.B(n_2098),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2354),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2308),
.B(n_2172),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2354),
.Y(n_2585)
);

BUFx3_ASAP7_75t_L g2586 ( 
.A(n_2305),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2343),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2439),
.A2(n_921),
.B1(n_741),
.B2(n_744),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2347),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_2297),
.Y(n_2590)
);

INVx2_ASAP7_75t_SL g2591 ( 
.A(n_2281),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_R g2592 ( 
.A(n_2377),
.B(n_2096),
.Y(n_2592)
);

OR2x6_ASAP7_75t_L g2593 ( 
.A(n_2275),
.B(n_2041),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2377),
.A2(n_2143),
.B(n_2098),
.Y(n_2594)
);

INVx4_ASAP7_75t_L g2595 ( 
.A(n_2485),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2351),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2475),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2441),
.B(n_2132),
.Y(n_2598)
);

BUFx6f_ASAP7_75t_L g2599 ( 
.A(n_2420),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2293),
.A2(n_2175),
.B(n_2143),
.Y(n_2600)
);

OAI21x1_ASAP7_75t_SL g2601 ( 
.A1(n_2273),
.A2(n_2148),
.B(n_2167),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2362),
.Y(n_2602)
);

O2A1O1Ixp33_ASAP7_75t_L g2603 ( 
.A1(n_2346),
.A2(n_2248),
.B(n_2307),
.C(n_2372),
.Y(n_2603)
);

AND2x4_ASAP7_75t_L g2604 ( 
.A(n_2479),
.B(n_2317),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2447),
.Y(n_2605)
);

INVx6_ASAP7_75t_L g2606 ( 
.A(n_2420),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2362),
.Y(n_2607)
);

BUFx2_ASAP7_75t_L g2608 ( 
.A(n_2505),
.Y(n_2608)
);

INVx2_ASAP7_75t_SL g2609 ( 
.A(n_2280),
.Y(n_2609)
);

INVx2_ASAP7_75t_SL g2610 ( 
.A(n_2280),
.Y(n_2610)
);

INVx3_ASAP7_75t_L g2611 ( 
.A(n_2447),
.Y(n_2611)
);

AOI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2266),
.A2(n_2175),
.B(n_2143),
.Y(n_2612)
);

INVx1_ASAP7_75t_SL g2613 ( 
.A(n_2259),
.Y(n_2613)
);

INVx4_ASAP7_75t_L g2614 ( 
.A(n_2294),
.Y(n_2614)
);

BUFx3_ASAP7_75t_L g2615 ( 
.A(n_2382),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2381),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2384),
.Y(n_2617)
);

OR2x2_ASAP7_75t_L g2618 ( 
.A(n_2474),
.B(n_2175),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2410),
.Y(n_2619)
);

INVx3_ASAP7_75t_L g2620 ( 
.A(n_2489),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2246),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2417),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2436),
.Y(n_2623)
);

HB1xp67_ASAP7_75t_L g2624 ( 
.A(n_2369),
.Y(n_2624)
);

AOI222xp33_ASAP7_75t_L g2625 ( 
.A1(n_2395),
.A2(n_753),
.B1(n_750),
.B2(n_754),
.C1(n_752),
.C2(n_740),
.Y(n_2625)
);

BUFx2_ASAP7_75t_L g2626 ( 
.A(n_2463),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_SL g2627 ( 
.A(n_2326),
.B(n_2225),
.Y(n_2627)
);

O2A1O1Ixp33_ASAP7_75t_SL g2628 ( 
.A1(n_2289),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2384),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2298),
.B(n_2225),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2462),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2332),
.B(n_2148),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2435),
.A2(n_2092),
.B1(n_2211),
.B2(n_759),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2270),
.B(n_2225),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2482),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2246),
.Y(n_2636)
);

OAI221xp5_ASAP7_75t_L g2637 ( 
.A1(n_2442),
.A2(n_763),
.B1(n_765),
.B2(n_760),
.C(n_755),
.Y(n_2637)
);

BUFx6f_ASAP7_75t_L g2638 ( 
.A(n_2246),
.Y(n_2638)
);

OAI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2254),
.A2(n_2196),
.B1(n_772),
.B2(n_774),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2308),
.B(n_2092),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2374),
.B(n_2196),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2498),
.Y(n_2642)
);

INVxp67_ASAP7_75t_SL g2643 ( 
.A(n_2369),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2388),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2317),
.B(n_2246),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2508),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2269),
.Y(n_2647)
);

OA22x2_ASAP7_75t_L g2648 ( 
.A1(n_2252),
.A2(n_777),
.B1(n_784),
.B2(n_770),
.Y(n_2648)
);

BUFx6f_ASAP7_75t_L g2649 ( 
.A(n_2258),
.Y(n_2649)
);

BUFx2_ASAP7_75t_L g2650 ( 
.A(n_2489),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2292),
.B(n_5),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2383),
.B(n_2196),
.Y(n_2652)
);

INVx3_ASAP7_75t_SL g2653 ( 
.A(n_2269),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2272),
.A2(n_788),
.B1(n_789),
.B2(n_786),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2254),
.A2(n_792),
.B1(n_793),
.B2(n_790),
.Y(n_2655)
);

NOR2x1_ASAP7_75t_SL g2656 ( 
.A(n_2317),
.B(n_1000),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2490),
.B(n_6),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2437),
.B(n_6),
.Y(n_2658)
);

BUFx2_ASAP7_75t_L g2659 ( 
.A(n_2294),
.Y(n_2659)
);

O2A1O1Ixp33_ASAP7_75t_L g2660 ( 
.A1(n_2307),
.A2(n_931),
.B(n_936),
.C(n_933),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2340),
.Y(n_2661)
);

AOI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2285),
.A2(n_2263),
.B(n_2251),
.Y(n_2662)
);

INVxp67_ASAP7_75t_L g2663 ( 
.A(n_2404),
.Y(n_2663)
);

INVx5_ASAP7_75t_L g2664 ( 
.A(n_2258),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2247),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2388),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2407),
.Y(n_2667)
);

O2A1O1Ixp33_ASAP7_75t_L g2668 ( 
.A1(n_2430),
.A2(n_931),
.B(n_936),
.C(n_933),
.Y(n_2668)
);

INVx3_ASAP7_75t_SL g2669 ( 
.A(n_2399),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2289),
.B(n_1000),
.Y(n_2670)
);

BUFx6f_ASAP7_75t_L g2671 ( 
.A(n_2258),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2258),
.Y(n_2672)
);

INVx2_ASAP7_75t_SL g2673 ( 
.A(n_2339),
.Y(n_2673)
);

NOR2xp67_ASAP7_75t_L g2674 ( 
.A(n_2502),
.B(n_937),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2407),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2306),
.B(n_937),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2506),
.B(n_938),
.Y(n_2677)
);

AOI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2251),
.A2(n_1519),
.B(n_1419),
.Y(n_2678)
);

OAI22xp5_ASAP7_75t_L g2679 ( 
.A1(n_2314),
.A2(n_798),
.B1(n_1481),
.B2(n_1473),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2378),
.A2(n_1519),
.B(n_1419),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_2339),
.Y(n_2681)
);

BUFx2_ASAP7_75t_L g2682 ( 
.A(n_2339),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2414),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2406),
.B(n_938),
.Y(n_2684)
);

INVx3_ASAP7_75t_L g2685 ( 
.A(n_2339),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2414),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2418),
.Y(n_2687)
);

BUFx2_ASAP7_75t_L g2688 ( 
.A(n_2379),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2418),
.Y(n_2689)
);

INVx4_ASAP7_75t_L g2690 ( 
.A(n_2399),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2350),
.B(n_943),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_2426),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2438),
.Y(n_2693)
);

AOI21x1_ASAP7_75t_L g2694 ( 
.A1(n_2404),
.A2(n_944),
.B(n_943),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2352),
.B(n_944),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2438),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2437),
.B(n_7),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2379),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_2457),
.A2(n_1420),
.B1(n_1431),
.B2(n_1417),
.Y(n_2699)
);

OAI21xp5_ASAP7_75t_L g2700 ( 
.A1(n_2510),
.A2(n_945),
.B(n_1444),
.Y(n_2700)
);

AND2x4_ASAP7_75t_L g2701 ( 
.A(n_2379),
.B(n_1000),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2279),
.B(n_945),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2468),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2302),
.B(n_1024),
.Y(n_2704)
);

BUFx3_ASAP7_75t_L g2705 ( 
.A(n_2379),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2403),
.B(n_1024),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2468),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2492),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2434),
.Y(n_2709)
);

INVx2_ASAP7_75t_SL g2710 ( 
.A(n_2400),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2370),
.B(n_8),
.Y(n_2711)
);

BUFx2_ASAP7_75t_L g2712 ( 
.A(n_2329),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2408),
.B(n_1024),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2278),
.B(n_1024),
.Y(n_2714)
);

BUFx2_ASAP7_75t_L g2715 ( 
.A(n_2329),
.Y(n_2715)
);

OR2x2_ASAP7_75t_L g2716 ( 
.A(n_2368),
.B(n_1024),
.Y(n_2716)
);

BUFx6f_ASAP7_75t_L g2717 ( 
.A(n_2329),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2300),
.B(n_1046),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2413),
.B(n_9),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2492),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_2451),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2443),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2357),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_2400),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2411),
.B(n_1046),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2319),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2448),
.Y(n_2727)
);

INVx2_ASAP7_75t_SL g2728 ( 
.A(n_2511),
.Y(n_2728)
);

OAI21x1_ASAP7_75t_L g2729 ( 
.A1(n_2250),
.A2(n_1431),
.B(n_1420),
.Y(n_2729)
);

NAND2x1p5_ASAP7_75t_L g2730 ( 
.A(n_2513),
.B(n_1434),
.Y(n_2730)
);

AND3x1_ASAP7_75t_SL g2731 ( 
.A(n_2493),
.B(n_9),
.C(n_10),
.Y(n_2731)
);

OR2x6_ASAP7_75t_L g2732 ( 
.A(n_2513),
.B(n_1434),
.Y(n_2732)
);

AND2x4_ASAP7_75t_L g2733 ( 
.A(n_2509),
.B(n_1046),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2397),
.Y(n_2734)
);

AOI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2385),
.A2(n_1519),
.B(n_1440),
.Y(n_2735)
);

OR2x6_ASAP7_75t_L g2736 ( 
.A(n_2386),
.B(n_1440),
.Y(n_2736)
);

INVx3_ASAP7_75t_L g2737 ( 
.A(n_2434),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_2451),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2444),
.B(n_2514),
.Y(n_2739)
);

INVx4_ASAP7_75t_L g2740 ( 
.A(n_2419),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2386),
.B(n_1046),
.Y(n_2741)
);

AND2x4_ASAP7_75t_L g2742 ( 
.A(n_2409),
.B(n_1046),
.Y(n_2742)
);

INVx4_ASAP7_75t_L g2743 ( 
.A(n_2419),
.Y(n_2743)
);

OAI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2402),
.A2(n_520),
.B1(n_530),
.B2(n_518),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_2457),
.A2(n_1058),
.B1(n_1067),
.B2(n_1057),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2328),
.B(n_1057),
.Y(n_2746)
);

OAI21x1_ASAP7_75t_SL g2747 ( 
.A1(n_2364),
.A2(n_974),
.B(n_10),
.Y(n_2747)
);

AO21x2_ASAP7_75t_L g2748 ( 
.A1(n_2387),
.A2(n_1058),
.B(n_1057),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2325),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_2355),
.Y(n_2750)
);

NAND3xp33_ASAP7_75t_L g2751 ( 
.A(n_2376),
.B(n_1058),
.C(n_1057),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2486),
.A2(n_1058),
.B1(n_1067),
.B2(n_1057),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2325),
.Y(n_2753)
);

AOI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2402),
.A2(n_2486),
.B1(n_2367),
.B2(n_2412),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2427),
.B(n_1058),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2325),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2448),
.Y(n_2757)
);

INVxp67_ASAP7_75t_SL g2758 ( 
.A(n_2247),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2409),
.B(n_1067),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2367),
.Y(n_2760)
);

OAI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2429),
.A2(n_539),
.B1(n_540),
.B2(n_531),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2366),
.A2(n_1427),
.B(n_1317),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2448),
.Y(n_2763)
);

BUFx6f_ASAP7_75t_L g2764 ( 
.A(n_2331),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2448),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2325),
.Y(n_2766)
);

INVx4_ASAP7_75t_L g2767 ( 
.A(n_2331),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2353),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2365),
.Y(n_2769)
);

INVxp67_ASAP7_75t_SL g2770 ( 
.A(n_2250),
.Y(n_2770)
);

BUFx2_ASAP7_75t_SL g2771 ( 
.A(n_2456),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2365),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2312),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_SL g2774 ( 
.A1(n_2316),
.A2(n_577),
.B1(n_583),
.B2(n_567),
.Y(n_2774)
);

INVx4_ASAP7_75t_L g2775 ( 
.A(n_2353),
.Y(n_2775)
);

INVx5_ASAP7_75t_L g2776 ( 
.A(n_2256),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2312),
.Y(n_2777)
);

OA21x2_ASAP7_75t_L g2778 ( 
.A1(n_2662),
.A2(n_2424),
.B(n_2268),
.Y(n_2778)
);

INVx4_ASAP7_75t_L g2779 ( 
.A(n_2579),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2583),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2552),
.B(n_2445),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2521),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2526),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2568),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2520),
.B(n_2356),
.Y(n_2785)
);

OAI21x1_ASAP7_75t_L g2786 ( 
.A1(n_2662),
.A2(n_2424),
.B(n_2268),
.Y(n_2786)
);

BUFx2_ASAP7_75t_R g2787 ( 
.A(n_2547),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2552),
.B(n_2471),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2515),
.B(n_2356),
.Y(n_2789)
);

CKINVDCx20_ASAP7_75t_R g2790 ( 
.A(n_2590),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2557),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2576),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2540),
.B(n_2390),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2585),
.Y(n_2794)
);

OAI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2774),
.A2(n_2422),
.B1(n_2394),
.B2(n_2390),
.Y(n_2795)
);

OAI21x1_ASAP7_75t_L g2796 ( 
.A1(n_2519),
.A2(n_2375),
.B(n_2318),
.Y(n_2796)
);

INVxp67_ASAP7_75t_SL g2797 ( 
.A(n_2536),
.Y(n_2797)
);

OAI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2603),
.A2(n_2405),
.B(n_2422),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2545),
.B(n_2476),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2602),
.Y(n_2800)
);

OAI21x1_ASAP7_75t_SL g2801 ( 
.A1(n_2609),
.A2(n_2464),
.B(n_2265),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2580),
.Y(n_2802)
);

NAND3xp33_ASAP7_75t_L g2803 ( 
.A(n_2572),
.B(n_2625),
.C(n_2603),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2587),
.Y(n_2804)
);

OAI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2639),
.A2(n_2432),
.B(n_2428),
.Y(n_2805)
);

OAI21x1_ASAP7_75t_L g2806 ( 
.A1(n_2519),
.A2(n_2318),
.B(n_2315),
.Y(n_2806)
);

INVx5_ASAP7_75t_L g2807 ( 
.A(n_2593),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2612),
.A2(n_2446),
.B(n_2440),
.Y(n_2808)
);

AOI21x1_ASAP7_75t_L g2809 ( 
.A1(n_2557),
.A2(n_2455),
.B(n_2428),
.Y(n_2809)
);

HB1xp67_ASAP7_75t_L g2810 ( 
.A(n_2597),
.Y(n_2810)
);

AO21x1_ASAP7_75t_L g2811 ( 
.A1(n_2639),
.A2(n_2481),
.B(n_2477),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2589),
.Y(n_2812)
);

AOI22x1_ASAP7_75t_L g2813 ( 
.A1(n_2538),
.A2(n_2556),
.B1(n_2533),
.B2(n_2614),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2774),
.A2(n_2524),
.B1(n_2637),
.B2(n_2541),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2553),
.Y(n_2815)
);

O2A1O1Ixp5_ASAP7_75t_L g2816 ( 
.A1(n_2630),
.A2(n_2458),
.B(n_2455),
.C(n_2478),
.Y(n_2816)
);

OAI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2655),
.A2(n_2398),
.B(n_2334),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2596),
.Y(n_2818)
);

OAI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2660),
.A2(n_2284),
.B(n_2458),
.Y(n_2819)
);

HB1xp67_ASAP7_75t_L g2820 ( 
.A(n_2597),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2545),
.B(n_2496),
.Y(n_2821)
);

INVxp67_ASAP7_75t_L g2822 ( 
.A(n_2750),
.Y(n_2822)
);

OAI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2660),
.A2(n_2284),
.B(n_2342),
.Y(n_2823)
);

OAI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2612),
.A2(n_2446),
.B(n_2440),
.Y(n_2824)
);

OAI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2744),
.A2(n_2637),
.B(n_2522),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2554),
.B(n_2286),
.Y(n_2826)
);

OA21x2_ASAP7_75t_L g2827 ( 
.A1(n_2536),
.A2(n_2283),
.B(n_2286),
.Y(n_2827)
);

OA21x2_ASAP7_75t_L g2828 ( 
.A1(n_2643),
.A2(n_2283),
.B(n_2336),
.Y(n_2828)
);

INVx2_ASAP7_75t_SL g2829 ( 
.A(n_2586),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2616),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2607),
.Y(n_2831)
);

AOI21x1_ASAP7_75t_L g2832 ( 
.A1(n_2630),
.A2(n_2507),
.B(n_2433),
.Y(n_2832)
);

OAI21x1_ASAP7_75t_L g2833 ( 
.A1(n_2600),
.A2(n_2694),
.B(n_2678),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2617),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2619),
.Y(n_2835)
);

OAI21x1_ASAP7_75t_L g2836 ( 
.A1(n_2600),
.A2(n_2465),
.B(n_2449),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2524),
.A2(n_2425),
.B1(n_2304),
.B2(n_2335),
.Y(n_2837)
);

OAI21x1_ASAP7_75t_L g2838 ( 
.A1(n_2678),
.A2(n_2323),
.B(n_2315),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2762),
.A2(n_2459),
.B(n_2421),
.Y(n_2839)
);

INVx2_ASAP7_75t_SL g2840 ( 
.A(n_2516),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2622),
.Y(n_2841)
);

OAI21x1_ASAP7_75t_L g2842 ( 
.A1(n_2729),
.A2(n_2324),
.B(n_2323),
.Y(n_2842)
);

OAI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2541),
.A2(n_2461),
.B1(n_2469),
.B2(n_2322),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2554),
.B(n_2344),
.Y(n_2844)
);

OAI21x1_ASAP7_75t_L g2845 ( 
.A1(n_2770),
.A2(n_2333),
.B(n_2324),
.Y(n_2845)
);

AO21x2_ASAP7_75t_L g2846 ( 
.A1(n_2643),
.A2(n_2393),
.B(n_2380),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2546),
.B(n_2309),
.Y(n_2847)
);

OR2x6_ASAP7_75t_L g2848 ( 
.A(n_2532),
.B(n_2499),
.Y(n_2848)
);

OAI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2522),
.A2(n_2345),
.B(n_2507),
.Y(n_2849)
);

A2O1A1Ixp33_ASAP7_75t_L g2850 ( 
.A1(n_2578),
.A2(n_2452),
.B(n_2453),
.C(n_2460),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2754),
.A2(n_2361),
.B1(n_2431),
.B2(n_2478),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2661),
.B(n_2290),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2658),
.A2(n_2484),
.B1(n_2499),
.B2(n_2491),
.Y(n_2853)
);

OAI21x1_ASAP7_75t_L g2854 ( 
.A1(n_2762),
.A2(n_2465),
.B(n_2449),
.Y(n_2854)
);

OAI21x1_ASAP7_75t_SL g2855 ( 
.A1(n_2610),
.A2(n_2267),
.B(n_2416),
.Y(n_2855)
);

OAI21x1_ASAP7_75t_L g2856 ( 
.A1(n_2770),
.A2(n_2333),
.B(n_2336),
.Y(n_2856)
);

BUFx6f_ASAP7_75t_L g2857 ( 
.A(n_2553),
.Y(n_2857)
);

AOI21x1_ASAP7_75t_L g2858 ( 
.A1(n_2670),
.A2(n_2484),
.B(n_2503),
.Y(n_2858)
);

INVx4_ASAP7_75t_L g2859 ( 
.A(n_2606),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2623),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2608),
.B(n_2309),
.Y(n_2861)
);

OAI21x1_ASAP7_75t_L g2862 ( 
.A1(n_2680),
.A2(n_2358),
.B(n_2338),
.Y(n_2862)
);

AOI21x1_ASAP7_75t_L g2863 ( 
.A1(n_2670),
.A2(n_2504),
.B(n_2396),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_2559),
.Y(n_2864)
);

OR2x2_ASAP7_75t_L g2865 ( 
.A(n_2570),
.B(n_2290),
.Y(n_2865)
);

CKINVDCx8_ASAP7_75t_R g2866 ( 
.A(n_2551),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2640),
.B(n_2537),
.Y(n_2867)
);

AO21x2_ASAP7_75t_L g2868 ( 
.A1(n_2749),
.A2(n_2393),
.B(n_2380),
.Y(n_2868)
);

INVx3_ASAP7_75t_L g2869 ( 
.A(n_2605),
.Y(n_2869)
);

OAI21x1_ASAP7_75t_L g2870 ( 
.A1(n_2680),
.A2(n_2358),
.B(n_2338),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2665),
.Y(n_2871)
);

AOI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2746),
.A2(n_2569),
.B(n_2594),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2746),
.A2(n_2415),
.B(n_2392),
.Y(n_2873)
);

OAI21x1_ASAP7_75t_L g2874 ( 
.A1(n_2735),
.A2(n_2282),
.B(n_2500),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2629),
.Y(n_2875)
);

AO21x2_ASAP7_75t_L g2876 ( 
.A1(n_2753),
.A2(n_2487),
.B(n_2282),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2631),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2644),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2517),
.B(n_2290),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2635),
.Y(n_2880)
);

INVx6_ASAP7_75t_L g2881 ( 
.A(n_2539),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2543),
.B(n_2290),
.Y(n_2882)
);

OAI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2735),
.A2(n_2480),
.B(n_2472),
.Y(n_2883)
);

NAND2x2_ASAP7_75t_L g2884 ( 
.A(n_2566),
.B(n_11),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2626),
.B(n_12),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2598),
.B(n_12),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2518),
.Y(n_2887)
);

OAI21x1_ASAP7_75t_L g2888 ( 
.A1(n_2601),
.A2(n_2480),
.B(n_2472),
.Y(n_2888)
);

O2A1O1Ixp33_ASAP7_75t_SL g2889 ( 
.A1(n_2544),
.A2(n_2488),
.B(n_2483),
.C(n_16),
.Y(n_2889)
);

AOI21xp5_ASAP7_75t_L g2890 ( 
.A1(n_2569),
.A2(n_2501),
.B(n_2495),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2642),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_L g2892 ( 
.A1(n_2594),
.A2(n_2512),
.B(n_2467),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2666),
.Y(n_2893)
);

OAI21x1_ASAP7_75t_L g2894 ( 
.A1(n_2709),
.A2(n_2512),
.B(n_2467),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2667),
.Y(n_2895)
);

OAI21x1_ASAP7_75t_L g2896 ( 
.A1(n_2709),
.A2(n_2737),
.B(n_2747),
.Y(n_2896)
);

AO21x2_ASAP7_75t_L g2897 ( 
.A1(n_2756),
.A2(n_2466),
.B(n_2494),
.Y(n_2897)
);

AOI21x1_ASAP7_75t_L g2898 ( 
.A1(n_2714),
.A2(n_2466),
.B(n_1067),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2646),
.B(n_13),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2529),
.B(n_1067),
.Y(n_2900)
);

AOI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_2697),
.A2(n_590),
.B1(n_593),
.B2(n_587),
.Y(n_2901)
);

OA21x2_ASAP7_75t_L g2902 ( 
.A1(n_2758),
.A2(n_599),
.B(n_595),
.Y(n_2902)
);

AOI21x1_ASAP7_75t_L g2903 ( 
.A1(n_2714),
.A2(n_1056),
.B(n_1005),
.Y(n_2903)
);

BUFx2_ASAP7_75t_L g2904 ( 
.A(n_2659),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2648),
.A2(n_609),
.B1(n_616),
.B2(n_604),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2665),
.Y(n_2906)
);

OAI21x1_ASAP7_75t_L g2907 ( 
.A1(n_2737),
.A2(n_1149),
.B(n_1148),
.Y(n_2907)
);

INVxp67_ASAP7_75t_L g2908 ( 
.A(n_2618),
.Y(n_2908)
);

OAI21x1_ASAP7_75t_L g2909 ( 
.A1(n_2718),
.A2(n_1166),
.B(n_1149),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2530),
.B(n_15),
.Y(n_2910)
);

BUFx2_ASAP7_75t_L g2911 ( 
.A(n_2539),
.Y(n_2911)
);

INVx4_ASAP7_75t_L g2912 ( 
.A(n_2606),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2687),
.Y(n_2913)
);

OAI21x1_ASAP7_75t_L g2914 ( 
.A1(n_2718),
.A2(n_1166),
.B(n_1149),
.Y(n_2914)
);

INVx4_ASAP7_75t_SL g2915 ( 
.A(n_2593),
.Y(n_2915)
);

O2A1O1Ixp33_ASAP7_75t_L g2916 ( 
.A1(n_2628),
.A2(n_19),
.B(n_15),
.C(n_18),
.Y(n_2916)
);

OAI22xp33_ASAP7_75t_L g2917 ( 
.A1(n_2648),
.A2(n_618),
.B1(n_619),
.B2(n_617),
.Y(n_2917)
);

OAI21x1_ASAP7_75t_L g2918 ( 
.A1(n_2773),
.A2(n_1167),
.B(n_1166),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2696),
.Y(n_2919)
);

INVxp33_ASAP7_75t_L g2920 ( 
.A(n_2584),
.Y(n_2920)
);

NOR2x1_ASAP7_75t_SL g2921 ( 
.A(n_2593),
.B(n_955),
.Y(n_2921)
);

CKINVDCx6p67_ASAP7_75t_R g2922 ( 
.A(n_2525),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2722),
.B(n_2581),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2531),
.Y(n_2924)
);

AOI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2627),
.A2(n_1427),
.B(n_1317),
.Y(n_2925)
);

BUFx6f_ASAP7_75t_L g2926 ( 
.A(n_2553),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2720),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2520),
.B(n_18),
.Y(n_2928)
);

O2A1O1Ixp33_ASAP7_75t_SL g2929 ( 
.A1(n_2640),
.A2(n_23),
.B(n_19),
.C(n_20),
.Y(n_2929)
);

OA21x2_ASAP7_75t_L g2930 ( 
.A1(n_2758),
.A2(n_634),
.B(n_628),
.Y(n_2930)
);

AOI22xp33_ASAP7_75t_SL g2931 ( 
.A1(n_2739),
.A2(n_662),
.B1(n_666),
.B2(n_650),
.Y(n_2931)
);

OAI21x1_ASAP7_75t_SL g2932 ( 
.A1(n_2614),
.A2(n_2591),
.B(n_2574),
.Y(n_2932)
);

OAI21x1_ASAP7_75t_L g2933 ( 
.A1(n_2777),
.A2(n_1167),
.B(n_1166),
.Y(n_2933)
);

BUFx2_ASAP7_75t_SL g2934 ( 
.A(n_2571),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2542),
.Y(n_2935)
);

AOI22xp33_ASAP7_75t_L g2936 ( 
.A1(n_2588),
.A2(n_680),
.B1(n_702),
.B2(n_677),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2581),
.B(n_20),
.Y(n_2937)
);

OAI221xp5_ASAP7_75t_L g2938 ( 
.A1(n_2654),
.A2(n_716),
.B1(n_721),
.B2(n_705),
.C(n_703),
.Y(n_2938)
);

OAI22xp33_ASAP7_75t_L g2939 ( 
.A1(n_2734),
.A2(n_773),
.B1(n_775),
.B2(n_766),
.Y(n_2939)
);

NAND3xp33_ASAP7_75t_L g2940 ( 
.A(n_2663),
.B(n_2627),
.C(n_2632),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2548),
.Y(n_2941)
);

INVxp67_ASAP7_75t_L g2942 ( 
.A(n_2527),
.Y(n_2942)
);

INVx4_ASAP7_75t_L g2943 ( 
.A(n_2606),
.Y(n_2943)
);

AOI21xp33_ASAP7_75t_L g2944 ( 
.A1(n_2663),
.A2(n_794),
.B(n_780),
.Y(n_2944)
);

NAND3xp33_ASAP7_75t_L g2945 ( 
.A(n_2632),
.B(n_799),
.C(n_796),
.Y(n_2945)
);

HB1xp67_ASAP7_75t_L g2946 ( 
.A(n_2769),
.Y(n_2946)
);

INVx4_ASAP7_75t_L g2947 ( 
.A(n_2599),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2633),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2534),
.Y(n_2949)
);

INVxp67_ASAP7_75t_SL g2950 ( 
.A(n_2624),
.Y(n_2950)
);

AO21x2_ASAP7_75t_L g2951 ( 
.A1(n_2766),
.A2(n_1056),
.B(n_1005),
.Y(n_2951)
);

OAI21x1_ASAP7_75t_L g2952 ( 
.A1(n_2772),
.A2(n_1178),
.B(n_1166),
.Y(n_2952)
);

BUFx6f_ASAP7_75t_L g2953 ( 
.A(n_2553),
.Y(n_2953)
);

OAI21x1_ASAP7_75t_L g2954 ( 
.A1(n_2704),
.A2(n_1215),
.B(n_1178),
.Y(n_2954)
);

HB1xp67_ASAP7_75t_L g2955 ( 
.A(n_2624),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2588),
.A2(n_1056),
.B1(n_1070),
.B2(n_1005),
.Y(n_2956)
);

INVxp67_ASAP7_75t_L g2957 ( 
.A(n_2582),
.Y(n_2957)
);

INVx4_ASAP7_75t_L g2958 ( 
.A(n_2599),
.Y(n_2958)
);

BUFx2_ASAP7_75t_R g2959 ( 
.A(n_2563),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2560),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2567),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2582),
.B(n_25),
.Y(n_2962)
);

AOI221xp5_ASAP7_75t_L g2963 ( 
.A1(n_2654),
.A2(n_975),
.B1(n_976),
.B2(n_960),
.C(n_955),
.Y(n_2963)
);

OR2x2_ASAP7_75t_L g2964 ( 
.A(n_2529),
.B(n_2535),
.Y(n_2964)
);

OAI22x1_ASAP7_75t_L g2965 ( 
.A1(n_2692),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2675),
.Y(n_2966)
);

AO31x2_ASAP7_75t_L g2967 ( 
.A1(n_2727),
.A2(n_1056),
.A3(n_1070),
.B(n_1005),
.Y(n_2967)
);

OAI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2578),
.A2(n_1056),
.B(n_1005),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2657),
.A2(n_1070),
.B1(n_1215),
.B2(n_1178),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2683),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_2647),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2599),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2686),
.Y(n_2973)
);

A2O1A1Ixp33_ASAP7_75t_L g2974 ( 
.A1(n_2711),
.A2(n_2719),
.B(n_2651),
.C(n_2745),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2689),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2584),
.B(n_27),
.Y(n_2976)
);

AOI22xp33_ASAP7_75t_L g2977 ( 
.A1(n_2674),
.A2(n_2728),
.B1(n_2752),
.B2(n_2745),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2760),
.B(n_28),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2634),
.B(n_29),
.Y(n_2979)
);

NAND2x1p5_ASAP7_75t_L g2980 ( 
.A(n_2532),
.B(n_1317),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2693),
.Y(n_2981)
);

OAI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2761),
.A2(n_1070),
.B(n_29),
.Y(n_2982)
);

BUFx4f_ASAP7_75t_L g2983 ( 
.A(n_2538),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_2615),
.Y(n_2984)
);

INVx6_ASAP7_75t_L g2985 ( 
.A(n_2561),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2732),
.A2(n_1427),
.B(n_1317),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2712),
.B(n_2715),
.Y(n_2987)
);

CKINVDCx20_ASAP7_75t_R g2988 ( 
.A(n_2653),
.Y(n_2988)
);

BUFx2_ASAP7_75t_L g2989 ( 
.A(n_2650),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2703),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2707),
.Y(n_2991)
);

BUFx3_ASAP7_75t_L g2992 ( 
.A(n_2518),
.Y(n_2992)
);

INVx4_ASAP7_75t_L g2993 ( 
.A(n_2653),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2708),
.Y(n_2994)
);

INVx3_ASAP7_75t_L g2995 ( 
.A(n_2605),
.Y(n_2995)
);

INVx4_ASAP7_75t_L g2996 ( 
.A(n_2669),
.Y(n_2996)
);

OAI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2726),
.A2(n_2668),
.B(n_2751),
.Y(n_2997)
);

OA21x2_ASAP7_75t_L g2998 ( 
.A1(n_2757),
.A2(n_1070),
.B(n_1178),
.Y(n_2998)
);

CKINVDCx16_ASAP7_75t_R g2999 ( 
.A(n_2592),
.Y(n_2999)
);

AND2x4_ASAP7_75t_L g3000 ( 
.A(n_2604),
.B(n_30),
.Y(n_3000)
);

OAI21xp33_ASAP7_75t_L g3001 ( 
.A1(n_2535),
.A2(n_30),
.B(n_31),
.Y(n_3001)
);

OAI21x1_ASAP7_75t_L g3002 ( 
.A1(n_2704),
.A2(n_1215),
.B(n_1178),
.Y(n_3002)
);

AND2x4_ASAP7_75t_L g3003 ( 
.A(n_2604),
.B(n_32),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2803),
.A2(n_2814),
.B1(n_2837),
.B2(n_2974),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2811),
.A2(n_2558),
.B1(n_2723),
.B2(n_2555),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2999),
.B(n_2592),
.Y(n_3006)
);

NAND2xp33_ASAP7_75t_SL g3007 ( 
.A(n_2779),
.B(n_2669),
.Y(n_3007)
);

NAND3xp33_ASAP7_75t_SL g3008 ( 
.A(n_2905),
.B(n_2613),
.C(n_2730),
.Y(n_3008)
);

AND2x4_ASAP7_75t_L g3009 ( 
.A(n_2847),
.B(n_2564),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2817),
.A2(n_2558),
.B1(n_2555),
.B2(n_2699),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2809),
.A2(n_2565),
.B(n_2564),
.Y(n_3011)
);

OAI21x1_ASAP7_75t_L g3012 ( 
.A1(n_2896),
.A2(n_2575),
.B(n_2565),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2837),
.A2(n_2752),
.B1(n_2699),
.B2(n_2732),
.Y(n_3013)
);

NAND3xp33_ASAP7_75t_SL g3014 ( 
.A(n_2905),
.B(n_2798),
.C(n_2825),
.Y(n_3014)
);

BUFx12f_ASAP7_75t_L g3015 ( 
.A(n_2864),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_2790),
.Y(n_3016)
);

OAI21x1_ASAP7_75t_L g3017 ( 
.A1(n_2872),
.A2(n_2903),
.B(n_2816),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2865),
.A2(n_2684),
.B1(n_2732),
.B2(n_2733),
.Y(n_3018)
);

INVx1_ASAP7_75t_SL g3019 ( 
.A(n_2904),
.Y(n_3019)
);

BUFx3_ASAP7_75t_L g3020 ( 
.A(n_2790),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2889),
.A2(n_2656),
.B(n_2528),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2917),
.A2(n_2684),
.B1(n_2733),
.B2(n_2717),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2917),
.A2(n_2948),
.B1(n_2902),
.B2(n_2930),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2889),
.A2(n_2839),
.B(n_2843),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2970),
.Y(n_3025)
);

AOI222xp33_ASAP7_75t_L g3026 ( 
.A1(n_2965),
.A2(n_2677),
.B1(n_2702),
.B2(n_2679),
.C1(n_2634),
.C2(n_2676),
.Y(n_3026)
);

OR2x6_ASAP7_75t_L g3027 ( 
.A(n_2848),
.B(n_2549),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2784),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2970),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2822),
.B(n_2641),
.Y(n_3030)
);

OA21x2_ASAP7_75t_L g3031 ( 
.A1(n_2797),
.A2(n_2765),
.B(n_2763),
.Y(n_3031)
);

INVx6_ASAP7_75t_L g3032 ( 
.A(n_2779),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_2902),
.A2(n_2717),
.B1(n_2677),
.B2(n_2702),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2994),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2792),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2802),
.Y(n_3036)
);

AOI22xp5_ASAP7_75t_L g3037 ( 
.A1(n_3001),
.A2(n_2731),
.B1(n_2730),
.B2(n_2577),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2974),
.A2(n_2575),
.B1(n_2731),
.B2(n_2710),
.Y(n_3038)
);

INVx4_ASAP7_75t_L g3039 ( 
.A(n_2983),
.Y(n_3039)
);

AOI221xp5_ASAP7_75t_L g3040 ( 
.A1(n_2939),
.A2(n_2668),
.B1(n_2676),
.B2(n_2695),
.C(n_2691),
.Y(n_3040)
);

CKINVDCx11_ASAP7_75t_R g3041 ( 
.A(n_2866),
.Y(n_3041)
);

CKINVDCx5p33_ASAP7_75t_R g3042 ( 
.A(n_2864),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_SL g3043 ( 
.A1(n_2902),
.A2(n_2771),
.B1(n_2717),
.B2(n_2577),
.Y(n_3043)
);

INVx4_ASAP7_75t_L g3044 ( 
.A(n_2983),
.Y(n_3044)
);

AND2x4_ASAP7_75t_L g3045 ( 
.A(n_2861),
.B(n_2989),
.Y(n_3045)
);

OAI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2884),
.A2(n_2523),
.B1(n_2518),
.B2(n_2776),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_2930),
.A2(n_2652),
.B1(n_2641),
.B2(n_2716),
.Y(n_3047)
);

CKINVDCx20_ASAP7_75t_R g3048 ( 
.A(n_2922),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2815),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2988),
.B(n_2595),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2987),
.B(n_2523),
.Y(n_3051)
);

OAI211xp5_ASAP7_75t_L g3052 ( 
.A1(n_2916),
.A2(n_2595),
.B(n_2690),
.C(n_2724),
.Y(n_3052)
);

AOI22xp5_ASAP7_75t_SL g3053 ( 
.A1(n_2988),
.A2(n_2523),
.B1(n_2562),
.B2(n_2561),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_R g3054 ( 
.A(n_2971),
.B(n_2561),
.Y(n_3054)
);

OR2x6_ASAP7_75t_L g3055 ( 
.A(n_2848),
.B(n_2549),
.Y(n_3055)
);

INVx3_ASAP7_75t_L g3056 ( 
.A(n_2996),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2804),
.Y(n_3057)
);

OAI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2884),
.A2(n_2690),
.B1(n_2652),
.B2(n_2620),
.Y(n_3058)
);

OAI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_2795),
.A2(n_2982),
.B1(n_2807),
.B2(n_2853),
.Y(n_3059)
);

AOI221x1_ASAP7_75t_L g3060 ( 
.A1(n_2885),
.A2(n_2685),
.B1(n_2724),
.B2(n_2695),
.C(n_2691),
.Y(n_3060)
);

OAI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_2822),
.A2(n_2620),
.B1(n_2611),
.B2(n_2776),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_2971),
.Y(n_3062)
);

OAI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2997),
.A2(n_2755),
.B(n_2725),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2957),
.B(n_2611),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2942),
.B(n_2682),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2812),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_2996),
.Y(n_3067)
);

OAI21x1_ASAP7_75t_L g3068 ( 
.A1(n_2816),
.A2(n_2685),
.B(n_2706),
.Y(n_3068)
);

CKINVDCx11_ASAP7_75t_R g3069 ( 
.A(n_2815),
.Y(n_3069)
);

OAI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2929),
.A2(n_2823),
.B(n_2930),
.Y(n_3070)
);

OAI22xp5_ASAP7_75t_L g3071 ( 
.A1(n_2977),
.A2(n_2776),
.B1(n_2706),
.B2(n_2713),
.Y(n_3071)
);

OAI22xp5_ASAP7_75t_L g3072 ( 
.A1(n_2977),
.A2(n_2776),
.B1(n_2713),
.B2(n_2755),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2818),
.Y(n_3073)
);

OAI21x1_ASAP7_75t_L g3074 ( 
.A1(n_2796),
.A2(n_2725),
.B(n_2700),
.Y(n_3074)
);

OAI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2807),
.A2(n_2736),
.B1(n_2664),
.B2(n_2740),
.Y(n_3075)
);

INVx1_ASAP7_75t_SL g3076 ( 
.A(n_2911),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_2942),
.B(n_2688),
.Y(n_3077)
);

AOI221xp5_ASAP7_75t_L g3078 ( 
.A1(n_2939),
.A2(n_2562),
.B1(n_2724),
.B2(n_2673),
.C(n_2705),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2994),
.Y(n_3079)
);

AND2x4_ASAP7_75t_L g3080 ( 
.A(n_2848),
.B(n_2573),
.Y(n_3080)
);

AOI21xp33_ASAP7_75t_L g3081 ( 
.A1(n_2797),
.A2(n_2736),
.B(n_2738),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2957),
.B(n_2638),
.Y(n_3082)
);

NAND2x1p5_ASAP7_75t_L g3083 ( 
.A(n_2807),
.B(n_2664),
.Y(n_3083)
);

INVxp67_ASAP7_75t_L g3084 ( 
.A(n_2867),
.Y(n_3084)
);

BUFx6f_ASAP7_75t_L g3085 ( 
.A(n_2815),
.Y(n_3085)
);

BUFx5_ASAP7_75t_L g3086 ( 
.A(n_2928),
.Y(n_3086)
);

AOI22xp33_ASAP7_75t_L g3087 ( 
.A1(n_2931),
.A2(n_2645),
.B1(n_2573),
.B2(n_2748),
.Y(n_3087)
);

AO21x2_ASAP7_75t_L g3088 ( 
.A1(n_2951),
.A2(n_2748),
.B(n_2742),
.Y(n_3088)
);

OAI21xp33_ASAP7_75t_SL g3089 ( 
.A1(n_2993),
.A2(n_2775),
.B(n_2767),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2781),
.B(n_2638),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2928),
.A2(n_2664),
.B1(n_2562),
.B2(n_2767),
.Y(n_3091)
);

NOR3xp33_ASAP7_75t_L g3092 ( 
.A(n_2940),
.B(n_2962),
.C(n_2937),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_2796),
.A2(n_2952),
.B(n_2855),
.Y(n_3093)
);

OAI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2928),
.A2(n_2664),
.B1(n_2775),
.B2(n_2736),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2931),
.A2(n_2645),
.B1(n_2621),
.B2(n_2636),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_SL g3096 ( 
.A1(n_2807),
.A2(n_2638),
.B1(n_2698),
.B2(n_2550),
.Y(n_3096)
);

BUFx3_ASAP7_75t_L g3097 ( 
.A(n_2984),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2830),
.Y(n_3098)
);

HB1xp67_ASAP7_75t_L g3099 ( 
.A(n_2791),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2788),
.B(n_2964),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_2879),
.B(n_2638),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2835),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2789),
.B(n_2698),
.Y(n_3103)
);

INVx4_ASAP7_75t_L g3104 ( 
.A(n_2815),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2799),
.B(n_2698),
.Y(n_3105)
);

AOI221xp5_ASAP7_75t_L g3106 ( 
.A1(n_2929),
.A2(n_2743),
.B1(n_2740),
.B2(n_2742),
.C(n_2741),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2841),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2860),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2780),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2877),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2780),
.Y(n_3111)
);

INVx4_ASAP7_75t_L g3112 ( 
.A(n_2857),
.Y(n_3112)
);

OR2x2_ASAP7_75t_L g3113 ( 
.A(n_2908),
.B(n_2698),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2880),
.Y(n_3114)
);

NAND2xp33_ASAP7_75t_R g3115 ( 
.A(n_2984),
.B(n_2550),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_L g3116 ( 
.A1(n_2936),
.A2(n_2636),
.B1(n_2649),
.B2(n_2621),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_2791),
.Y(n_3117)
);

OR2x6_ASAP7_75t_L g3118 ( 
.A(n_2785),
.B(n_2621),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2794),
.Y(n_3119)
);

OAI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_2805),
.A2(n_2759),
.B(n_2741),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2794),
.Y(n_3121)
);

OAI21x1_ASAP7_75t_L g3122 ( 
.A1(n_2952),
.A2(n_2743),
.B(n_2721),
.Y(n_3122)
);

BUFx12f_ASAP7_75t_L g3123 ( 
.A(n_2978),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_SL g3124 ( 
.A1(n_3000),
.A2(n_2649),
.B1(n_2671),
.B2(n_2636),
.Y(n_3124)
);

OR2x2_ASAP7_75t_L g3125 ( 
.A(n_2908),
.B(n_2923),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2800),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2821),
.B(n_2721),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2891),
.Y(n_3128)
);

AOI221xp5_ASAP7_75t_L g3129 ( 
.A1(n_2936),
.A2(n_2759),
.B1(n_2672),
.B2(n_2681),
.C(n_2671),
.Y(n_3129)
);

AOI22xp33_ASAP7_75t_L g3130 ( 
.A1(n_2969),
.A2(n_2671),
.B1(n_2672),
.B2(n_2649),
.Y(n_3130)
);

BUFx12f_ASAP7_75t_L g3131 ( 
.A(n_2976),
.Y(n_3131)
);

OAI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_2920),
.A2(n_2721),
.B1(n_2681),
.B2(n_2672),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2782),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2783),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2924),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_2852),
.B(n_2681),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2859),
.B(n_2912),
.Y(n_3137)
);

INVx4_ASAP7_75t_L g3138 ( 
.A(n_2857),
.Y(n_3138)
);

OAI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_3000),
.A2(n_3003),
.B1(n_2920),
.B2(n_2886),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2935),
.Y(n_3140)
);

A2O1A1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_2901),
.A2(n_2721),
.B(n_2768),
.C(n_2764),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2800),
.Y(n_3142)
);

NOR3xp33_ASAP7_75t_SL g3143 ( 
.A(n_2899),
.B(n_32),
.C(n_33),
.Y(n_3143)
);

OAI22xp33_ASAP7_75t_L g3144 ( 
.A1(n_2968),
.A2(n_2764),
.B1(n_2768),
.B2(n_2701),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2941),
.Y(n_3145)
);

AOI22xp33_ASAP7_75t_L g3146 ( 
.A1(n_2969),
.A2(n_2701),
.B1(n_2768),
.B2(n_2764),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2793),
.B(n_34),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2867),
.B(n_34),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2831),
.Y(n_3149)
);

BUFx6f_ASAP7_75t_L g3150 ( 
.A(n_2857),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2840),
.B(n_2882),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_2851),
.A2(n_1219),
.B1(n_1234),
.B2(n_1215),
.Y(n_3152)
);

AND2x4_ASAP7_75t_L g3153 ( 
.A(n_2785),
.B(n_2915),
.Y(n_3153)
);

OR2x6_ASAP7_75t_L g3154 ( 
.A(n_2785),
.B(n_1215),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2966),
.Y(n_3155)
);

AOI21x1_ASAP7_75t_L g3156 ( 
.A1(n_2810),
.A2(n_35),
.B(n_37),
.Y(n_3156)
);

BUFx2_ASAP7_75t_L g3157 ( 
.A(n_2993),
.Y(n_3157)
);

HB1xp67_ASAP7_75t_L g3158 ( 
.A(n_2810),
.Y(n_3158)
);

AND2x4_ASAP7_75t_SL g3159 ( 
.A(n_3000),
.B(n_955),
.Y(n_3159)
);

AND2x4_ASAP7_75t_L g3160 ( 
.A(n_2915),
.B(n_37),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_3003),
.A2(n_1234),
.B1(n_1239),
.B2(n_1219),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_2829),
.B(n_38),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2890),
.A2(n_1427),
.B(n_1317),
.Y(n_3163)
);

BUFx2_ASAP7_75t_L g3164 ( 
.A(n_2992),
.Y(n_3164)
);

BUFx3_ASAP7_75t_L g3165 ( 
.A(n_2992),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_2934),
.B(n_38),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2973),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2985),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2975),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_R g3170 ( 
.A(n_2881),
.B(n_2985),
.Y(n_3170)
);

CKINVDCx11_ASAP7_75t_R g3171 ( 
.A(n_2857),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_3003),
.A2(n_1234),
.B1(n_1239),
.B2(n_1219),
.Y(n_3172)
);

CKINVDCx20_ASAP7_75t_R g3173 ( 
.A(n_2985),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2831),
.Y(n_3174)
);

AOI22xp5_ASAP7_75t_L g3175 ( 
.A1(n_2945),
.A2(n_1234),
.B1(n_1239),
.B2(n_1219),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2981),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2990),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2991),
.Y(n_3178)
);

AOI221xp5_ASAP7_75t_SL g3179 ( 
.A1(n_2979),
.A2(n_2910),
.B1(n_2944),
.B2(n_2938),
.C(n_2844),
.Y(n_3179)
);

AOI221xp5_ASAP7_75t_L g3180 ( 
.A1(n_2950),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.C(n_43),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_2787),
.B(n_43),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2820),
.Y(n_3182)
);

OAI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2819),
.A2(n_44),
.B(n_45),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2820),
.Y(n_3184)
);

BUFx2_ASAP7_75t_L g3185 ( 
.A(n_2859),
.Y(n_3185)
);

INVx6_ASAP7_75t_L g3186 ( 
.A(n_2926),
.Y(n_3186)
);

OAI21xp5_ASAP7_75t_SL g3187 ( 
.A1(n_2926),
.A2(n_46),
.B(n_47),
.Y(n_3187)
);

OR2x2_ASAP7_75t_L g3188 ( 
.A(n_2826),
.B(n_48),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2955),
.B(n_48),
.Y(n_3189)
);

OAI22xp5_ASAP7_75t_L g3190 ( 
.A1(n_2881),
.A2(n_53),
.B1(n_49),
.B2(n_50),
.Y(n_3190)
);

OR2x6_ASAP7_75t_L g3191 ( 
.A(n_2849),
.B(n_1219),
.Y(n_3191)
);

AOI221xp5_ASAP7_75t_L g3192 ( 
.A1(n_2950),
.A2(n_53),
.B1(n_49),
.B2(n_50),
.C(n_54),
.Y(n_3192)
);

NAND2x1p5_ASAP7_75t_L g3193 ( 
.A(n_2912),
.B(n_1317),
.Y(n_3193)
);

CKINVDCx11_ASAP7_75t_R g3194 ( 
.A(n_2926),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2955),
.B(n_54),
.Y(n_3195)
);

INVx1_ASAP7_75t_SL g3196 ( 
.A(n_2881),
.Y(n_3196)
);

HB1xp67_ASAP7_75t_L g3197 ( 
.A(n_2871),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2949),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_2960),
.A2(n_2961),
.B1(n_2956),
.B2(n_2963),
.Y(n_3199)
);

AOI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_2956),
.A2(n_1239),
.B1(n_1259),
.B2(n_1234),
.Y(n_3200)
);

OAI22xp5_ASAP7_75t_L g3201 ( 
.A1(n_2850),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_L g3202 ( 
.A(n_2959),
.B(n_2943),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3182),
.Y(n_3203)
);

INVxp67_ASAP7_75t_L g3204 ( 
.A(n_3065),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3184),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3099),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_3117),
.Y(n_3207)
);

BUFx2_ASAP7_75t_L g3208 ( 
.A(n_3170),
.Y(n_3208)
);

BUFx10_ASAP7_75t_L g3209 ( 
.A(n_3160),
.Y(n_3209)
);

INVx2_ASAP7_75t_SL g3210 ( 
.A(n_3032),
.Y(n_3210)
);

BUFx2_ASAP7_75t_L g3211 ( 
.A(n_3197),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3031),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_3093),
.Y(n_3213)
);

HB1xp67_ASAP7_75t_L g3214 ( 
.A(n_3158),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_3031),
.Y(n_3215)
);

OAI21x1_ASAP7_75t_L g3216 ( 
.A1(n_3017),
.A2(n_2786),
.B(n_2806),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_3041),
.Y(n_3217)
);

NOR2x1_ASAP7_75t_R g3218 ( 
.A(n_3039),
.B(n_2943),
.Y(n_3218)
);

OR2x6_ASAP7_75t_L g3219 ( 
.A(n_3027),
.B(n_2873),
.Y(n_3219)
);

INVx2_ASAP7_75t_SL g3220 ( 
.A(n_3032),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_3025),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3135),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3140),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3145),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3155),
.Y(n_3225)
);

HB1xp67_ASAP7_75t_L g3226 ( 
.A(n_3030),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_3153),
.B(n_2869),
.Y(n_3227)
);

BUFx2_ASAP7_75t_L g3228 ( 
.A(n_3045),
.Y(n_3228)
);

HB1xp67_ASAP7_75t_L g3229 ( 
.A(n_3030),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3029),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3034),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_3079),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3109),
.Y(n_3233)
);

BUFx2_ASAP7_75t_L g3234 ( 
.A(n_3045),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3167),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_3012),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3111),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3119),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3169),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_3151),
.B(n_2871),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3176),
.Y(n_3241)
);

HB1xp67_ASAP7_75t_L g3242 ( 
.A(n_3195),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3019),
.B(n_2906),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3177),
.Y(n_3244)
);

INVx3_ASAP7_75t_L g3245 ( 
.A(n_3086),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_3100),
.B(n_2906),
.Y(n_3246)
);

BUFx6f_ASAP7_75t_L g3247 ( 
.A(n_3160),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_3153),
.B(n_2869),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3121),
.Y(n_3249)
);

OR2x6_ASAP7_75t_L g3250 ( 
.A(n_3027),
.B(n_2806),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3084),
.B(n_2946),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3068),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3178),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3028),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_3126),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3142),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3149),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3035),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3174),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3036),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_3086),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3133),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3198),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3057),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_3086),
.Y(n_3265)
);

BUFx2_ASAP7_75t_L g3266 ( 
.A(n_3007),
.Y(n_3266)
);

OR2x2_ASAP7_75t_L g3267 ( 
.A(n_3125),
.B(n_3019),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3066),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3073),
.Y(n_3269)
);

OR2x2_ASAP7_75t_L g3270 ( 
.A(n_3113),
.B(n_2946),
.Y(n_3270)
);

BUFx2_ASAP7_75t_L g3271 ( 
.A(n_3173),
.Y(n_3271)
);

AO21x2_ASAP7_75t_L g3272 ( 
.A1(n_3070),
.A2(n_2951),
.B(n_2898),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3077),
.B(n_3076),
.Y(n_3273)
);

BUFx6f_ASAP7_75t_L g3274 ( 
.A(n_3015),
.Y(n_3274)
);

OAI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_3014),
.A2(n_2850),
.B(n_2887),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_3195),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3098),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3102),
.Y(n_3278)
);

AO21x2_ASAP7_75t_L g3279 ( 
.A1(n_3070),
.A2(n_3183),
.B(n_3004),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_3076),
.B(n_2995),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3107),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3108),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3110),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3114),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3128),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_3136),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_3042),
.B(n_2947),
.Y(n_3287)
);

OA21x2_ASAP7_75t_L g3288 ( 
.A1(n_3024),
.A2(n_2786),
.B(n_2845),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3134),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_3080),
.B(n_2995),
.Y(n_3290)
);

AO21x2_ASAP7_75t_L g3291 ( 
.A1(n_3183),
.A2(n_2846),
.B(n_2868),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3189),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3188),
.B(n_2900),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3105),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3092),
.B(n_2972),
.Y(n_3295)
);

AND2x4_ASAP7_75t_L g3296 ( 
.A(n_3080),
.B(n_2915),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3064),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3090),
.Y(n_3298)
);

CKINVDCx20_ASAP7_75t_R g3299 ( 
.A(n_3048),
.Y(n_3299)
);

BUFx2_ASAP7_75t_L g3300 ( 
.A(n_3157),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_3049),
.Y(n_3301)
);

AO21x1_ASAP7_75t_SL g3302 ( 
.A1(n_3120),
.A2(n_2932),
.B(n_2813),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3196),
.B(n_3127),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3101),
.Y(n_3304)
);

NOR2xp33_ASAP7_75t_L g3305 ( 
.A(n_3016),
.B(n_2947),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3051),
.B(n_2827),
.Y(n_3306)
);

INVx4_ASAP7_75t_L g3307 ( 
.A(n_3039),
.Y(n_3307)
);

OA21x2_ASAP7_75t_L g3308 ( 
.A1(n_3011),
.A2(n_2856),
.B(n_2845),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3082),
.Y(n_3309)
);

AO21x2_ASAP7_75t_L g3310 ( 
.A1(n_3004),
.A2(n_2846),
.B(n_2868),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3101),
.Y(n_3311)
);

OR2x2_ASAP7_75t_L g3312 ( 
.A(n_3164),
.B(n_2827),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3185),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3009),
.Y(n_3314)
);

AO21x2_ASAP7_75t_L g3315 ( 
.A1(n_3059),
.A2(n_3008),
.B(n_3201),
.Y(n_3315)
);

OAI21x1_ASAP7_75t_L g3316 ( 
.A1(n_3122),
.A2(n_2856),
.B(n_2833),
.Y(n_3316)
);

BUFx4f_ASAP7_75t_L g3317 ( 
.A(n_3193),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3086),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3009),
.B(n_2827),
.Y(n_3319)
);

AND2x2_ASAP7_75t_L g3320 ( 
.A(n_3103),
.B(n_2972),
.Y(n_3320)
);

INVx3_ASAP7_75t_L g3321 ( 
.A(n_3086),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3154),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3154),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3154),
.Y(n_3324)
);

OAI21x1_ASAP7_75t_L g3325 ( 
.A1(n_3071),
.A2(n_2933),
.B(n_2894),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3118),
.Y(n_3326)
);

OA21x2_ASAP7_75t_L g3327 ( 
.A1(n_3060),
.A2(n_2933),
.B(n_2838),
.Y(n_3327)
);

HB1xp67_ASAP7_75t_L g3328 ( 
.A(n_3196),
.Y(n_3328)
);

OAI21x1_ASAP7_75t_L g3329 ( 
.A1(n_3071),
.A2(n_2838),
.B(n_2874),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3165),
.B(n_2972),
.Y(n_3330)
);

INVx3_ASAP7_75t_L g3331 ( 
.A(n_3104),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3074),
.Y(n_3332)
);

BUFx2_ASAP7_75t_L g3333 ( 
.A(n_3056),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3156),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3118),
.Y(n_3335)
);

INVx3_ASAP7_75t_L g3336 ( 
.A(n_3104),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3118),
.Y(n_3337)
);

INVx4_ASAP7_75t_L g3338 ( 
.A(n_3044),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3027),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3061),
.Y(n_3340)
);

BUFx2_ASAP7_75t_L g3341 ( 
.A(n_3056),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3061),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3055),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3062),
.B(n_2958),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3067),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3067),
.B(n_3168),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3191),
.B(n_3147),
.Y(n_3347)
);

OR2x2_ASAP7_75t_SL g3348 ( 
.A(n_3148),
.B(n_2926),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3055),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3055),
.Y(n_3350)
);

HB1xp67_ASAP7_75t_L g3351 ( 
.A(n_3139),
.Y(n_3351)
);

INVxp67_ASAP7_75t_SL g3352 ( 
.A(n_3139),
.Y(n_3352)
);

INVxp67_ASAP7_75t_SL g3353 ( 
.A(n_3115),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3088),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3191),
.Y(n_3355)
);

AND2x4_ASAP7_75t_L g3356 ( 
.A(n_3053),
.B(n_2958),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3191),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3088),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3186),
.Y(n_3359)
);

OA21x2_ASAP7_75t_L g3360 ( 
.A1(n_3063),
.A2(n_3002),
.B(n_2954),
.Y(n_3360)
);

OA21x2_ASAP7_75t_L g3361 ( 
.A1(n_3063),
.A2(n_3002),
.B(n_2954),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3097),
.B(n_2972),
.Y(n_3362)
);

OAI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3038),
.A2(n_2832),
.B(n_2925),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3131),
.B(n_2953),
.Y(n_3364)
);

INVx2_ASAP7_75t_SL g3365 ( 
.A(n_3186),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3179),
.B(n_2953),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_SL g3367 ( 
.A1(n_3279),
.A2(n_3038),
.B1(n_3201),
.B2(n_3013),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3222),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3352),
.A2(n_3023),
.B1(n_3187),
.B2(n_3058),
.Y(n_3369)
);

AOI221x1_ASAP7_75t_SL g3370 ( 
.A1(n_3292),
.A2(n_3166),
.B1(n_3181),
.B2(n_3190),
.C(n_3058),
.Y(n_3370)
);

OAI221xp5_ASAP7_75t_L g3371 ( 
.A1(n_3275),
.A2(n_3179),
.B1(n_3143),
.B2(n_3043),
.C(n_3187),
.Y(n_3371)
);

AOI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3279),
.A2(n_3046),
.B(n_3137),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3279),
.A2(n_3315),
.B(n_3353),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3242),
.B(n_3276),
.Y(n_3374)
);

OAI21x1_ASAP7_75t_L g3375 ( 
.A1(n_3236),
.A2(n_3213),
.B(n_3331),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3351),
.A2(n_3037),
.B1(n_3124),
.B2(n_3005),
.Y(n_3376)
);

OA21x2_ASAP7_75t_L g3377 ( 
.A1(n_3212),
.A2(n_3047),
.B(n_3120),
.Y(n_3377)
);

INVx3_ASAP7_75t_L g3378 ( 
.A(n_3356),
.Y(n_3378)
);

AOI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_3315),
.A2(n_3006),
.B(n_3091),
.Y(n_3379)
);

OA21x2_ASAP7_75t_L g3380 ( 
.A1(n_3212),
.A2(n_3081),
.B(n_3033),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_SL g3381 ( 
.A1(n_3315),
.A2(n_3013),
.B1(n_3072),
.B2(n_3123),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3268),
.Y(n_3382)
);

AOI222xp33_ASAP7_75t_L g3383 ( 
.A1(n_3292),
.A2(n_3180),
.B1(n_3192),
.B2(n_3072),
.C1(n_3010),
.C2(n_3190),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3228),
.B(n_3202),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3222),
.Y(n_3385)
);

INVx2_ASAP7_75t_SL g3386 ( 
.A(n_3271),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3223),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3228),
.B(n_3050),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3268),
.Y(n_3389)
);

BUFx3_ASAP7_75t_L g3390 ( 
.A(n_3299),
.Y(n_3390)
);

BUFx3_ASAP7_75t_L g3391 ( 
.A(n_3217),
.Y(n_3391)
);

OAI221xp5_ASAP7_75t_L g3392 ( 
.A1(n_3366),
.A2(n_3052),
.B1(n_3095),
.B2(n_3026),
.C(n_3022),
.Y(n_3392)
);

OA21x2_ASAP7_75t_L g3393 ( 
.A1(n_3215),
.A2(n_3081),
.B(n_3021),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_SL g3394 ( 
.A1(n_3310),
.A2(n_3091),
.B1(n_3094),
.B2(n_3162),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3223),
.Y(n_3395)
);

OAI21x1_ASAP7_75t_L g3396 ( 
.A1(n_3236),
.A2(n_3083),
.B(n_3094),
.Y(n_3396)
);

AOI221xp5_ASAP7_75t_L g3397 ( 
.A1(n_3334),
.A2(n_3040),
.B1(n_3087),
.B2(n_3078),
.C(n_3018),
.Y(n_3397)
);

OAI221xp5_ASAP7_75t_L g3398 ( 
.A1(n_3334),
.A2(n_3026),
.B1(n_3141),
.B2(n_3116),
.C(n_3129),
.Y(n_3398)
);

OAI22xp5_ASAP7_75t_SL g3399 ( 
.A1(n_3208),
.A2(n_3044),
.B1(n_3020),
.B2(n_3054),
.Y(n_3399)
);

AOI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3310),
.A2(n_3159),
.B1(n_3144),
.B2(n_3146),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3234),
.B(n_3069),
.Y(n_3401)
);

AO31x2_ASAP7_75t_L g3402 ( 
.A1(n_3354),
.A2(n_2921),
.A3(n_2875),
.B(n_2878),
.Y(n_3402)
);

AOI221xp5_ASAP7_75t_SL g3403 ( 
.A1(n_3295),
.A2(n_3089),
.B1(n_3132),
.B2(n_3106),
.C(n_3152),
.Y(n_3403)
);

NAND3xp33_ASAP7_75t_L g3404 ( 
.A(n_3340),
.B(n_3175),
.C(n_3130),
.Y(n_3404)
);

OR2x2_ASAP7_75t_L g3405 ( 
.A(n_3246),
.B(n_3112),
.Y(n_3405)
);

AOI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3310),
.A2(n_3199),
.B1(n_2801),
.B2(n_3172),
.Y(n_3406)
);

AOI221xp5_ASAP7_75t_L g3407 ( 
.A1(n_3291),
.A2(n_3363),
.B1(n_3229),
.B2(n_3226),
.C(n_3332),
.Y(n_3407)
);

AND2x4_ASAP7_75t_L g3408 ( 
.A(n_3208),
.B(n_3112),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3234),
.B(n_3273),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3273),
.B(n_3171),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_3274),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3224),
.Y(n_3412)
);

OR2x2_ASAP7_75t_SL g3413 ( 
.A(n_3247),
.B(n_2953),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_3356),
.Y(n_3414)
);

OR2x2_ASAP7_75t_L g3415 ( 
.A(n_3246),
.B(n_3138),
.Y(n_3415)
);

AOI22xp33_ASAP7_75t_L g3416 ( 
.A1(n_3291),
.A2(n_3161),
.B1(n_2876),
.B2(n_2828),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_L g3417 ( 
.A1(n_3291),
.A2(n_2876),
.B1(n_2828),
.B2(n_3096),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3224),
.Y(n_3418)
);

OAI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_3348),
.A2(n_3138),
.B1(n_2953),
.B2(n_3085),
.Y(n_3419)
);

OAI221xp5_ASAP7_75t_L g3420 ( 
.A1(n_3349),
.A2(n_3219),
.B1(n_3250),
.B2(n_3293),
.C(n_3339),
.Y(n_3420)
);

OAI211xp5_ASAP7_75t_L g3421 ( 
.A1(n_3266),
.A2(n_3194),
.B(n_3049),
.C(n_3150),
.Y(n_3421)
);

AOI22xp33_ASAP7_75t_L g3422 ( 
.A1(n_3219),
.A2(n_2828),
.B1(n_2897),
.B2(n_3075),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3225),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3225),
.Y(n_3424)
);

OR2x2_ASAP7_75t_L g3425 ( 
.A(n_3267),
.B(n_3049),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3235),
.Y(n_3426)
);

INVx4_ASAP7_75t_L g3427 ( 
.A(n_3274),
.Y(n_3427)
);

CKINVDCx5p33_ASAP7_75t_R g3428 ( 
.A(n_3274),
.Y(n_3428)
);

OAI22xp5_ASAP7_75t_SL g3429 ( 
.A1(n_3266),
.A2(n_3083),
.B1(n_3150),
.B2(n_3085),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3235),
.Y(n_3430)
);

AOI22xp5_ASAP7_75t_SL g3431 ( 
.A1(n_3271),
.A2(n_3150),
.B1(n_3085),
.B2(n_3193),
.Y(n_3431)
);

OAI221xp5_ASAP7_75t_L g3432 ( 
.A1(n_3349),
.A2(n_3163),
.B1(n_2878),
.B2(n_2893),
.C(n_2875),
.Y(n_3432)
);

NAND3xp33_ASAP7_75t_L g3433 ( 
.A(n_3340),
.B(n_2778),
.C(n_3200),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3283),
.Y(n_3434)
);

OAI22xp5_ASAP7_75t_L g3435 ( 
.A1(n_3348),
.A2(n_2858),
.B1(n_2863),
.B2(n_2980),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3267),
.A2(n_2980),
.B1(n_2778),
.B2(n_2986),
.Y(n_3436)
);

AOI221xp5_ASAP7_75t_L g3437 ( 
.A1(n_3332),
.A2(n_2895),
.B1(n_2913),
.B2(n_2893),
.C(n_2834),
.Y(n_3437)
);

NOR2x1_ASAP7_75t_SL g3438 ( 
.A(n_3302),
.B(n_2897),
.Y(n_3438)
);

OAI22xp5_ASAP7_75t_L g3439 ( 
.A1(n_3204),
.A2(n_2778),
.B1(n_2895),
.B2(n_2834),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3227),
.B(n_2909),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3283),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3239),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3219),
.A2(n_2919),
.B1(n_2927),
.B2(n_2913),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_L g3444 ( 
.A1(n_3219),
.A2(n_3347),
.B1(n_3247),
.B2(n_3302),
.Y(n_3444)
);

OAI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3219),
.A2(n_2927),
.B1(n_2919),
.B2(n_2998),
.Y(n_3445)
);

NAND3xp33_ASAP7_75t_L g3446 ( 
.A(n_3342),
.B(n_2998),
.C(n_960),
.Y(n_3446)
);

INVxp67_ASAP7_75t_SL g3447 ( 
.A(n_3252),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3239),
.Y(n_3448)
);

OAI21x1_ASAP7_75t_L g3449 ( 
.A1(n_3236),
.A2(n_2836),
.B(n_2824),
.Y(n_3449)
);

HB1xp67_ASAP7_75t_L g3450 ( 
.A(n_3211),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3289),
.Y(n_3451)
);

NAND3xp33_ASAP7_75t_L g3452 ( 
.A(n_3342),
.B(n_2998),
.C(n_960),
.Y(n_3452)
);

AO21x2_ASAP7_75t_L g3453 ( 
.A1(n_3252),
.A2(n_2914),
.B(n_2918),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3347),
.A2(n_2888),
.B1(n_2907),
.B2(n_2808),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_3247),
.A2(n_2862),
.B1(n_2870),
.B2(n_2892),
.Y(n_3455)
);

BUFx12f_ASAP7_75t_L g3456 ( 
.A(n_3274),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_SL g3457 ( 
.A1(n_3209),
.A2(n_2854),
.B1(n_2883),
.B2(n_2842),
.Y(n_3457)
);

OAI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3251),
.A2(n_2842),
.B(n_55),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_3247),
.A2(n_3272),
.B1(n_3298),
.B2(n_3294),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3241),
.Y(n_3460)
);

AOI22xp33_ASAP7_75t_L g3461 ( 
.A1(n_3247),
.A2(n_1259),
.B1(n_1277),
.B2(n_1239),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3272),
.A2(n_1277),
.B1(n_1259),
.B2(n_60),
.Y(n_3462)
);

OR2x2_ASAP7_75t_L g3463 ( 
.A(n_3207),
.B(n_2967),
.Y(n_3463)
);

OA21x2_ASAP7_75t_L g3464 ( 
.A1(n_3215),
.A2(n_2967),
.B(n_58),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_3272),
.A2(n_1277),
.B1(n_1259),
.B2(n_61),
.Y(n_3465)
);

OAI221xp5_ASAP7_75t_L g3466 ( 
.A1(n_3250),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.C(n_64),
.Y(n_3466)
);

OAI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3243),
.A2(n_59),
.B(n_62),
.Y(n_3467)
);

OAI211xp5_ASAP7_75t_L g3468 ( 
.A1(n_3300),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_3468)
);

INVx1_ASAP7_75t_SL g3469 ( 
.A(n_3364),
.Y(n_3469)
);

AO21x2_ASAP7_75t_L g3470 ( 
.A1(n_3252),
.A2(n_2967),
.B(n_65),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_L g3471 ( 
.A1(n_3294),
.A2(n_1277),
.B1(n_1259),
.B2(n_71),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3289),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3286),
.Y(n_3473)
);

BUFx2_ASAP7_75t_L g3474 ( 
.A(n_3300),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3298),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_3475)
);

AOI21xp33_ASAP7_75t_L g3476 ( 
.A1(n_3322),
.A2(n_72),
.B(n_73),
.Y(n_3476)
);

AOI22xp33_ASAP7_75t_L g3477 ( 
.A1(n_3209),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_3210),
.B(n_75),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_SL g3479 ( 
.A1(n_3209),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3297),
.B(n_2967),
.Y(n_3480)
);

AND2x2_ASAP7_75t_L g3481 ( 
.A(n_3227),
.B(n_78),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3209),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3241),
.Y(n_3483)
);

BUFx2_ASAP7_75t_L g3484 ( 
.A(n_3280),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3227),
.B(n_79),
.Y(n_3485)
);

OAI221xp5_ASAP7_75t_L g3486 ( 
.A1(n_3250),
.A2(n_84),
.B1(n_80),
.B2(n_83),
.C(n_85),
.Y(n_3486)
);

AOI221xp5_ASAP7_75t_L g3487 ( 
.A1(n_3297),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.C(n_87),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3286),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_3488)
);

AOI221xp5_ASAP7_75t_L g3489 ( 
.A1(n_3306),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.C(n_94),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3262),
.Y(n_3490)
);

OAI211xp5_ASAP7_75t_L g3491 ( 
.A1(n_3307),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_3491)
);

AND2x4_ASAP7_75t_L g3492 ( 
.A(n_3210),
.B(n_3220),
.Y(n_3492)
);

OAI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3317),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3493)
);

OAI221xp5_ASAP7_75t_L g3494 ( 
.A1(n_3250),
.A2(n_3350),
.B1(n_3343),
.B2(n_3339),
.C(n_3323),
.Y(n_3494)
);

AOI221xp5_ASAP7_75t_L g3495 ( 
.A1(n_3306),
.A2(n_100),
.B1(n_96),
.B2(n_98),
.C(n_101),
.Y(n_3495)
);

OAI211xp5_ASAP7_75t_L g3496 ( 
.A1(n_3307),
.A2(n_102),
.B(n_98),
.C(n_101),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3220),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_3497)
);

AOI221xp5_ASAP7_75t_L g3498 ( 
.A1(n_3263),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.C(n_107),
.Y(n_3498)
);

AOI22x1_ASAP7_75t_L g3499 ( 
.A1(n_3307),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_3499)
);

INVxp67_ASAP7_75t_SL g3500 ( 
.A(n_3373),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3374),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3444),
.B(n_3243),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3444),
.B(n_3314),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3370),
.B(n_3367),
.Y(n_3504)
);

AOI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3367),
.A2(n_3350),
.B1(n_3343),
.B2(n_3337),
.Y(n_3505)
);

BUFx2_ASAP7_75t_L g3506 ( 
.A(n_3411),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3378),
.B(n_3314),
.Y(n_3507)
);

BUFx2_ASAP7_75t_L g3508 ( 
.A(n_3411),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3368),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_3456),
.B(n_3274),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3403),
.B(n_3211),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3378),
.B(n_3414),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3385),
.Y(n_3513)
);

OAI221xp5_ASAP7_75t_L g3514 ( 
.A1(n_3381),
.A2(n_3250),
.B1(n_3312),
.B2(n_3319),
.C(n_3322),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3387),
.B(n_3214),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3414),
.B(n_3333),
.Y(n_3516)
);

OR2x6_ASAP7_75t_SL g3517 ( 
.A(n_3428),
.B(n_3313),
.Y(n_3517)
);

OR2x2_ASAP7_75t_L g3518 ( 
.A(n_3395),
.B(n_3206),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3409),
.B(n_3333),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3383),
.B(n_3206),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_3390),
.Y(n_3521)
);

OR2x2_ASAP7_75t_L g3522 ( 
.A(n_3412),
.B(n_3203),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3490),
.Y(n_3523)
);

BUFx8_ASAP7_75t_SL g3524 ( 
.A(n_3391),
.Y(n_3524)
);

HB1xp67_ASAP7_75t_L g3525 ( 
.A(n_3450),
.Y(n_3525)
);

BUFx3_ASAP7_75t_L g3526 ( 
.A(n_3427),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3418),
.Y(n_3527)
);

OR2x2_ASAP7_75t_L g3528 ( 
.A(n_3423),
.B(n_3203),
.Y(n_3528)
);

OR2x2_ASAP7_75t_L g3529 ( 
.A(n_3424),
.B(n_3205),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3426),
.Y(n_3530)
);

AND2x4_ASAP7_75t_L g3531 ( 
.A(n_3408),
.B(n_3356),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3484),
.B(n_3341),
.Y(n_3532)
);

INVxp67_ASAP7_75t_SL g3533 ( 
.A(n_3438),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_3430),
.B(n_3205),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3408),
.B(n_3341),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3369),
.B(n_3244),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3382),
.Y(n_3537)
);

INVx1_ASAP7_75t_SL g3538 ( 
.A(n_3384),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3401),
.B(n_3319),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3492),
.B(n_3346),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_3389),
.Y(n_3541)
);

BUFx2_ASAP7_75t_L g3542 ( 
.A(n_3427),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3442),
.B(n_3262),
.Y(n_3543)
);

AND2x4_ASAP7_75t_SL g3544 ( 
.A(n_3388),
.B(n_3307),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3492),
.B(n_3346),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3450),
.B(n_3244),
.Y(n_3546)
);

INVx3_ASAP7_75t_L g3547 ( 
.A(n_3375),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3448),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3474),
.B(n_3253),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3460),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3483),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3434),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3386),
.B(n_3253),
.Y(n_3553)
);

AND2x2_ASAP7_75t_L g3554 ( 
.A(n_3469),
.B(n_3290),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3396),
.Y(n_3555)
);

NOR2x1_ASAP7_75t_L g3556 ( 
.A(n_3481),
.B(n_3338),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3410),
.B(n_3290),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3431),
.B(n_3290),
.Y(n_3558)
);

INVx3_ASAP7_75t_L g3559 ( 
.A(n_3393),
.Y(n_3559)
);

OAI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_3381),
.A2(n_3338),
.B1(n_3356),
.B2(n_3261),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3440),
.B(n_3290),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3407),
.B(n_3254),
.Y(n_3562)
);

NAND3xp33_ASAP7_75t_L g3563 ( 
.A(n_3433),
.B(n_3357),
.C(n_3355),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3441),
.Y(n_3564)
);

OR2x2_ASAP7_75t_L g3565 ( 
.A(n_3451),
.B(n_3262),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3405),
.B(n_3280),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3472),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3415),
.B(n_3227),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3464),
.Y(n_3569)
);

BUFx2_ASAP7_75t_L g3570 ( 
.A(n_3413),
.Y(n_3570)
);

INVx3_ASAP7_75t_L g3571 ( 
.A(n_3393),
.Y(n_3571)
);

OR2x2_ASAP7_75t_L g3572 ( 
.A(n_3376),
.B(n_3263),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3404),
.Y(n_3573)
);

INVxp67_ASAP7_75t_SL g3574 ( 
.A(n_3379),
.Y(n_3574)
);

HB1xp67_ASAP7_75t_L g3575 ( 
.A(n_3425),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3394),
.B(n_3248),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3464),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3464),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3447),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3485),
.B(n_3254),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3394),
.B(n_3248),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3447),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3377),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3377),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3372),
.B(n_3248),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3473),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3371),
.A2(n_3406),
.B1(n_3458),
.B2(n_3466),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3421),
.B(n_3248),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3377),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3399),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3393),
.B(n_3240),
.Y(n_3591)
);

BUFx2_ASAP7_75t_L g3592 ( 
.A(n_3429),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3397),
.B(n_3258),
.Y(n_3593)
);

INVx2_ASAP7_75t_SL g3594 ( 
.A(n_3463),
.Y(n_3594)
);

NOR2x1_ASAP7_75t_L g3595 ( 
.A(n_3478),
.B(n_3338),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3419),
.B(n_3240),
.Y(n_3596)
);

AOI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3392),
.A2(n_3337),
.B1(n_3326),
.B2(n_3324),
.Y(n_3597)
);

HB1xp67_ASAP7_75t_L g3598 ( 
.A(n_3439),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3480),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3478),
.B(n_3258),
.Y(n_3600)
);

BUFx2_ASAP7_75t_L g3601 ( 
.A(n_3467),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3380),
.Y(n_3602)
);

INVx3_ASAP7_75t_L g3603 ( 
.A(n_3449),
.Y(n_3603)
);

INVx2_ASAP7_75t_SL g3604 ( 
.A(n_3380),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3470),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3457),
.B(n_3328),
.Y(n_3606)
);

HB1xp67_ASAP7_75t_L g3607 ( 
.A(n_3486),
.Y(n_3607)
);

AND2x4_ASAP7_75t_L g3608 ( 
.A(n_3422),
.B(n_3338),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3470),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3406),
.B(n_3260),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3453),
.Y(n_3611)
);

INVxp67_ASAP7_75t_SL g3612 ( 
.A(n_3454),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3398),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3462),
.B(n_3260),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_3453),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3494),
.Y(n_3616)
);

OR2x2_ASAP7_75t_L g3617 ( 
.A(n_3436),
.B(n_3264),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3457),
.B(n_3313),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3455),
.B(n_3365),
.Y(n_3619)
);

NOR2xp67_ASAP7_75t_L g3620 ( 
.A(n_3420),
.B(n_3245),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3400),
.Y(n_3621)
);

OR2x2_ASAP7_75t_L g3622 ( 
.A(n_3459),
.B(n_3264),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3432),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3459),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3455),
.B(n_3365),
.Y(n_3625)
);

OAI22xp5_ASAP7_75t_L g3626 ( 
.A1(n_3462),
.A2(n_3261),
.B1(n_3265),
.B2(n_3245),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_L g3627 ( 
.A(n_3524),
.B(n_3287),
.Y(n_3627)
);

OAI22xp5_ASAP7_75t_L g3628 ( 
.A1(n_3574),
.A2(n_3422),
.B1(n_3465),
.B2(n_3479),
.Y(n_3628)
);

OR2x2_ASAP7_75t_L g3629 ( 
.A(n_3520),
.B(n_3270),
.Y(n_3629)
);

OR2x2_ASAP7_75t_L g3630 ( 
.A(n_3538),
.B(n_3270),
.Y(n_3630)
);

OAI22xp33_ASAP7_75t_L g3631 ( 
.A1(n_3514),
.A2(n_3435),
.B1(n_3445),
.B2(n_3312),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3613),
.A2(n_3416),
.B1(n_3465),
.B2(n_3417),
.Y(n_3632)
);

AOI222xp33_ASAP7_75t_L g3633 ( 
.A1(n_3504),
.A2(n_3495),
.B1(n_3489),
.B2(n_3487),
.C1(n_3416),
.C2(n_3498),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3509),
.Y(n_3634)
);

AOI222xp33_ASAP7_75t_L g3635 ( 
.A1(n_3587),
.A2(n_3468),
.B1(n_3417),
.B2(n_3488),
.C1(n_3497),
.C2(n_3437),
.Y(n_3635)
);

NAND2xp33_ASAP7_75t_R g3636 ( 
.A(n_3601),
.B(n_3296),
.Y(n_3636)
);

OAI211xp5_ASAP7_75t_L g3637 ( 
.A1(n_3590),
.A2(n_3479),
.B(n_3496),
.C(n_3491),
.Y(n_3637)
);

BUFx3_ASAP7_75t_L g3638 ( 
.A(n_3524),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_3575),
.Y(n_3639)
);

AOI22xp33_ASAP7_75t_SL g3640 ( 
.A1(n_3500),
.A2(n_3499),
.B1(n_3288),
.B2(n_3213),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3512),
.Y(n_3641)
);

AND4x1_ASAP7_75t_L g3642 ( 
.A(n_3595),
.B(n_3477),
.C(n_3482),
.D(n_3488),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3601),
.B(n_3269),
.Y(n_3643)
);

OAI21x1_ASAP7_75t_L g3644 ( 
.A1(n_3555),
.A2(n_3236),
.B(n_3213),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3557),
.B(n_3362),
.Y(n_3645)
);

OAI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3560),
.A2(n_3511),
.B(n_3593),
.Y(n_3646)
);

AOI22xp33_ASAP7_75t_L g3647 ( 
.A1(n_3624),
.A2(n_3443),
.B1(n_3288),
.B2(n_3335),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3512),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3569),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3569),
.Y(n_3650)
);

OAI221xp5_ASAP7_75t_L g3651 ( 
.A1(n_3607),
.A2(n_3477),
.B1(n_3482),
.B2(n_3475),
.C(n_3476),
.Y(n_3651)
);

BUFx6f_ASAP7_75t_L g3652 ( 
.A(n_3526),
.Y(n_3652)
);

AND2x2_ASAP7_75t_SL g3653 ( 
.A(n_3592),
.B(n_3317),
.Y(n_3653)
);

AO21x2_ASAP7_75t_L g3654 ( 
.A1(n_3602),
.A2(n_3493),
.B(n_3358),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3577),
.Y(n_3655)
);

OAI211xp5_ASAP7_75t_L g3656 ( 
.A1(n_3590),
.A2(n_3475),
.B(n_3213),
.C(n_3288),
.Y(n_3656)
);

NAND2xp33_ASAP7_75t_SL g3657 ( 
.A(n_3540),
.B(n_3364),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3513),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3527),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3577),
.Y(n_3660)
);

NAND4xp25_ASAP7_75t_L g3661 ( 
.A(n_3618),
.B(n_3305),
.C(n_3344),
.D(n_3345),
.Y(n_3661)
);

NAND4xp25_ASAP7_75t_L g3662 ( 
.A(n_3618),
.B(n_3345),
.C(n_3362),
.D(n_3336),
.Y(n_3662)
);

OAI31xp33_ASAP7_75t_L g3663 ( 
.A1(n_3563),
.A2(n_3493),
.A3(n_3443),
.B(n_3452),
.Y(n_3663)
);

OAI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_3592),
.A2(n_3261),
.B1(n_3265),
.B2(n_3245),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3621),
.A2(n_3288),
.B1(n_3335),
.B2(n_3326),
.Y(n_3665)
);

OAI21x1_ASAP7_75t_L g3666 ( 
.A1(n_3555),
.A2(n_3571),
.B(n_3559),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3578),
.Y(n_3667)
);

AND2x4_ASAP7_75t_L g3668 ( 
.A(n_3557),
.B(n_3245),
.Y(n_3668)
);

HB1xp67_ASAP7_75t_L g3669 ( 
.A(n_3525),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3530),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3573),
.B(n_3269),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3614),
.B(n_3277),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_3521),
.Y(n_3673)
);

AOI221xp5_ASAP7_75t_L g3674 ( 
.A1(n_3610),
.A2(n_3471),
.B1(n_3358),
.B2(n_3354),
.C(n_3357),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3578),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3600),
.B(n_3277),
.Y(n_3676)
);

AO21x2_ASAP7_75t_L g3677 ( 
.A1(n_3602),
.A2(n_3281),
.B(n_3278),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3566),
.Y(n_3678)
);

INVxp67_ASAP7_75t_SL g3679 ( 
.A(n_3559),
.Y(n_3679)
);

AOI33xp33_ASAP7_75t_L g3680 ( 
.A1(n_3606),
.A2(n_3471),
.A3(n_3309),
.B1(n_3284),
.B2(n_3281),
.B3(n_3285),
.Y(n_3680)
);

OAI33xp33_ASAP7_75t_L g3681 ( 
.A1(n_3562),
.A2(n_3285),
.A3(n_3282),
.B1(n_3284),
.B2(n_3278),
.B3(n_3309),
.Y(n_3681)
);

NAND4xp25_ASAP7_75t_L g3682 ( 
.A(n_3608),
.B(n_3336),
.C(n_3331),
.D(n_3265),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3501),
.B(n_3282),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3604),
.A2(n_3324),
.B1(n_3323),
.B2(n_3446),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_SL g3685 ( 
.A(n_3510),
.B(n_3218),
.Y(n_3685)
);

NAND4xp25_ASAP7_75t_L g3686 ( 
.A(n_3608),
.B(n_3336),
.C(n_3331),
.D(n_3265),
.Y(n_3686)
);

OAI33xp33_ASAP7_75t_L g3687 ( 
.A1(n_3536),
.A2(n_3355),
.A3(n_3303),
.B1(n_3359),
.B2(n_3318),
.B3(n_3304),
.Y(n_3687)
);

OAI211xp5_ASAP7_75t_L g3688 ( 
.A1(n_3612),
.A2(n_3329),
.B(n_3308),
.C(n_3321),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_R g3689 ( 
.A(n_3526),
.B(n_3331),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3580),
.B(n_3318),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3548),
.Y(n_3691)
);

OAI221xp5_ASAP7_75t_L g3692 ( 
.A1(n_3597),
.A2(n_3327),
.B1(n_3461),
.B2(n_3361),
.C(n_3360),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3550),
.Y(n_3693)
);

NAND3xp33_ASAP7_75t_L g3694 ( 
.A(n_3606),
.B(n_3308),
.C(n_3461),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3566),
.Y(n_3695)
);

AND3x1_ASAP7_75t_L g3696 ( 
.A(n_3556),
.B(n_3321),
.C(n_3261),
.Y(n_3696)
);

INVxp67_ASAP7_75t_L g3697 ( 
.A(n_3506),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3604),
.A2(n_3304),
.B1(n_3311),
.B2(n_3296),
.Y(n_3698)
);

OAI211xp5_ASAP7_75t_SL g3699 ( 
.A1(n_3559),
.A2(n_3336),
.B(n_3321),
.C(n_3359),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3553),
.B(n_3321),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3540),
.B(n_3330),
.Y(n_3701)
);

AOI31xp33_ASAP7_75t_L g3702 ( 
.A1(n_3576),
.A2(n_3218),
.A3(n_3330),
.B(n_3296),
.Y(n_3702)
);

INVxp67_ASAP7_75t_L g3703 ( 
.A(n_3506),
.Y(n_3703)
);

OAI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3517),
.A2(n_3317),
.B1(n_3301),
.B2(n_3311),
.Y(n_3704)
);

NOR4xp25_ASAP7_75t_SL g3705 ( 
.A(n_3570),
.B(n_3301),
.C(n_3296),
.D(n_3329),
.Y(n_3705)
);

AOI221xp5_ASAP7_75t_L g3706 ( 
.A1(n_3598),
.A2(n_3301),
.B1(n_3231),
.B2(n_3232),
.C(n_3230),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_L g3707 ( 
.A1(n_3623),
.A2(n_3327),
.B1(n_3221),
.B2(n_3231),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3519),
.B(n_3549),
.Y(n_3708)
);

OAI211xp5_ASAP7_75t_L g3709 ( 
.A1(n_3571),
.A2(n_3308),
.B(n_3301),
.C(n_3216),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3551),
.Y(n_3710)
);

NAND4xp25_ASAP7_75t_L g3711 ( 
.A(n_3608),
.B(n_3320),
.C(n_3216),
.D(n_3308),
.Y(n_3711)
);

AOI22xp33_ASAP7_75t_L g3712 ( 
.A1(n_3583),
.A2(n_3327),
.B1(n_3230),
.B2(n_3232),
.Y(n_3712)
);

NAND2xp33_ASAP7_75t_R g3713 ( 
.A(n_3508),
.B(n_108),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3522),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3554),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_L g3716 ( 
.A(n_3544),
.B(n_3320),
.Y(n_3716)
);

AOI221xp5_ASAP7_75t_L g3717 ( 
.A1(n_3571),
.A2(n_3301),
.B1(n_3221),
.B2(n_3237),
.C(n_3238),
.Y(n_3717)
);

OAI33xp33_ASAP7_75t_L g3718 ( 
.A1(n_3572),
.A2(n_109),
.A3(n_110),
.B1(n_111),
.B2(n_112),
.B3(n_113),
.Y(n_3718)
);

OAI33xp33_ASAP7_75t_L g3719 ( 
.A1(n_3572),
.A2(n_3622),
.A3(n_3579),
.B1(n_3582),
.B2(n_3599),
.B3(n_3616),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3519),
.B(n_3360),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3545),
.B(n_3316),
.Y(n_3721)
);

AO21x2_ASAP7_75t_L g3722 ( 
.A1(n_3582),
.A2(n_3316),
.B(n_3325),
.Y(n_3722)
);

AOI22xp33_ASAP7_75t_L g3723 ( 
.A1(n_3583),
.A2(n_3327),
.B1(n_3237),
.B2(n_3238),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3554),
.Y(n_3724)
);

INVxp67_ASAP7_75t_L g3725 ( 
.A(n_3517),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3576),
.A2(n_3361),
.B(n_3360),
.Y(n_3726)
);

OR2x6_ASAP7_75t_L g3727 ( 
.A(n_3570),
.B(n_3325),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3584),
.A2(n_3249),
.B1(n_3255),
.B2(n_3233),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_SL g3729 ( 
.A1(n_3505),
.A2(n_3361),
.B(n_3360),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3532),
.B(n_3361),
.Y(n_3730)
);

OAI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3622),
.A2(n_3249),
.B1(n_3255),
.B2(n_3233),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3522),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3528),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_R g3734 ( 
.A(n_3508),
.B(n_109),
.Y(n_3734)
);

INVx1_ASAP7_75t_SL g3735 ( 
.A(n_3544),
.Y(n_3735)
);

NAND2xp33_ASAP7_75t_SL g3736 ( 
.A(n_3545),
.B(n_3256),
.Y(n_3736)
);

OR2x2_ASAP7_75t_L g3737 ( 
.A(n_3515),
.B(n_3256),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3539),
.B(n_3257),
.Y(n_3738)
);

AOI22xp33_ASAP7_75t_L g3739 ( 
.A1(n_3584),
.A2(n_3259),
.B1(n_3257),
.B2(n_3402),
.Y(n_3739)
);

OAI22xp33_ASAP7_75t_L g3740 ( 
.A1(n_3581),
.A2(n_3617),
.B1(n_3585),
.B2(n_3555),
.Y(n_3740)
);

AOI211xp5_ASAP7_75t_SL g3741 ( 
.A1(n_3581),
.A2(n_113),
.B(n_110),
.C(n_112),
.Y(n_3741)
);

OR2x2_ASAP7_75t_L g3742 ( 
.A(n_3629),
.B(n_3515),
.Y(n_3742)
);

AOI22xp33_ASAP7_75t_L g3743 ( 
.A1(n_3719),
.A2(n_3589),
.B1(n_3609),
.B2(n_3605),
.Y(n_3743)
);

BUFx2_ASAP7_75t_L g3744 ( 
.A(n_3673),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3677),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3645),
.B(n_3539),
.Y(n_3746)
);

NOR2xp33_ASAP7_75t_L g3747 ( 
.A(n_3638),
.B(n_3585),
.Y(n_3747)
);

OR2x2_ASAP7_75t_L g3748 ( 
.A(n_3639),
.B(n_3546),
.Y(n_3748)
);

OR2x2_ASAP7_75t_L g3749 ( 
.A(n_3671),
.B(n_3518),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3652),
.Y(n_3750)
);

OA211x2_ASAP7_75t_L g3751 ( 
.A1(n_3685),
.A2(n_3542),
.B(n_3533),
.C(n_3531),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3741),
.B(n_3532),
.Y(n_3752)
);

BUFx3_ASAP7_75t_L g3753 ( 
.A(n_3652),
.Y(n_3753)
);

AND2x4_ASAP7_75t_L g3754 ( 
.A(n_3652),
.B(n_3531),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3701),
.B(n_3627),
.Y(n_3755)
);

INVx2_ASAP7_75t_SL g3756 ( 
.A(n_3734),
.Y(n_3756)
);

NAND3xp33_ASAP7_75t_L g3757 ( 
.A(n_3640),
.B(n_3656),
.C(n_3633),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3669),
.Y(n_3758)
);

NAND2x1p5_ASAP7_75t_L g3759 ( 
.A(n_3653),
.B(n_3542),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3719),
.B(n_3531),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3678),
.B(n_3535),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3695),
.B(n_3535),
.Y(n_3762)
);

OAI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3637),
.A2(n_3591),
.B(n_3502),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3715),
.B(n_3502),
.Y(n_3764)
);

NAND3xp33_ASAP7_75t_L g3765 ( 
.A(n_3640),
.B(n_3656),
.C(n_3637),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3649),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3680),
.B(n_3591),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3650),
.Y(n_3768)
);

AO21x2_ASAP7_75t_L g3769 ( 
.A1(n_3679),
.A2(n_3646),
.B(n_3740),
.Y(n_3769)
);

NOR3xp33_ASAP7_75t_SL g3770 ( 
.A(n_3713),
.B(n_3626),
.C(n_3547),
.Y(n_3770)
);

NAND3xp33_ASAP7_75t_L g3771 ( 
.A(n_3642),
.B(n_3628),
.C(n_3635),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3724),
.B(n_3594),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3697),
.B(n_3594),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3655),
.Y(n_3774)
);

NAND3xp33_ASAP7_75t_L g3775 ( 
.A(n_3674),
.B(n_3609),
.C(n_3605),
.Y(n_3775)
);

OR2x2_ASAP7_75t_L g3776 ( 
.A(n_3643),
.B(n_3518),
.Y(n_3776)
);

XOR2x2_ASAP7_75t_L g3777 ( 
.A(n_3651),
.B(n_3588),
.Y(n_3777)
);

NAND3xp33_ASAP7_75t_L g3778 ( 
.A(n_3674),
.B(n_3589),
.C(n_3619),
.Y(n_3778)
);

HB1xp67_ASAP7_75t_L g3779 ( 
.A(n_3697),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3725),
.B(n_3568),
.Y(n_3780)
);

HB1xp67_ASAP7_75t_L g3781 ( 
.A(n_3703),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3630),
.B(n_3528),
.Y(n_3782)
);

AOI211xp5_ASAP7_75t_L g3783 ( 
.A1(n_3631),
.A2(n_3625),
.B(n_3619),
.C(n_3620),
.Y(n_3783)
);

NOR3xp33_ASAP7_75t_L g3784 ( 
.A(n_3718),
.B(n_3603),
.C(n_3547),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3681),
.B(n_3588),
.Y(n_3785)
);

NOR2x1_ASAP7_75t_L g3786 ( 
.A(n_3702),
.B(n_3654),
.Y(n_3786)
);

NOR2x1_ASAP7_75t_L g3787 ( 
.A(n_3654),
.B(n_3547),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3677),
.Y(n_3788)
);

OA211x2_ASAP7_75t_L g3789 ( 
.A1(n_3663),
.A2(n_3558),
.B(n_3503),
.C(n_3625),
.Y(n_3789)
);

CKINVDCx5p33_ASAP7_75t_R g3790 ( 
.A(n_3689),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3735),
.B(n_3568),
.Y(n_3791)
);

NAND3xp33_ASAP7_75t_L g3792 ( 
.A(n_3694),
.B(n_3617),
.C(n_3503),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3666),
.Y(n_3793)
);

AOI22xp33_ASAP7_75t_L g3794 ( 
.A1(n_3718),
.A2(n_3615),
.B1(n_3611),
.B2(n_3537),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3641),
.B(n_3507),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3648),
.B(n_3507),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_3681),
.B(n_3558),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3703),
.B(n_3516),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3660),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3687),
.B(n_3529),
.Y(n_3800)
);

AOI22xp33_ASAP7_75t_L g3801 ( 
.A1(n_3632),
.A2(n_3615),
.B1(n_3611),
.B2(n_3537),
.Y(n_3801)
);

NOR3xp33_ASAP7_75t_SL g3802 ( 
.A(n_3682),
.B(n_3603),
.C(n_3516),
.Y(n_3802)
);

OR2x2_ASAP7_75t_L g3803 ( 
.A(n_3672),
.B(n_3529),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3667),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3675),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3716),
.B(n_3596),
.Y(n_3806)
);

AOI221xp5_ASAP7_75t_L g3807 ( 
.A1(n_3687),
.A2(n_3603),
.B1(n_3523),
.B2(n_3552),
.C(n_3567),
.Y(n_3807)
);

OR2x2_ASAP7_75t_L g3808 ( 
.A(n_3676),
.B(n_3534),
.Y(n_3808)
);

NAND3xp33_ASAP7_75t_L g3809 ( 
.A(n_3692),
.B(n_3564),
.C(n_3523),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3714),
.B(n_3732),
.Y(n_3810)
);

AOI211xp5_ASAP7_75t_L g3811 ( 
.A1(n_3688),
.A2(n_3596),
.B(n_3561),
.C(n_3543),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3683),
.B(n_3708),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3668),
.B(n_3561),
.Y(n_3813)
);

AO21x2_ASAP7_75t_L g3814 ( 
.A1(n_3726),
.A2(n_3541),
.B(n_3586),
.Y(n_3814)
);

NOR3xp33_ASAP7_75t_L g3815 ( 
.A(n_3651),
.B(n_3534),
.C(n_3543),
.Y(n_3815)
);

AOI211xp5_ASAP7_75t_L g3816 ( 
.A1(n_3688),
.A2(n_3541),
.B(n_3565),
.C(n_116),
.Y(n_3816)
);

NAND3xp33_ASAP7_75t_L g3817 ( 
.A(n_3692),
.B(n_3565),
.C(n_3259),
.Y(n_3817)
);

NOR3xp33_ASAP7_75t_L g3818 ( 
.A(n_3709),
.B(n_114),
.C(n_115),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_L g3819 ( 
.A(n_3661),
.B(n_116),
.Y(n_3819)
);

NOR3xp33_ASAP7_75t_L g3820 ( 
.A(n_3709),
.B(n_117),
.C(n_118),
.Y(n_3820)
);

OR2x2_ASAP7_75t_L g3821 ( 
.A(n_3733),
.B(n_3402),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3738),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3668),
.B(n_3402),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3721),
.B(n_3402),
.Y(n_3824)
);

NAND3xp33_ASAP7_75t_L g3825 ( 
.A(n_3726),
.B(n_117),
.C(n_119),
.Y(n_3825)
);

AOI211x1_ASAP7_75t_L g3826 ( 
.A1(n_3711),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3737),
.Y(n_3827)
);

NAND3xp33_ASAP7_75t_L g3828 ( 
.A(n_3706),
.B(n_120),
.C(n_121),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3704),
.B(n_122),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_3707),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3644),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3710),
.B(n_125),
.Y(n_3832)
);

AND2x2_ASAP7_75t_SL g3833 ( 
.A(n_3696),
.B(n_125),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3744),
.B(n_3634),
.Y(n_3834)
);

INVx1_ASAP7_75t_SL g3835 ( 
.A(n_3755),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3814),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3814),
.Y(n_3837)
);

OR2x2_ASAP7_75t_L g3838 ( 
.A(n_3742),
.B(n_3658),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3779),
.Y(n_3839)
);

INVx3_ASAP7_75t_L g3840 ( 
.A(n_3833),
.Y(n_3840)
);

OAI221xp5_ASAP7_75t_L g3841 ( 
.A1(n_3757),
.A2(n_3647),
.B1(n_3665),
.B2(n_3636),
.C(n_3712),
.Y(n_3841)
);

OAI22xp5_ASAP7_75t_L g3842 ( 
.A1(n_3765),
.A2(n_3705),
.B1(n_3727),
.B2(n_3698),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3826),
.A2(n_3727),
.B1(n_3720),
.B2(n_3730),
.Y(n_3843)
);

OAI221xp5_ASAP7_75t_L g3844 ( 
.A1(n_3763),
.A2(n_3723),
.B1(n_3706),
.B2(n_3727),
.C(n_3662),
.Y(n_3844)
);

AOI211xp5_ASAP7_75t_L g3845 ( 
.A1(n_3771),
.A2(n_3686),
.B(n_3664),
.C(n_3699),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3787),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3832),
.B(n_3659),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3786),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3833),
.B(n_3670),
.Y(n_3849)
);

NAND3xp33_ASAP7_75t_L g3850 ( 
.A(n_3818),
.B(n_3693),
.C(n_3691),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3779),
.Y(n_3851)
);

AOI322xp5_ASAP7_75t_L g3852 ( 
.A1(n_3767),
.A2(n_3736),
.A3(n_3731),
.B1(n_3739),
.B2(n_3717),
.C1(n_3684),
.C2(n_3728),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3746),
.B(n_3690),
.Y(n_3853)
);

AOI221x1_ASAP7_75t_L g3854 ( 
.A1(n_3818),
.A2(n_3657),
.B1(n_3699),
.B2(n_3729),
.C(n_3700),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3769),
.Y(n_3855)
);

OAI211xp5_ASAP7_75t_L g3856 ( 
.A1(n_3760),
.A2(n_3717),
.B(n_3722),
.C(n_128),
.Y(n_3856)
);

OAI321xp33_ASAP7_75t_L g3857 ( 
.A1(n_3783),
.A2(n_3722),
.A3(n_127),
.B1(n_129),
.B2(n_130),
.C(n_131),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3764),
.B(n_126),
.Y(n_3858)
);

NAND3xp33_ASAP7_75t_L g3859 ( 
.A(n_3820),
.B(n_126),
.C(n_127),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3781),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3769),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_SL g3862 ( 
.A(n_3820),
.B(n_130),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3781),
.Y(n_3863)
);

AND2x4_ASAP7_75t_L g3864 ( 
.A(n_3754),
.B(n_131),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3747),
.B(n_132),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3782),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3758),
.Y(n_3867)
);

INVx3_ASAP7_75t_L g3868 ( 
.A(n_3754),
.Y(n_3868)
);

INVx2_ASAP7_75t_SL g3869 ( 
.A(n_3750),
.Y(n_3869)
);

INVx2_ASAP7_75t_SL g3870 ( 
.A(n_3750),
.Y(n_3870)
);

AOI221xp5_ASAP7_75t_L g3871 ( 
.A1(n_3785),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.C(n_136),
.Y(n_3871)
);

HB1xp67_ASAP7_75t_L g3872 ( 
.A(n_3780),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3747),
.B(n_133),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3825),
.A2(n_134),
.B(n_135),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_L g3875 ( 
.A1(n_3789),
.A2(n_960),
.B1(n_975),
.B2(n_955),
.Y(n_3875)
);

OR2x2_ASAP7_75t_L g3876 ( 
.A(n_3792),
.B(n_136),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3819),
.B(n_137),
.Y(n_3877)
);

HB1xp67_ASAP7_75t_L g3878 ( 
.A(n_3753),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3745),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3788),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3819),
.B(n_3785),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3766),
.Y(n_3882)
);

AOI33xp33_ASAP7_75t_L g3883 ( 
.A1(n_3816),
.A2(n_139),
.A3(n_140),
.B1(n_141),
.B2(n_142),
.B3(n_143),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3753),
.B(n_140),
.Y(n_3884)
);

AOI221xp5_ASAP7_75t_L g3885 ( 
.A1(n_3797),
.A2(n_3800),
.B1(n_3815),
.B2(n_3760),
.C(n_3784),
.Y(n_3885)
);

NAND3xp33_ASAP7_75t_L g3886 ( 
.A(n_3770),
.B(n_141),
.C(n_142),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_L g3887 ( 
.A1(n_3778),
.A2(n_960),
.B1(n_975),
.B2(n_955),
.Y(n_3887)
);

INVx1_ASAP7_75t_SL g3888 ( 
.A(n_3752),
.Y(n_3888)
);

OR2x2_ASAP7_75t_L g3889 ( 
.A(n_3812),
.B(n_144),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3797),
.A2(n_976),
.B1(n_975),
.B2(n_147),
.Y(n_3890)
);

OAI21xp33_ASAP7_75t_L g3891 ( 
.A1(n_3800),
.A2(n_145),
.B(n_146),
.Y(n_3891)
);

BUFx2_ASAP7_75t_L g3892 ( 
.A(n_3759),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3770),
.B(n_145),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3756),
.Y(n_3894)
);

INVxp67_ASAP7_75t_L g3895 ( 
.A(n_3798),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3768),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3774),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3791),
.B(n_146),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3777),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3795),
.Y(n_3900)
);

AOI221xp5_ASAP7_75t_L g3901 ( 
.A1(n_3815),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_3901)
);

NOR2xp33_ASAP7_75t_L g3902 ( 
.A(n_3790),
.B(n_150),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3813),
.B(n_151),
.Y(n_3903)
);

AND2x4_ASAP7_75t_SL g3904 ( 
.A(n_3761),
.B(n_152),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3806),
.B(n_153),
.Y(n_3905)
);

HB1xp67_ASAP7_75t_L g3906 ( 
.A(n_3793),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3796),
.B(n_154),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3799),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3822),
.B(n_154),
.Y(n_3909)
);

INVx6_ASAP7_75t_L g3910 ( 
.A(n_3829),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3759),
.B(n_155),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3762),
.B(n_155),
.Y(n_3912)
);

INVx1_ASAP7_75t_SL g3913 ( 
.A(n_3748),
.Y(n_3913)
);

INVx2_ASAP7_75t_SL g3914 ( 
.A(n_3773),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_R g3915 ( 
.A(n_3810),
.B(n_157),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3802),
.B(n_158),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3804),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3802),
.B(n_158),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3803),
.Y(n_3919)
);

BUFx3_ASAP7_75t_L g3920 ( 
.A(n_3805),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3808),
.Y(n_3921)
);

INVxp67_ASAP7_75t_SL g3922 ( 
.A(n_3828),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3784),
.B(n_3827),
.Y(n_3923)
);

HB1xp67_ASAP7_75t_L g3924 ( 
.A(n_3772),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3749),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3868),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3903),
.B(n_3776),
.Y(n_3927)
);

NAND2x1_ASAP7_75t_L g3928 ( 
.A(n_3868),
.B(n_3831),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3836),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3903),
.B(n_3811),
.Y(n_3930)
);

OR2x2_ASAP7_75t_L g3931 ( 
.A(n_3872),
.B(n_3743),
.Y(n_3931)
);

OAI32xp33_ASAP7_75t_L g3932 ( 
.A1(n_3840),
.A2(n_3809),
.A3(n_3743),
.B1(n_3830),
.B2(n_3801),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3836),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3905),
.B(n_3830),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3868),
.Y(n_3935)
);

NOR2x1p5_ASAP7_75t_L g3936 ( 
.A(n_3840),
.B(n_3751),
.Y(n_3936)
);

AOI22xp5_ASAP7_75t_L g3937 ( 
.A1(n_3885),
.A2(n_3801),
.B1(n_3775),
.B2(n_3794),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3905),
.B(n_3807),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3837),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3898),
.B(n_3807),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3904),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3837),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3898),
.B(n_3794),
.Y(n_3943)
);

CKINVDCx16_ASAP7_75t_R g3944 ( 
.A(n_3915),
.Y(n_3944)
);

AOI22xp5_ASAP7_75t_L g3945 ( 
.A1(n_3862),
.A2(n_3817),
.B1(n_3821),
.B2(n_3824),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3835),
.B(n_3823),
.Y(n_3946)
);

OAI22xp33_ASAP7_75t_L g3947 ( 
.A1(n_3841),
.A2(n_164),
.B1(n_159),
.B2(n_160),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3907),
.Y(n_3948)
);

OAI22xp5_ASAP7_75t_L g3949 ( 
.A1(n_3881),
.A2(n_164),
.B1(n_159),
.B2(n_160),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3904),
.Y(n_3950)
);

OAI32xp33_ASAP7_75t_L g3951 ( 
.A1(n_3840),
.A2(n_165),
.A3(n_166),
.B1(n_167),
.B2(n_170),
.Y(n_3951)
);

INVx3_ASAP7_75t_SL g3952 ( 
.A(n_3864),
.Y(n_3952)
);

OR2x2_ASAP7_75t_L g3953 ( 
.A(n_3913),
.B(n_165),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3912),
.Y(n_3954)
);

OR2x2_ASAP7_75t_L g3955 ( 
.A(n_3919),
.B(n_166),
.Y(n_3955)
);

OAI21xp33_ASAP7_75t_SL g3956 ( 
.A1(n_3855),
.A2(n_167),
.B(n_170),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3855),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3907),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3912),
.Y(n_3959)
);

AND2x4_ASAP7_75t_L g3960 ( 
.A(n_3869),
.B(n_173),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3839),
.Y(n_3961)
);

NOR2xp33_ASAP7_75t_L g3962 ( 
.A(n_3864),
.B(n_174),
.Y(n_3962)
);

AOI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3862),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3851),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3860),
.Y(n_3965)
);

OA222x2_ASAP7_75t_L g3966 ( 
.A1(n_3861),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.C1(n_179),
.C2(n_180),
.Y(n_3966)
);

AND2x2_ASAP7_75t_L g3967 ( 
.A(n_3853),
.B(n_179),
.Y(n_3967)
);

OAI33xp33_ASAP7_75t_L g3968 ( 
.A1(n_3923),
.A2(n_181),
.A3(n_182),
.B1(n_183),
.B2(n_184),
.B3(n_186),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3865),
.B(n_181),
.Y(n_3969)
);

OR2x2_ASAP7_75t_L g3970 ( 
.A(n_3919),
.B(n_182),
.Y(n_3970)
);

INVxp67_ASAP7_75t_L g3971 ( 
.A(n_3878),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3863),
.Y(n_3972)
);

OAI22xp33_ASAP7_75t_SL g3973 ( 
.A1(n_3861),
.A2(n_3893),
.B1(n_3848),
.B2(n_3876),
.Y(n_3973)
);

OR2x6_ASAP7_75t_L g3974 ( 
.A(n_3894),
.B(n_183),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3864),
.Y(n_3975)
);

NAND2x2_ASAP7_75t_L g3976 ( 
.A(n_3869),
.B(n_184),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3889),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3838),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3884),
.Y(n_3979)
);

OA222x2_ASAP7_75t_L g3980 ( 
.A1(n_3848),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.C1(n_190),
.C2(n_191),
.Y(n_3980)
);

AOI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3891),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3906),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3834),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3834),
.Y(n_3984)
);

OAI32xp33_ASAP7_75t_L g3985 ( 
.A1(n_3886),
.A2(n_193),
.A3(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3866),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3858),
.Y(n_3987)
);

HB1xp67_ASAP7_75t_L g3988 ( 
.A(n_3915),
.Y(n_3988)
);

AOI22xp5_ASAP7_75t_L g3989 ( 
.A1(n_3893),
.A2(n_198),
.B1(n_195),
.B2(n_197),
.Y(n_3989)
);

OR2x2_ASAP7_75t_L g3990 ( 
.A(n_3921),
.B(n_197),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3879),
.Y(n_3991)
);

OAI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3890),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3884),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3879),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3880),
.Y(n_3995)
);

NAND4xp25_ASAP7_75t_L g3996 ( 
.A(n_3871),
.B(n_202),
.C(n_199),
.D(n_200),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3853),
.B(n_3894),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3900),
.B(n_202),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3880),
.Y(n_3999)
);

OR2x2_ASAP7_75t_L g4000 ( 
.A(n_3921),
.B(n_203),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3865),
.B(n_204),
.Y(n_4001)
);

AND2x4_ASAP7_75t_SL g4002 ( 
.A(n_3900),
.B(n_204),
.Y(n_4002)
);

INVx2_ASAP7_75t_SL g4003 ( 
.A(n_3870),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3873),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3873),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3910),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3888),
.B(n_205),
.Y(n_4007)
);

HB1xp67_ASAP7_75t_L g4008 ( 
.A(n_3870),
.Y(n_4008)
);

INVx2_ASAP7_75t_SL g4009 ( 
.A(n_3911),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3925),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3909),
.Y(n_4011)
);

INVxp67_ASAP7_75t_SL g4012 ( 
.A(n_3902),
.Y(n_4012)
);

OR2x2_ASAP7_75t_L g4013 ( 
.A(n_3876),
.B(n_205),
.Y(n_4013)
);

OAI33xp33_ASAP7_75t_L g4014 ( 
.A1(n_3842),
.A2(n_206),
.A3(n_207),
.B1(n_208),
.B2(n_210),
.B3(n_211),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3883),
.B(n_207),
.Y(n_4015)
);

BUFx2_ASAP7_75t_L g4016 ( 
.A(n_3997),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3988),
.Y(n_4017)
);

BUFx2_ASAP7_75t_L g4018 ( 
.A(n_3960),
.Y(n_4018)
);

INVx1_ASAP7_75t_SL g4019 ( 
.A(n_3944),
.Y(n_4019)
);

NAND4xp25_ASAP7_75t_L g4020 ( 
.A(n_3937),
.B(n_3845),
.C(n_3854),
.D(n_3892),
.Y(n_4020)
);

AND2x4_ASAP7_75t_L g4021 ( 
.A(n_4006),
.B(n_3920),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3936),
.B(n_3911),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3960),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3937),
.B(n_3922),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3967),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3927),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3946),
.B(n_3924),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3983),
.B(n_3916),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_4004),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_4012),
.B(n_3916),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_4005),
.Y(n_4031)
);

NOR2xp33_ASAP7_75t_SL g4032 ( 
.A(n_4008),
.B(n_3902),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3948),
.Y(n_4033)
);

NOR2xp33_ASAP7_75t_L g4034 ( 
.A(n_3952),
.B(n_3910),
.Y(n_4034)
);

INVx1_ASAP7_75t_SL g4035 ( 
.A(n_4002),
.Y(n_4035)
);

NAND2xp33_ASAP7_75t_R g4036 ( 
.A(n_3974),
.B(n_3918),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3958),
.Y(n_4037)
);

OR2x2_ASAP7_75t_L g4038 ( 
.A(n_3984),
.B(n_3914),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3973),
.A2(n_3857),
.B(n_3856),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_4009),
.B(n_3883),
.Y(n_4040)
);

NOR2xp33_ASAP7_75t_L g4041 ( 
.A(n_3968),
.B(n_3910),
.Y(n_4041)
);

OR2x2_ASAP7_75t_L g4042 ( 
.A(n_3931),
.B(n_3914),
.Y(n_4042)
);

OR2x2_ASAP7_75t_L g4043 ( 
.A(n_3959),
.B(n_3847),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_4003),
.B(n_3918),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3954),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3969),
.Y(n_4046)
);

HB1xp67_ASAP7_75t_L g4047 ( 
.A(n_3974),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3963),
.B(n_3849),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_4001),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_4013),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3930),
.B(n_3849),
.Y(n_4051)
);

NOR2xp33_ASAP7_75t_L g4052 ( 
.A(n_3975),
.B(n_3877),
.Y(n_4052)
);

INVxp67_ASAP7_75t_SL g4053 ( 
.A(n_3973),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3953),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3955),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_3978),
.B(n_3895),
.Y(n_4056)
);

INVx1_ASAP7_75t_SL g4057 ( 
.A(n_4007),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3970),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3926),
.B(n_3867),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3979),
.B(n_3920),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3993),
.B(n_3998),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3935),
.B(n_3850),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3990),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3971),
.B(n_3843),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3963),
.B(n_3901),
.Y(n_4065)
);

INVxp67_ASAP7_75t_L g4066 ( 
.A(n_3962),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_3941),
.B(n_3882),
.Y(n_4067)
);

AND2x2_ASAP7_75t_SL g4068 ( 
.A(n_3940),
.B(n_3875),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3950),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_4000),
.Y(n_4070)
);

CKINVDCx16_ASAP7_75t_R g4071 ( 
.A(n_3977),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3976),
.Y(n_4072)
);

NOR2xp67_ASAP7_75t_L g4073 ( 
.A(n_3982),
.B(n_3844),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_3986),
.B(n_3896),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_3989),
.B(n_3859),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3929),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_4010),
.B(n_3897),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3961),
.B(n_3908),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3938),
.B(n_3846),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_L g4080 ( 
.A(n_3989),
.B(n_3846),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3987),
.B(n_3917),
.Y(n_4081)
);

OR2x2_ASAP7_75t_L g4082 ( 
.A(n_3943),
.B(n_3874),
.Y(n_4082)
);

OAI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_3956),
.A2(n_3899),
.B(n_3852),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_4011),
.B(n_3899),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3957),
.B(n_3887),
.Y(n_4085)
);

OAI322xp33_ASAP7_75t_L g4086 ( 
.A1(n_3945),
.A2(n_212),
.A3(n_213),
.B1(n_215),
.B2(n_216),
.C1(n_217),
.C2(n_218),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3933),
.Y(n_4087)
);

OAI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_3956),
.A2(n_215),
.B(n_216),
.Y(n_4088)
);

OAI33xp33_ASAP7_75t_L g4089 ( 
.A1(n_3947),
.A2(n_217),
.A3(n_218),
.B1(n_219),
.B2(n_220),
.B3(n_222),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3928),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3939),
.Y(n_4091)
);

NOR2xp33_ASAP7_75t_L g4092 ( 
.A(n_4014),
.B(n_219),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3964),
.B(n_220),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3934),
.B(n_223),
.Y(n_4094)
);

BUFx2_ASAP7_75t_L g4095 ( 
.A(n_3965),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3942),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3981),
.B(n_224),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_3972),
.B(n_224),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_3991),
.B(n_225),
.Y(n_4099)
);

INVx1_ASAP7_75t_SL g4100 ( 
.A(n_4016),
.Y(n_4100)
);

NOR2xp33_ASAP7_75t_L g4101 ( 
.A(n_4019),
.B(n_3932),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4053),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_4019),
.B(n_4015),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_4071),
.B(n_4026),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_4032),
.B(n_3999),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_L g4106 ( 
.A(n_4024),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4018),
.Y(n_4107)
);

INVx1_ASAP7_75t_SL g4108 ( 
.A(n_4051),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4032),
.B(n_3981),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_4021),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4047),
.Y(n_4111)
);

AND2x2_ASAP7_75t_L g4112 ( 
.A(n_4027),
.B(n_3945),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_4021),
.B(n_3949),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4023),
.B(n_3996),
.Y(n_4114)
);

INVx2_ASAP7_75t_SL g4115 ( 
.A(n_4069),
.Y(n_4115)
);

OAI21xp33_ASAP7_75t_L g4116 ( 
.A1(n_4020),
.A2(n_3985),
.B(n_3992),
.Y(n_4116)
);

INVxp67_ASAP7_75t_SL g4117 ( 
.A(n_4024),
.Y(n_4117)
);

OR2x2_ASAP7_75t_L g4118 ( 
.A(n_4042),
.B(n_3994),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4022),
.B(n_3966),
.Y(n_4119)
);

INVx2_ASAP7_75t_SL g4120 ( 
.A(n_4090),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_4025),
.B(n_3951),
.Y(n_4121)
);

INVx1_ASAP7_75t_SL g4122 ( 
.A(n_4035),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_4044),
.B(n_4028),
.Y(n_4123)
);

OR2x2_ASAP7_75t_L g4124 ( 
.A(n_4038),
.B(n_3995),
.Y(n_4124)
);

OR2x2_ASAP7_75t_L g4125 ( 
.A(n_4030),
.B(n_3966),
.Y(n_4125)
);

OAI21xp5_ASAP7_75t_SL g4126 ( 
.A1(n_4039),
.A2(n_3980),
.B(n_225),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4099),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_4061),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_4035),
.B(n_3980),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_4030),
.B(n_227),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4093),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_4034),
.B(n_227),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_4099),
.B(n_4098),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_4052),
.B(n_229),
.Y(n_4134)
);

NOR2x1_ASAP7_75t_L g4135 ( 
.A(n_4060),
.B(n_231),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4095),
.Y(n_4136)
);

NOR2x1p5_ASAP7_75t_L g4137 ( 
.A(n_4017),
.B(n_231),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_4056),
.B(n_232),
.Y(n_4138)
);

CKINVDCx5p33_ASAP7_75t_R g4139 ( 
.A(n_4057),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4094),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4050),
.Y(n_4141)
);

AOI322xp5_ASAP7_75t_L g4142 ( 
.A1(n_4079),
.A2(n_4041),
.A3(n_4048),
.B1(n_4084),
.B2(n_4075),
.C1(n_4080),
.C2(n_4072),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_4057),
.B(n_232),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4059),
.Y(n_4144)
);

OAI31xp33_ASAP7_75t_L g4145 ( 
.A1(n_4079),
.A2(n_4048),
.A3(n_4080),
.B(n_4082),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_4092),
.B(n_233),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4054),
.B(n_234),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_4063),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_4064),
.B(n_234),
.Y(n_4149)
);

NAND2x1_ASAP7_75t_SL g4150 ( 
.A(n_4062),
.B(n_235),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4067),
.B(n_236),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4067),
.B(n_237),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_4078),
.B(n_237),
.Y(n_4153)
);

AND2x2_ASAP7_75t_L g4154 ( 
.A(n_4029),
.B(n_238),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4043),
.Y(n_4155)
);

INVx1_ASAP7_75t_SL g4156 ( 
.A(n_4040),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4046),
.B(n_238),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4055),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4049),
.B(n_239),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4058),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4066),
.B(n_240),
.Y(n_4161)
);

AND2x4_ASAP7_75t_L g4162 ( 
.A(n_4045),
.B(n_4031),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4068),
.B(n_240),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4033),
.B(n_241),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_4037),
.B(n_241),
.Y(n_4165)
);

OR2x2_ASAP7_75t_L g4166 ( 
.A(n_4074),
.B(n_242),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4139),
.Y(n_4167)
);

OAI221xp5_ASAP7_75t_L g4168 ( 
.A1(n_4102),
.A2(n_4083),
.B1(n_4073),
.B2(n_4036),
.C(n_4065),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_4115),
.B(n_4108),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4139),
.Y(n_4170)
);

AND2x2_ASAP7_75t_SL g4171 ( 
.A(n_4112),
.B(n_4084),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_4117),
.A2(n_4086),
.B(n_4083),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_4150),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4115),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_4100),
.B(n_4077),
.Y(n_4175)
);

AOI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_4101),
.A2(n_4065),
.B1(n_4070),
.B2(n_4091),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4110),
.Y(n_4177)
);

O2A1O1Ixp33_ASAP7_75t_L g4178 ( 
.A1(n_4106),
.A2(n_4097),
.B(n_4096),
.C(n_4087),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4106),
.B(n_4088),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4110),
.Y(n_4180)
);

NAND3xp33_ASAP7_75t_L g4181 ( 
.A(n_4145),
.B(n_4076),
.C(n_4088),
.Y(n_4181)
);

AOI31xp33_ASAP7_75t_L g4182 ( 
.A1(n_4122),
.A2(n_4081),
.A3(n_4089),
.B(n_4085),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4104),
.Y(n_4183)
);

NOR4xp25_ASAP7_75t_L g4184 ( 
.A(n_4117),
.B(n_4081),
.C(n_4085),
.D(n_244),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4153),
.B(n_4138),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4163),
.Y(n_4186)
);

OR4x1_ASAP7_75t_L g4187 ( 
.A(n_4120),
.B(n_242),
.C(n_243),
.D(n_245),
.Y(n_4187)
);

O2A1O1Ixp33_ASAP7_75t_L g4188 ( 
.A1(n_4105),
.A2(n_243),
.B(n_247),
.C(n_250),
.Y(n_4188)
);

OAI221xp5_ASAP7_75t_L g4189 ( 
.A1(n_4101),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.C(n_254),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4151),
.B(n_251),
.Y(n_4190)
);

INVx2_ASAP7_75t_SL g4191 ( 
.A(n_4152),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4118),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_4135),
.B(n_253),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4105),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4127),
.B(n_254),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_4127),
.B(n_4149),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4156),
.A2(n_976),
.B1(n_975),
.B2(n_1427),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4119),
.B(n_256),
.Y(n_4198)
);

AOI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_4109),
.A2(n_256),
.B(n_257),
.Y(n_4199)
);

AOI211xp5_ASAP7_75t_L g4200 ( 
.A1(n_4112),
.A2(n_258),
.B(n_259),
.C(n_261),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_4126),
.B(n_258),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4123),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_4116),
.A2(n_259),
.B(n_265),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4137),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4166),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_4103),
.A2(n_976),
.B1(n_1427),
.B2(n_267),
.Y(n_4206)
);

INVx1_ASAP7_75t_SL g4207 ( 
.A(n_4124),
.Y(n_4207)
);

AOI21xp33_ASAP7_75t_L g4208 ( 
.A1(n_4129),
.A2(n_265),
.B(n_266),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4154),
.Y(n_4209)
);

OAI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_4107),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4125),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4134),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4162),
.Y(n_4213)
);

A2O1A1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_4142),
.A2(n_270),
.B(n_271),
.C(n_272),
.Y(n_4214)
);

OR2x2_ASAP7_75t_L g4215 ( 
.A(n_4144),
.B(n_271),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4162),
.Y(n_4216)
);

AOI221xp5_ASAP7_75t_L g4217 ( 
.A1(n_4129),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.C(n_275),
.Y(n_4217)
);

HB1xp67_ASAP7_75t_L g4218 ( 
.A(n_4162),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4148),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_4155),
.B(n_275),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4148),
.Y(n_4221)
);

NAND3xp33_ASAP7_75t_L g4222 ( 
.A(n_4136),
.B(n_276),
.C(n_277),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_4133),
.B(n_276),
.Y(n_4223)
);

NAND4xp25_ASAP7_75t_SL g4224 ( 
.A(n_4113),
.B(n_277),
.C(n_278),
.D(n_279),
.Y(n_4224)
);

INVx1_ASAP7_75t_SL g4225 ( 
.A(n_4132),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4132),
.B(n_4128),
.Y(n_4226)
);

AO22x1_ASAP7_75t_L g4227 ( 
.A1(n_4120),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4143),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_SL g4229 ( 
.A1(n_4111),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4130),
.Y(n_4230)
);

OAI33xp33_ASAP7_75t_L g4231 ( 
.A1(n_4121),
.A2(n_283),
.A3(n_285),
.B1(n_286),
.B2(n_287),
.B3(n_288),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4131),
.Y(n_4232)
);

OAI22xp5_ASAP7_75t_L g4233 ( 
.A1(n_4207),
.A2(n_4141),
.B1(n_4160),
.B2(n_4158),
.Y(n_4233)
);

XOR2x2_ASAP7_75t_L g4234 ( 
.A(n_4171),
.B(n_4114),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4225),
.B(n_4140),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4218),
.Y(n_4236)
);

HB1xp67_ASAP7_75t_L g4237 ( 
.A(n_4168),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4207),
.B(n_4164),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_4225),
.B(n_4165),
.Y(n_4239)
);

XNOR2x2_ASAP7_75t_L g4240 ( 
.A(n_4181),
.B(n_4146),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4202),
.B(n_4147),
.Y(n_4241)
);

BUFx3_ASAP7_75t_L g4242 ( 
.A(n_4213),
.Y(n_4242)
);

OAI322xp33_ASAP7_75t_L g4243 ( 
.A1(n_4172),
.A2(n_4159),
.A3(n_4157),
.B1(n_4161),
.B2(n_291),
.C1(n_292),
.C2(n_293),
.Y(n_4243)
);

AND2x2_ASAP7_75t_L g4244 ( 
.A(n_4169),
.B(n_287),
.Y(n_4244)
);

INVxp67_ASAP7_75t_L g4245 ( 
.A(n_4226),
.Y(n_4245)
);

INVxp67_ASAP7_75t_L g4246 ( 
.A(n_4196),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_4227),
.B(n_289),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_L g4248 ( 
.A(n_4231),
.B(n_289),
.Y(n_4248)
);

AOI221xp5_ASAP7_75t_L g4249 ( 
.A1(n_4184),
.A2(n_290),
.B1(n_292),
.B2(n_294),
.C(n_296),
.Y(n_4249)
);

OAI22xp33_ASAP7_75t_L g4250 ( 
.A1(n_4182),
.A2(n_290),
.B1(n_294),
.B2(n_297),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4184),
.B(n_297),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4200),
.B(n_298),
.Y(n_4252)
);

NAND4xp25_ASAP7_75t_L g4253 ( 
.A(n_4175),
.B(n_298),
.C(n_299),
.D(n_301),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4200),
.B(n_299),
.Y(n_4254)
);

XNOR2x2_ASAP7_75t_L g4255 ( 
.A(n_4181),
.B(n_301),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4187),
.Y(n_4256)
);

OA22x2_ASAP7_75t_L g4257 ( 
.A1(n_4176),
.A2(n_302),
.B1(n_305),
.B2(n_306),
.Y(n_4257)
);

INVx1_ASAP7_75t_SL g4258 ( 
.A(n_4179),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4192),
.B(n_302),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4216),
.B(n_4180),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_4191),
.B(n_305),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_4219),
.B(n_308),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_SL g4263 ( 
.A(n_4221),
.B(n_308),
.Y(n_4263)
);

OAI21xp33_ASAP7_75t_L g4264 ( 
.A1(n_4167),
.A2(n_4170),
.B(n_4211),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4177),
.Y(n_4265)
);

INVx1_ASAP7_75t_SL g4266 ( 
.A(n_4185),
.Y(n_4266)
);

AOI321xp33_ASAP7_75t_R g4267 ( 
.A1(n_4178),
.A2(n_309),
.A3(n_310),
.B1(n_311),
.B2(n_312),
.C(n_313),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4174),
.B(n_310),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4198),
.Y(n_4269)
);

XNOR2xp5_ASAP7_75t_L g4270 ( 
.A(n_4173),
.B(n_312),
.Y(n_4270)
);

AOI21xp33_ASAP7_75t_L g4271 ( 
.A1(n_4204),
.A2(n_314),
.B(n_316),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_4215),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4220),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4183),
.B(n_316),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4194),
.B(n_317),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4193),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4190),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4230),
.Y(n_4278)
);

OAI221xp5_ASAP7_75t_SL g4279 ( 
.A1(n_4214),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.C(n_320),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4205),
.B(n_318),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4209),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4195),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4232),
.B(n_319),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4229),
.B(n_4201),
.Y(n_4284)
);

AND2x2_ASAP7_75t_L g4285 ( 
.A(n_4223),
.B(n_321),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4212),
.B(n_321),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4222),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4257),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4256),
.B(n_4199),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_4242),
.B(n_4186),
.Y(n_4290)
);

AOI22xp5_ASAP7_75t_L g4291 ( 
.A1(n_4258),
.A2(n_4228),
.B1(n_4217),
.B2(n_4224),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4260),
.B(n_4222),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4256),
.B(n_4203),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4242),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4245),
.B(n_4188),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4245),
.B(n_4210),
.Y(n_4296)
);

NOR2x1_ASAP7_75t_L g4297 ( 
.A(n_4236),
.B(n_4189),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_4266),
.B(n_4208),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_L g4299 ( 
.A(n_4246),
.B(n_4206),
.Y(n_4299)
);

INVx1_ASAP7_75t_SL g4300 ( 
.A(n_4234),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4257),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4255),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_4250),
.B(n_4197),
.Y(n_4303)
);

HB1xp67_ASAP7_75t_L g4304 ( 
.A(n_4246),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4251),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4270),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4244),
.B(n_323),
.Y(n_4307)
);

OR2x2_ASAP7_75t_L g4308 ( 
.A(n_4235),
.B(n_327),
.Y(n_4308)
);

XNOR2xp5_ASAP7_75t_L g4309 ( 
.A(n_4240),
.B(n_329),
.Y(n_4309)
);

AND4x1_ASAP7_75t_L g4310 ( 
.A(n_4239),
.B(n_330),
.C(n_331),
.D(n_332),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4275),
.Y(n_4311)
);

XNOR2xp5_ASAP7_75t_L g4312 ( 
.A(n_4250),
.B(n_333),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4238),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4274),
.Y(n_4314)
);

AOI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4239),
.A2(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_4285),
.B(n_336),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4247),
.Y(n_4317)
);

OAI211xp5_ASAP7_75t_L g4318 ( 
.A1(n_4264),
.A2(n_337),
.B(n_338),
.C(n_340),
.Y(n_4318)
);

XNOR2xp5_ASAP7_75t_L g4319 ( 
.A(n_4267),
.B(n_337),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4273),
.Y(n_4320)
);

OR2x6_ASAP7_75t_L g4321 ( 
.A(n_4281),
.B(n_338),
.Y(n_4321)
);

OAI211xp5_ASAP7_75t_L g4322 ( 
.A1(n_4237),
.A2(n_4265),
.B(n_4241),
.C(n_4287),
.Y(n_4322)
);

AOI21xp33_ASAP7_75t_SL g4323 ( 
.A1(n_4262),
.A2(n_340),
.B(n_341),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4273),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4237),
.B(n_4268),
.Y(n_4325)
);

O2A1O1Ixp33_ASAP7_75t_L g4326 ( 
.A1(n_4262),
.A2(n_341),
.B(n_342),
.C(n_343),
.Y(n_4326)
);

BUFx2_ASAP7_75t_L g4327 ( 
.A(n_4281),
.Y(n_4327)
);

NAND4xp25_ASAP7_75t_L g4328 ( 
.A(n_4284),
.B(n_342),
.C(n_343),
.D(n_344),
.Y(n_4328)
);

AOI211x1_ASAP7_75t_L g4329 ( 
.A1(n_4322),
.A2(n_4233),
.B(n_4278),
.C(n_4263),
.Y(n_4329)
);

AOI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_4327),
.A2(n_4263),
.B(n_4261),
.Y(n_4330)
);

NOR2xp33_ASAP7_75t_L g4331 ( 
.A(n_4294),
.B(n_4243),
.Y(n_4331)
);

OAI21xp33_ASAP7_75t_SL g4332 ( 
.A1(n_4300),
.A2(n_4249),
.B(n_4269),
.Y(n_4332)
);

NOR3xp33_ASAP7_75t_L g4333 ( 
.A(n_4325),
.B(n_4280),
.C(n_4276),
.Y(n_4333)
);

INVx1_ASAP7_75t_SL g4334 ( 
.A(n_4292),
.Y(n_4334)
);

NOR2x1_ASAP7_75t_L g4335 ( 
.A(n_4290),
.B(n_4253),
.Y(n_4335)
);

BUFx12f_ASAP7_75t_L g4336 ( 
.A(n_4290),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_4304),
.B(n_4279),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4309),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4289),
.A2(n_4279),
.B(n_4252),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_4302),
.B(n_4323),
.Y(n_4340)
);

INVxp67_ASAP7_75t_L g4341 ( 
.A(n_4321),
.Y(n_4341)
);

OAI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_4313),
.A2(n_4248),
.B1(n_4254),
.B2(n_4259),
.Y(n_4342)
);

INVx2_ASAP7_75t_SL g4343 ( 
.A(n_4308),
.Y(n_4343)
);

NOR3x1_ASAP7_75t_L g4344 ( 
.A(n_4296),
.B(n_4318),
.C(n_4293),
.Y(n_4344)
);

OA22x2_ASAP7_75t_L g4345 ( 
.A1(n_4291),
.A2(n_4272),
.B1(n_4277),
.B2(n_4283),
.Y(n_4345)
);

AOI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_4295),
.A2(n_4248),
.B(n_4271),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4320),
.B(n_4286),
.Y(n_4347)
);

AOI22xp5_ASAP7_75t_L g4348 ( 
.A1(n_4317),
.A2(n_4282),
.B1(n_347),
.B2(n_348),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4297),
.A2(n_346),
.B(n_349),
.Y(n_4349)
);

OAI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4324),
.A2(n_4298),
.B1(n_4319),
.B2(n_4297),
.Y(n_4350)
);

AOI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_4305),
.A2(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_SL g4352 ( 
.A(n_4323),
.B(n_352),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_L g4353 ( 
.A(n_4310),
.B(n_353),
.Y(n_4353)
);

AOI22xp33_ASAP7_75t_L g4354 ( 
.A1(n_4333),
.A2(n_4288),
.B1(n_4301),
.B2(n_4311),
.Y(n_4354)
);

AOI311xp33_ASAP7_75t_L g4355 ( 
.A1(n_4331),
.A2(n_4299),
.A3(n_4306),
.B(n_4314),
.C(n_4303),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4336),
.Y(n_4356)
);

NOR2x1_ASAP7_75t_SL g4357 ( 
.A(n_4337),
.B(n_4321),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4347),
.Y(n_4358)
);

AOI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4334),
.A2(n_4307),
.B1(n_4316),
.B2(n_4328),
.Y(n_4359)
);

OA22x2_ASAP7_75t_L g4360 ( 
.A1(n_4348),
.A2(n_4312),
.B1(n_4315),
.B2(n_4326),
.Y(n_4360)
);

AOI222xp33_ASAP7_75t_L g4361 ( 
.A1(n_4350),
.A2(n_353),
.B1(n_354),
.B2(n_356),
.C1(n_357),
.C2(n_358),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4329),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4335),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_4340),
.A2(n_4330),
.B(n_4352),
.Y(n_4364)
);

XNOR2xp5_ASAP7_75t_L g4365 ( 
.A(n_4345),
.B(n_354),
.Y(n_4365)
);

OAI32xp33_ASAP7_75t_L g4366 ( 
.A1(n_4332),
.A2(n_356),
.A3(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_SL g4367 ( 
.A(n_4349),
.B(n_360),
.Y(n_4367)
);

A2O1A1Ixp33_ASAP7_75t_SL g4368 ( 
.A1(n_4338),
.A2(n_361),
.B(n_362),
.C(n_363),
.Y(n_4368)
);

OAI31xp33_ASAP7_75t_L g4369 ( 
.A1(n_4342),
.A2(n_361),
.A3(n_363),
.B(n_364),
.Y(n_4369)
);

XOR2xp5_ASAP7_75t_L g4370 ( 
.A(n_4356),
.B(n_4346),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_4362),
.A2(n_4353),
.B1(n_4343),
.B2(n_4341),
.Y(n_4371)
);

NOR2x1_ASAP7_75t_L g4372 ( 
.A(n_4358),
.B(n_4363),
.Y(n_4372)
);

AOI22xp5_ASAP7_75t_L g4373 ( 
.A1(n_4359),
.A2(n_4339),
.B1(n_4351),
.B2(n_4344),
.Y(n_4373)
);

AOI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4354),
.A2(n_976),
.B1(n_372),
.B2(n_375),
.Y(n_4374)
);

AOI22xp5_ASAP7_75t_L g4375 ( 
.A1(n_4360),
.A2(n_366),
.B1(n_376),
.B2(n_378),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4365),
.Y(n_4376)
);

AOI221xp5_ASAP7_75t_L g4377 ( 
.A1(n_4364),
.A2(n_379),
.B1(n_380),
.B2(n_382),
.C(n_383),
.Y(n_4377)
);

AOI22xp5_ASAP7_75t_L g4378 ( 
.A1(n_4367),
.A2(n_385),
.B1(n_388),
.B2(n_389),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4357),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4366),
.Y(n_4380)
);

INVxp33_ASAP7_75t_L g4381 ( 
.A(n_4372),
.Y(n_4381)
);

AOI322xp5_ASAP7_75t_L g4382 ( 
.A1(n_4376),
.A2(n_4355),
.A3(n_4368),
.B1(n_4369),
.B2(n_4361),
.C1(n_399),
.C2(n_401),
.Y(n_4382)
);

AOI322xp5_ASAP7_75t_L g4383 ( 
.A1(n_4379),
.A2(n_489),
.A3(n_394),
.B1(n_395),
.B2(n_397),
.C1(n_406),
.C2(n_407),
.Y(n_4383)
);

INVxp33_ASAP7_75t_L g4384 ( 
.A(n_4370),
.Y(n_4384)
);

OR2x2_ASAP7_75t_L g4385 ( 
.A(n_4380),
.B(n_391),
.Y(n_4385)
);

BUFx2_ASAP7_75t_L g4386 ( 
.A(n_4373),
.Y(n_4386)
);

AOI22xp5_ASAP7_75t_L g4387 ( 
.A1(n_4371),
.A2(n_409),
.B1(n_411),
.B2(n_414),
.Y(n_4387)
);

NOR2x1p5_ASAP7_75t_L g4388 ( 
.A(n_4385),
.B(n_4381),
.Y(n_4388)
);

NOR2x1_ASAP7_75t_L g4389 ( 
.A(n_4386),
.B(n_4374),
.Y(n_4389)
);

AND4x1_ASAP7_75t_L g4390 ( 
.A(n_4387),
.B(n_4375),
.C(n_4378),
.D(n_4377),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4384),
.Y(n_4391)
);

NOR2x1_ASAP7_75t_L g4392 ( 
.A(n_4382),
.B(n_415),
.Y(n_4392)
);

O2A1O1Ixp33_ASAP7_75t_L g4393 ( 
.A1(n_4391),
.A2(n_4383),
.B(n_417),
.C(n_418),
.Y(n_4393)
);

OAI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4392),
.A2(n_416),
.B1(n_422),
.B2(n_423),
.Y(n_4394)
);

INVx4_ASAP7_75t_L g4395 ( 
.A(n_4394),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4393),
.B(n_4388),
.Y(n_4396)
);

HB1xp67_ASAP7_75t_L g4397 ( 
.A(n_4396),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_4397),
.B(n_4389),
.Y(n_4398)
);

NAND4xp75_ASAP7_75t_L g4399 ( 
.A(n_4398),
.B(n_4395),
.C(n_4390),
.D(n_432),
.Y(n_4399)
);

OAI22x1_ASAP7_75t_L g4400 ( 
.A1(n_4399),
.A2(n_427),
.B1(n_429),
.B2(n_437),
.Y(n_4400)
);

INVx1_ASAP7_75t_SL g4401 ( 
.A(n_4400),
.Y(n_4401)
);

AOI222xp33_ASAP7_75t_SL g4402 ( 
.A1(n_4401),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.C1(n_444),
.C2(n_447),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4402),
.Y(n_4403)
);

AOI221xp5_ASAP7_75t_L g4404 ( 
.A1(n_4403),
.A2(n_449),
.B1(n_450),
.B2(n_453),
.C(n_456),
.Y(n_4404)
);

AOI31xp33_ASAP7_75t_L g4405 ( 
.A1(n_4403),
.A2(n_458),
.A3(n_460),
.B(n_461),
.Y(n_4405)
);

AOI22xp5_ASAP7_75t_SL g4406 ( 
.A1(n_4405),
.A2(n_463),
.B1(n_464),
.B2(n_468),
.Y(n_4406)
);

AOI22xp33_ASAP7_75t_L g4407 ( 
.A1(n_4404),
.A2(n_469),
.B1(n_471),
.B2(n_474),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4406),
.Y(n_4408)
);

AOI21xp5_ASAP7_75t_L g4409 ( 
.A1(n_4408),
.A2(n_4407),
.B(n_478),
.Y(n_4409)
);

AOI211xp5_ASAP7_75t_L g4410 ( 
.A1(n_4409),
.A2(n_475),
.B(n_479),
.C(n_488),
.Y(n_4410)
);


endmodule