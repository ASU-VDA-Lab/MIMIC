module real_jpeg_20524_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_1),
.A2(n_5),
.B1(n_24),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_3),
.B1(n_39),
.B2(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_5),
.B1(n_24),
.B2(n_39),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_44),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_2),
.B(n_65),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_2),
.B(n_46),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_2),
.A2(n_33),
.B(n_48),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_8),
.B1(n_37),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_3),
.A2(n_39),
.B(n_61),
.C(n_108),
.Y(n_107)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_22),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_5),
.A2(n_7),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_5),
.A2(n_10),
.B1(n_24),
.B2(n_34),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_8),
.B1(n_24),
.B2(n_37),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_56),
.B(n_59),
.C(n_62),
.Y(n_58)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_61),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_116),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_114),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_15),
.B(n_95),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_78),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_67),
.B2(n_68),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_40),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_20),
.A2(n_29),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_21),
.B(n_26),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_23),
.A2(n_26),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_26),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_26),
.B(n_39),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_29),
.A2(n_102),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_29),
.B(n_109),
.C(n_166),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_29),
.A2(n_102),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_29),
.B(n_183),
.C(n_190),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_30),
.B(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_33),
.A2(n_34),
.B(n_39),
.C(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_70),
.B(n_71),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_35),
.B(n_39),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_39),
.A2(n_44),
.B(n_49),
.C(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_54),
.B2(n_66),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_41),
.A2(n_42),
.B1(n_123),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_41),
.A2(n_42),
.B1(n_85),
.B2(n_86),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_42),
.B(n_93),
.C(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_42),
.B(n_86),
.C(n_172),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_50),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_43),
.Y(n_113)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_47),
.B(n_48),
.C(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_47),
.A2(n_51),
.B1(n_52),
.B2(n_113),
.Y(n_112)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_105),
.C(n_111),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_66),
.B1(n_111),
.B2(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_63),
.B2(n_65),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_65),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_64),
.Y(n_94)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_76),
.B(n_82),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.C(n_93),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_85),
.B1(n_86),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_81),
.A2(n_110),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_85),
.A2(n_86),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_86),
.B(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_98),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.C(n_103),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_103),
.A2(n_104),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_158),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_134),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_112),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_136),
.C(n_138),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_141),
.B(n_198),
.C(n_204),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_128),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_118),
.B(n_128),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_120),
.B(n_122),
.C(n_126),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.C(n_135),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_135),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_148),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_197),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_192),
.B(n_196),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_180),
.B(n_191),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_169),
.B(n_179),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_161),
.B(n_168),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_153),
.B(n_160),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B(n_159),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_173),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_182),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_189),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);


endmodule