module fake_jpeg_25059_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_38),
.B1(n_40),
.B2(n_36),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_23),
.B1(n_22),
.B2(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_35),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_16),
.B1(n_32),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_19),
.B1(n_21),
.B2(n_42),
.Y(n_90)
);

AND2x4_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_17),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_35),
.B(n_29),
.C(n_34),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_63),
.Y(n_68)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_85),
.B1(n_16),
.B2(n_21),
.Y(n_117)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_54),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_84),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_87),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_83),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_40),
.B1(n_34),
.B2(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_49),
.B1(n_62),
.B2(n_50),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_31),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_43),
.B1(n_41),
.B2(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_115),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_54),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_112),
.C(n_114),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_54),
.B1(n_47),
.B2(n_50),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_98),
.B1(n_107),
.B2(n_117),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_76),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_62),
.B1(n_50),
.B2(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_108),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_71),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_55),
.C(n_56),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_27),
.C(n_20),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_70),
.B1(n_66),
.B2(n_78),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_121),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_70),
.B1(n_78),
.B2(n_77),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_83),
.B1(n_90),
.B2(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_129),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_89),
.B1(n_82),
.B2(n_88),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_133),
.B1(n_137),
.B2(n_99),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_77),
.B1(n_57),
.B2(n_60),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_134),
.B(n_80),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_67),
.B1(n_81),
.B2(n_43),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_41),
.B1(n_42),
.B2(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_138),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_107),
.B1(n_105),
.B2(n_112),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

CKINVDCx12_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_141),
.Y(n_152)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_71),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_97),
.B(n_96),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_120),
.B(n_133),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_111),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_94),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_158),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_91),
.C(n_71),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_132),
.B1(n_123),
.B2(n_99),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_15),
.C(n_13),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_167),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_172),
.C(n_143),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_119),
.B1(n_135),
.B2(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_119),
.B1(n_137),
.B2(n_124),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_175),
.C(n_181),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_126),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_143),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_192),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_132),
.B(n_27),
.C(n_18),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_144),
.B(n_156),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_127),
.B1(n_122),
.B2(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_166),
.Y(n_199)
);

CKINVDCx10_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_191),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_160),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_145),
.B(n_165),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_184),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_208),
.B1(n_214),
.B2(n_180),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_171),
.B(n_157),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_30),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_151),
.B(n_13),
.C(n_15),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_27),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_26),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_175),
.B(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_219),
.B1(n_221),
.B2(n_206),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_170),
.B1(n_177),
.B2(n_185),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_168),
.B1(n_171),
.B2(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_168),
.C(n_188),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_225),
.C(n_226),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_191),
.C(n_116),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_20),
.C(n_24),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_24),
.C(n_80),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_214),
.C(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_237),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_196),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_243),
.B1(n_213),
.B2(n_197),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_198),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_193),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_255),
.Y(n_268)
);

OAI322xp33_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_231),
.A3(n_208),
.B1(n_233),
.B2(n_227),
.C1(n_228),
.C2(n_215),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_242),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

FAx1_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_220),
.CI(n_227),
.CON(n_257),
.SN(n_257)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_0),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_204),
.B1(n_229),
.B2(n_199),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_211),
.B1(n_41),
.B2(n_16),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_240),
.C(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_265),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_205),
.B(n_241),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_205),
.B(n_213),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_270),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_30),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_18),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_9),
.B(n_12),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_257),
.B1(n_259),
.B2(n_2),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_262),
.B(n_257),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_7),
.B(n_12),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_24),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_80),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_42),
.B1(n_24),
.B2(n_18),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_269),
.C(n_271),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_287),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_6),
.B(n_12),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_11),
.B(n_10),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_6),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_273),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_285),
.B(n_7),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_273),
.A3(n_26),
.B1(n_6),
.B2(n_8),
.C1(n_11),
.C2(n_5),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

AOI222xp33_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_289),
.B1(n_290),
.B2(n_7),
.C1(n_3),
.C2(n_0),
.Y(n_295)
);

AOI321xp33_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_294),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_1),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_1),
.C(n_3),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_1),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_1),
.B(n_4),
.C(n_26),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_4),
.Y(n_300)
);


endmodule