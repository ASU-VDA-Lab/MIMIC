module fake_jpeg_14784_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_24),
.B1(n_27),
.B2(n_20),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_42),
.B1(n_21),
.B2(n_14),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_15),
.B1(n_25),
.B2(n_21),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_27),
.B(n_20),
.C(n_25),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_14),
.B(n_28),
.C(n_17),
.Y(n_63)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_24),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_36),
.Y(n_55)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_20),
.B1(n_17),
.B2(n_28),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_61),
.B1(n_19),
.B2(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_63),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_33),
.B1(n_31),
.B2(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_65),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_40),
.B(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_40),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_76),
.B1(n_85),
.B2(n_90),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_48),
.B1(n_44),
.B2(n_50),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_60),
.B(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_71),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_33),
.B1(n_31),
.B2(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_63),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_55),
.C(n_60),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_99),
.C(n_33),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_101),
.B(n_109),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_59),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_110),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_92),
.B(n_72),
.C(n_76),
.D(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_66),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_29),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_74),
.B1(n_86),
.B2(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_115),
.B1(n_123),
.B2(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_90),
.B1(n_75),
.B2(n_52),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_26),
.B(n_16),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_96),
.B1(n_111),
.B2(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_16),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_109),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_136),
.C(n_98),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_95),
.Y(n_138)
);

BUFx16f_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_142),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_119),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_103),
.B1(n_6),
.B2(n_8),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_145),
.C(n_133),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_121),
.A3(n_113),
.B1(n_123),
.B2(n_112),
.C1(n_122),
.C2(n_120),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_120),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_98),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_139),
.B1(n_141),
.B2(n_5),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_136),
.C(n_137),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_156),
.C(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_159),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_8),
.B(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_9),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_9),
.Y(n_160)
);

AOI21x1_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_146),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_143),
.C(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.C(n_162),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_155),
.C(n_10),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_164),
.B(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_170),
.B(n_12),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_12),
.C(n_13),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_175),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_8),
.Y(n_180)
);


endmodule