module fake_jpeg_24899_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_7),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_2),
.Y(n_44)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_18),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_21),
.B(n_20),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_14),
.B1(n_17),
.B2(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_42),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_23),
.B(n_12),
.C(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_54),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_15),
.B1(n_18),
.B2(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_18),
.B1(n_33),
.B2(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_44),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_73),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_41),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_61),
.B1(n_46),
.B2(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_61),
.B1(n_46),
.B2(n_36),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_68),
.B(n_72),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_12),
.B(n_66),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_57),
.B1(n_54),
.B2(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_56),
.B1(n_41),
.B2(n_14),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_81),
.B(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_56),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_3),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_49),
.B1(n_17),
.B2(n_23),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_63),
.C(n_67),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_86),
.B(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_75),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_89),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_100),
.C(n_80),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_76),
.B(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_74),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.C(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

OAI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_107),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_108),
.Y(n_111)
);


endmodule