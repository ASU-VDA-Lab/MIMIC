module fake_jpeg_22514_n_60 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_10),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_5),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_6),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_31),
.B1(n_27),
.B2(n_43),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_51),
.B1(n_14),
.B2(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_52),
.B(n_19),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_22),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_23),
.Y(n_60)
);


endmodule