module fake_jpeg_711_n_131 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_6),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_41),
.Y(n_47)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_15),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_44),
.Y(n_68)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_43),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_13),
.B(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_65),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_30),
.A2(n_22),
.B1(n_12),
.B2(n_25),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_61),
.B1(n_65),
.B2(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_25),
.B1(n_16),
.B2(n_21),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_64),
.B1(n_70),
.B2(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_46),
.B1(n_43),
.B2(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_33),
.A2(n_16),
.B1(n_21),
.B2(n_12),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_31),
.A2(n_20),
.B1(n_23),
.B2(n_15),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_70),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_2),
.B1(n_20),
.B2(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_47),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_81),
.B(n_49),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_59),
.B1(n_61),
.B2(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_56),
.C(n_50),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_86),
.C(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_64),
.C(n_58),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_98),
.C(n_87),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_77),
.B1(n_73),
.B2(n_86),
.Y(n_101)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_93),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_102),
.B1(n_92),
.B2(n_93),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_71),
.B1(n_87),
.B2(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_98),
.C(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_90),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_116),
.B(n_98),
.C(n_87),
.D(n_96),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_114),
.B1(n_90),
.B2(n_96),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_118),
.B(n_79),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_106),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_115),
.B(n_116),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_118),
.A3(n_89),
.B1(n_104),
.B2(n_95),
.C1(n_99),
.C2(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_89),
.Y(n_128)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_99),
.B(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);


endmodule