module fake_jpeg_5459_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_28),
.CON(n_52),
.SN(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_16),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_12),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_62),
.B1(n_25),
.B2(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_28),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_59),
.B(n_37),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_53),
.B(n_60),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_31),
.B(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_31),
.B1(n_26),
.B2(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_37),
.B1(n_25),
.B2(n_17),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_67),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_18),
.B(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_26),
.B1(n_27),
.B2(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_21),
.B1(n_19),
.B2(n_27),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_60),
.B1(n_62),
.B2(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_22),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_85),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_80),
.B(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_56),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_64),
.B1(n_62),
.B2(n_66),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_90),
.B1(n_61),
.B2(n_66),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_92),
.Y(n_108)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_0),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_57),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_59),
.C(n_53),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_95),
.A2(n_107),
.B(n_112),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_54),
.B(n_53),
.C(n_47),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_78),
.B(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_46),
.B1(n_54),
.B2(n_36),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_103),
.B1(n_88),
.B2(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_111),
.B1(n_115),
.B2(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_84),
.B(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_67),
.B1(n_65),
.B2(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_57),
.B1(n_49),
.B2(n_63),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_49),
.B1(n_57),
.B2(n_63),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_73),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_86),
.Y(n_137)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_71),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_121),
.B1(n_94),
.B2(n_99),
.Y(n_161)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_74),
.C(n_79),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_33),
.C(n_40),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_131),
.B1(n_103),
.B2(n_100),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_85),
.B1(n_79),
.B2(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_1),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_134),
.B(n_117),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_104),
.B1(n_106),
.B2(n_96),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_85),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_144),
.B(n_145),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_98),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_58),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_165),
.B(n_130),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_155),
.B1(n_120),
.B2(n_139),
.Y(n_173)
);

NAND2x1_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_111),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_159),
.B(n_161),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_105),
.B1(n_112),
.B2(n_119),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_119),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_162),
.C(n_163),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_94),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_167),
.Y(n_188)
);

OAI22x1_ASAP7_75t_R g159 ( 
.A1(n_128),
.A2(n_109),
.B1(n_40),
.B2(n_33),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_58),
.C(n_33),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_136),
.B(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_58),
.C(n_40),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_172),
.C(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_72),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_126),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_58),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_181),
.B1(n_187),
.B2(n_196),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_179),
.C(n_186),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_198),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_185),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_134),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_184),
.B(n_193),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_139),
.B1(n_166),
.B2(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_133),
.B(n_131),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_127),
.C(n_143),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_170),
.B(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_127),
.C(n_132),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.C(n_172),
.Y(n_202)
);

NAND2x1p5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_140),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_123),
.B(n_18),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_170),
.B1(n_150),
.B2(n_158),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_123),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_125),
.B1(n_122),
.B2(n_76),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_18),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_205),
.C(n_214),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_209),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_164),
.C(n_161),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_168),
.B1(n_151),
.B2(n_157),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_217),
.B1(n_187),
.B2(n_178),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_164),
.C(n_165),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_148),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_198),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_174),
.B(n_165),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_181),
.Y(n_231)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_150),
.C(n_169),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_202),
.C(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_183),
.B1(n_194),
.B2(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_24),
.B1(n_17),
.B2(n_3),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_227),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_201),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_219),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_180),
.B1(n_192),
.B2(n_188),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_182),
.C(n_101),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_118),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_77),
.C(n_92),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_241),
.C(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_213),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_92),
.C(n_25),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_25),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_242),
.Y(n_248)
);

AO221x1_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_256),
.B1(n_255),
.B2(n_246),
.C(n_258),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_212),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_259),
.C(n_260),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_209),
.B1(n_200),
.B2(n_216),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_231),
.A3(n_223),
.B1(n_237),
.B2(n_232),
.C1(n_241),
.C2(n_236),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_204),
.C(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_257),
.C(n_261),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_216),
.Y(n_256)
);

XOR2x1_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_252),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_222),
.C(n_200),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_243),
.B(n_15),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_24),
.C(n_17),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_262),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_271),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_269),
.CI(n_263),
.CON(n_285),
.SN(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_229),
.C(n_15),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_251),
.C(n_247),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_24),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_14),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_247),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_14),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_4),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_1),
.C(n_3),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_284),
.C(n_287),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_3),
.C(n_4),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_4),
.C(n_5),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_271),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_295),
.B(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_264),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

AOI222xp33_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_267),
.B1(n_270),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_299),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_11),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_10),
.C2(n_4),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_284),
.Y(n_304)
);

AOI31xp33_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_6),
.A3(n_7),
.B(n_10),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_302),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_288),
.B(n_287),
.C(n_280),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_10),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_6),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.C(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_10),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_302),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_307),
.Y(n_317)
);


endmodule