module real_aes_7001_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g168 ( .A1(n_0), .A2(n_169), .B(n_172), .C(n_176), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_1), .B(n_160), .Y(n_179) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_2), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g445 ( .A(n_2), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_3), .B(n_170), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_4), .A2(n_133), .B(n_136), .C(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_5), .A2(n_128), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_6), .A2(n_128), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_7), .B(n_160), .Y(n_549) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_8), .A2(n_162), .B(n_234), .Y(n_233) );
AND2x6_ASAP7_75t_L g133 ( .A(n_9), .B(n_134), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_10), .A2(n_133), .B(n_136), .C(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g509 ( .A(n_11), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_12), .B(n_40), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_12), .B(n_40), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_13), .B(n_175), .Y(n_520) );
INVx1_ASAP7_75t_L g154 ( .A(n_14), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_15), .B(n_170), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_16), .A2(n_171), .B(n_529), .C(n_531), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_17), .B(n_160), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_18), .B(n_148), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_19), .A2(n_136), .B(n_139), .C(n_147), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_20), .A2(n_174), .B(n_242), .C(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_21), .B(n_175), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_22), .A2(n_75), .B1(n_452), .B2(n_740), .C1(n_743), .C2(n_744), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_23), .B(n_175), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_24), .Y(n_490) );
INVx1_ASAP7_75t_L g470 ( .A(n_25), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_26), .A2(n_136), .B(n_147), .C(n_237), .Y(n_236) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_27), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_28), .Y(n_516) );
INVx1_ASAP7_75t_L g484 ( .A(n_29), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_30), .A2(n_128), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g131 ( .A(n_31), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_32), .A2(n_186), .B(n_187), .C(n_191), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_33), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_34), .A2(n_174), .B(n_546), .C(n_548), .Y(n_545) );
INVxp67_ASAP7_75t_L g485 ( .A(n_35), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_36), .A2(n_100), .B1(n_109), .B2(n_748), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_37), .B(n_239), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_38), .A2(n_136), .B(n_147), .C(n_469), .Y(n_468) );
CKINVDCx14_ASAP7_75t_R g544 ( .A(n_39), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_41), .A2(n_176), .B(n_507), .C(n_508), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_42), .B(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_43), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_44), .B(n_170), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_45), .B(n_128), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_46), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_47), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_48), .B(n_448), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_49), .A2(n_186), .B(n_191), .C(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g173 ( .A(n_50), .Y(n_173) );
INVx1_ASAP7_75t_L g217 ( .A(n_51), .Y(n_217) );
INVx1_ASAP7_75t_L g557 ( .A(n_52), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_53), .B(n_128), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_54), .Y(n_156) );
CKINVDCx14_ASAP7_75t_R g505 ( .A(n_55), .Y(n_505) );
INVx1_ASAP7_75t_L g134 ( .A(n_56), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_57), .B(n_128), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_58), .B(n_160), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_59), .A2(n_146), .B(n_202), .C(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
INVx1_ASAP7_75t_SL g547 ( .A(n_61), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_62), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_63), .B(n_170), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_64), .B(n_160), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_65), .B(n_171), .Y(n_252) );
INVx1_ASAP7_75t_L g493 ( .A(n_66), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g166 ( .A(n_67), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_68), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_69), .A2(n_136), .B(n_191), .C(n_200), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_70), .Y(n_226) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_72), .A2(n_128), .B(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_73), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_74), .A2(n_128), .B(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_75), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_76), .A2(n_127), .B(n_480), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_77), .Y(n_467) );
INVx1_ASAP7_75t_L g527 ( .A(n_78), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_79), .B(n_144), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_80), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_81), .A2(n_128), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g530 ( .A(n_82), .Y(n_530) );
INVx2_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
INVx1_ASAP7_75t_L g519 ( .A(n_84), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_85), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_86), .B(n_175), .Y(n_253) );
INVx2_ASAP7_75t_L g105 ( .A(n_87), .Y(n_105) );
OR2x2_ASAP7_75t_L g442 ( .A(n_87), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g455 ( .A(n_87), .B(n_444), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_88), .A2(n_136), .B(n_191), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_89), .B(n_128), .Y(n_184) );
INVx1_ASAP7_75t_L g188 ( .A(n_90), .Y(n_188) );
INVxp67_ASAP7_75t_L g229 ( .A(n_91), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_92), .A2(n_116), .B1(n_438), .B2(n_439), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_92), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_93), .B(n_162), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_94), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g201 ( .A(n_95), .Y(n_201) );
INVx1_ASAP7_75t_L g248 ( .A(n_96), .Y(n_248) );
INVx2_ASAP7_75t_L g560 ( .A(n_97), .Y(n_560) );
AND2x2_ASAP7_75t_L g219 ( .A(n_98), .B(n_150), .Y(n_219) );
INVx2_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g749 ( .A(n_101), .Y(n_749) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
OR2x2_ASAP7_75t_L g459 ( .A(n_105), .B(n_444), .Y(n_459) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_105), .B(n_443), .Y(n_746) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_450), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g747 ( .A(n_111), .Y(n_747) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI21xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_440), .B(n_447), .Y(n_114) );
INVx1_ASAP7_75t_L g439 ( .A(n_116), .Y(n_439) );
INVx2_ASAP7_75t_L g456 ( .A(n_116), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_116), .A2(n_453), .B1(n_741), .B2(n_742), .Y(n_740) );
AND2x2_ASAP7_75t_SL g116 ( .A(n_117), .B(n_393), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_328), .Y(n_117) );
NAND4xp25_ASAP7_75t_SL g118 ( .A(n_119), .B(n_273), .C(n_297), .D(n_320), .Y(n_118) );
AOI221xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_210), .B1(n_244), .B2(n_257), .C(n_260), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_180), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_122), .A2(n_158), .B1(n_211), .B2(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_122), .B(n_181), .Y(n_331) );
AND2x2_ASAP7_75t_L g350 ( .A(n_122), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_122), .B(n_334), .Y(n_420) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_158), .Y(n_122) );
AND2x2_ASAP7_75t_L g288 ( .A(n_123), .B(n_181), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_123), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g311 ( .A(n_123), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_123), .B(n_159), .Y(n_316) );
INVx2_ASAP7_75t_L g348 ( .A(n_123), .Y(n_348) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_123), .Y(n_392) );
AND2x2_ASAP7_75t_L g409 ( .A(n_123), .B(n_286), .Y(n_409) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g327 ( .A(n_124), .B(n_286), .Y(n_327) );
AND2x4_ASAP7_75t_L g341 ( .A(n_124), .B(n_158), .Y(n_341) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_124), .Y(n_345) );
AND2x2_ASAP7_75t_L g365 ( .A(n_124), .B(n_280), .Y(n_365) );
AND2x2_ASAP7_75t_L g415 ( .A(n_124), .B(n_182), .Y(n_415) );
AND2x2_ASAP7_75t_L g425 ( .A(n_124), .B(n_159), .Y(n_425) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_155), .Y(n_124) );
AOI21xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_135), .B(n_148), .Y(n_125) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g249 ( .A(n_129), .B(n_133), .Y(n_249) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g146 ( .A(n_130), .Y(n_146) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g243 ( .A(n_131), .Y(n_243) );
INVx1_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
INVx3_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
INVx1_ASAP7_75t_L g239 ( .A(n_132), .Y(n_239) );
BUFx3_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
INVx4_ASAP7_75t_SL g178 ( .A(n_133), .Y(n_178) );
INVx5_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx3_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_145), .Y(n_139) );
INVx2_ASAP7_75t_L g144 ( .A(n_141), .Y(n_144) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_144), .A2(n_188), .B(n_189), .C(n_190), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_144), .A2(n_190), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_144), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_L g518 ( .A1(n_144), .A2(n_495), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_145), .A2(n_170), .B(n_470), .C(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_146), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_149), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_150), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_150), .A2(n_214), .B(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_150), .A2(n_249), .B(n_467), .C(n_468), .Y(n_466) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_150), .A2(n_503), .B(n_510), .Y(n_502) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_L g163 ( .A(n_151), .B(n_152), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_157), .A2(n_515), .B(n_521), .Y(n_514) );
AND2x2_ASAP7_75t_L g281 ( .A(n_158), .B(n_181), .Y(n_281) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_158), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_158), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g371 ( .A(n_158), .Y(n_371) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g259 ( .A(n_159), .B(n_196), .Y(n_259) );
AND2x2_ASAP7_75t_L g286 ( .A(n_159), .B(n_197), .Y(n_286) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_164), .B(n_179), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_161), .B(n_193), .Y(n_192) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_161), .A2(n_198), .B(n_208), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_161), .B(n_209), .Y(n_208) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_161), .A2(n_247), .B(n_254), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_161), .B(n_473), .Y(n_472) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_161), .A2(n_489), .B(n_496), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_161), .B(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_162), .A2(n_235), .B(n_236), .Y(n_234) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g256 ( .A(n_163), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_178), .Y(n_165) );
INVx2_ASAP7_75t_L g186 ( .A(n_167), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_167), .A2(n_178), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_167), .A2(n_178), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_167), .A2(n_178), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g526 ( .A1(n_167), .A2(n_178), .B(n_527), .C(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_167), .A2(n_178), .B(n_544), .C(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_SL g556 ( .A1(n_167), .A2(n_178), .B(n_557), .C(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_170), .B(n_229), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_170), .A2(n_203), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_171), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_174), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g507 ( .A(n_175), .Y(n_507) );
INVx2_ASAP7_75t_L g495 ( .A(n_176), .Y(n_495) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_177), .Y(n_190) );
INVx1_ASAP7_75t_L g531 ( .A(n_177), .Y(n_531) );
INVx1_ASAP7_75t_L g191 ( .A(n_178), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_180), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_194), .Y(n_180) );
OR2x2_ASAP7_75t_L g312 ( .A(n_181), .B(n_195), .Y(n_312) );
AND2x2_ASAP7_75t_L g349 ( .A(n_181), .B(n_259), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_181), .B(n_280), .Y(n_360) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_181), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_181), .B(n_316), .Y(n_433) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx2_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
AND2x2_ASAP7_75t_L g267 ( .A(n_182), .B(n_195), .Y(n_267) );
AND2x2_ASAP7_75t_L g383 ( .A(n_182), .B(n_278), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_182), .B(n_316), .Y(n_405) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_192), .Y(n_182) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_195), .Y(n_351) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_196), .Y(n_303) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_207), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_204), .C(n_205), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_203), .B(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_203), .B(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g548 ( .A(n_206), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_220), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_211), .B(n_293), .Y(n_412) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_212), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g264 ( .A(n_212), .B(n_265), .Y(n_264) );
INVx5_ASAP7_75t_SL g272 ( .A(n_212), .Y(n_272) );
OR2x2_ASAP7_75t_L g295 ( .A(n_212), .B(n_265), .Y(n_295) );
OR2x2_ASAP7_75t_L g305 ( .A(n_212), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g368 ( .A(n_212), .B(n_222), .Y(n_368) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_212), .B(n_221), .Y(n_406) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_212), .B(n_348), .C(n_428), .D(n_429), .Y(n_427) );
AND2x2_ASAP7_75t_L g437 ( .A(n_212), .B(n_269), .Y(n_437) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_219), .Y(n_212) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g262 ( .A(n_221), .B(n_258), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_221), .B(n_264), .Y(n_431) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_231), .Y(n_221) );
OR2x2_ASAP7_75t_L g271 ( .A(n_222), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_222), .B(n_246), .Y(n_290) );
INVxp67_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_222), .B(n_265), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_222), .B(n_232), .Y(n_359) );
AND2x2_ASAP7_75t_L g374 ( .A(n_222), .B(n_269), .Y(n_374) );
OR2x2_ASAP7_75t_L g403 ( .A(n_222), .B(n_232), .Y(n_403) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_230), .Y(n_222) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_223), .A2(n_525), .B(n_532), .Y(n_524) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_223), .A2(n_542), .B(n_549), .Y(n_541) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_223), .A2(n_555), .B(n_561), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_231), .B(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_231), .B(n_272), .Y(n_411) );
OR2x2_ASAP7_75t_L g432 ( .A(n_231), .B(n_309), .Y(n_432) );
INVx1_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g245 ( .A(n_232), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g269 ( .A(n_232), .B(n_265), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_232), .B(n_246), .Y(n_284) );
AND2x2_ASAP7_75t_L g354 ( .A(n_232), .B(n_278), .Y(n_354) );
AND2x2_ASAP7_75t_L g388 ( .A(n_232), .B(n_272), .Y(n_388) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_233), .B(n_272), .Y(n_291) );
AND2x2_ASAP7_75t_L g319 ( .A(n_233), .B(n_246), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B(n_241), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_241), .A2(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_244), .B(n_327), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_245), .A2(n_334), .B1(n_370), .B2(n_387), .C(n_389), .Y(n_386) );
INVx5_ASAP7_75t_SL g265 ( .A(n_246), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_250), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_249), .A2(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_249), .A2(n_516), .B(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g478 ( .A(n_256), .Y(n_478) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OAI33xp33_ASAP7_75t_L g285 ( .A1(n_258), .A2(n_286), .A3(n_287), .B1(n_289), .B2(n_292), .B3(n_296), .Y(n_285) );
OR2x2_ASAP7_75t_L g301 ( .A(n_258), .B(n_302), .Y(n_301) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_258), .A2(n_327), .A3(n_334), .B1(n_411), .B2(n_412), .C1(n_413), .C2(n_416), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_258), .B(n_286), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_SL g434 ( .A1(n_258), .A2(n_286), .B(n_435), .C(n_437), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_259), .A2(n_274), .B1(n_279), .B2(n_282), .C(n_285), .Y(n_273) );
INVx1_ASAP7_75t_L g366 ( .A(n_259), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_259), .B(n_415), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B1(n_266), .B2(n_268), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g343 ( .A(n_264), .B(n_278), .Y(n_343) );
AND2x2_ASAP7_75t_L g401 ( .A(n_264), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_272), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_265), .B(n_278), .Y(n_337) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_267), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_267), .B(n_345), .Y(n_399) );
OAI321xp33_ASAP7_75t_L g418 ( .A1(n_267), .A2(n_340), .A3(n_419), .B1(n_420), .B2(n_421), .C(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g385 ( .A(n_268), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g324 ( .A(n_269), .B(n_272), .Y(n_324) );
AOI321xp33_ASAP7_75t_L g382 ( .A1(n_269), .A2(n_286), .A3(n_383), .B1(n_384), .B2(n_385), .C(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_284), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_272), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_272), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_272), .B(n_358), .Y(n_395) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g318 ( .A(n_276), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g283 ( .A(n_277), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g391 ( .A(n_278), .Y(n_391) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_281), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g314 ( .A(n_286), .Y(n_314) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_288), .B(n_323), .Y(n_372) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g336 ( .A(n_291), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g381 ( .A(n_291), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_292), .A2(n_339), .B1(n_342), .B2(n_344), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g436 ( .A(n_295), .B(n_359), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_300), .B1(n_304), .B2(n_310), .C(n_313), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_SL g380 ( .A(n_306), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_308), .B(n_358), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_308), .A2(n_376), .B(n_378), .Y(n_375) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g421 ( .A(n_309), .B(n_403), .Y(n_421) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g323 ( .A(n_312), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_368), .Y(n_367) );
INVxp67_ASAP7_75t_L g429 ( .A(n_319), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .B(n_325), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_323), .B(n_341), .Y(n_377) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g398 ( .A(n_327), .Y(n_398) );
NAND5xp2_ASAP7_75t_L g328 ( .A(n_329), .B(n_346), .C(n_355), .D(n_375), .E(n_382), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_335), .C(n_338), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_342), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_350), .B(n_352), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_347), .A2(n_401), .B1(n_404), .B2(n_406), .C(n_407), .Y(n_400) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AOI321xp33_ASAP7_75t_L g355 ( .A1(n_348), .A2(n_356), .A3(n_360), .B1(n_361), .B2(n_367), .C(n_369), .Y(n_355) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g426 ( .A(n_360), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_366), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g378 ( .A(n_363), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NOR2xp67_ASAP7_75t_SL g390 ( .A(n_364), .B(n_371), .Y(n_390) );
AOI321xp33_ASAP7_75t_SL g422 ( .A1(n_367), .A2(n_423), .A3(n_424), .B1(n_425), .B2(n_426), .C(n_427), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_372), .C(n_373), .Y(n_369) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_380), .B(n_388), .Y(n_417) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .C(n_392), .Y(n_389) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_418), .C(n_430), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_396), .B(n_400), .C(n_410), .Y(n_394) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_399), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_431), .B1(n_432), .B2(n_433), .C(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g419 ( .A(n_401), .Y(n_419) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g423 ( .A(n_421), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_442), .Y(n_449) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_447), .A2(n_451), .B(n_747), .Y(n_450) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .B1(n_457), .B2(n_460), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g742 ( .A(n_458), .Y(n_742) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g741 ( .A(n_460), .Y(n_741) );
OR4x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_630), .C(n_677), .D(n_717), .Y(n_460) );
NAND3xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_576), .C(n_605), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_498), .B(n_533), .C(n_569), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_463), .A2(n_589), .B(n_606), .C(n_610), .Y(n_605) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_474), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_465), .B(n_568), .Y(n_567) );
INVx3_ASAP7_75t_SL g572 ( .A(n_465), .Y(n_572) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_465), .Y(n_584) );
AND2x4_ASAP7_75t_L g588 ( .A(n_465), .B(n_540), .Y(n_588) );
AND2x2_ASAP7_75t_L g599 ( .A(n_465), .B(n_488), .Y(n_599) );
OR2x2_ASAP7_75t_L g623 ( .A(n_465), .B(n_536), .Y(n_623) );
AND2x2_ASAP7_75t_L g636 ( .A(n_465), .B(n_541), .Y(n_636) );
AND2x2_ASAP7_75t_L g676 ( .A(n_465), .B(n_662), .Y(n_676) );
AND2x2_ASAP7_75t_L g683 ( .A(n_465), .B(n_646), .Y(n_683) );
AND2x2_ASAP7_75t_L g713 ( .A(n_465), .B(n_475), .Y(n_713) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_474), .B(n_640), .Y(n_652) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_487), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_475), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g590 ( .A(n_475), .B(n_487), .Y(n_590) );
BUFx3_ASAP7_75t_L g598 ( .A(n_475), .Y(n_598) );
OR2x2_ASAP7_75t_L g619 ( .A(n_475), .B(n_501), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_475), .B(n_640), .Y(n_730) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_486), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_477), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g537 ( .A(n_479), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_486), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_487), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g583 ( .A(n_487), .Y(n_583) );
AND2x2_ASAP7_75t_L g646 ( .A(n_487), .B(n_541), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_487), .A2(n_649), .B1(n_651), .B2(n_653), .C(n_654), .Y(n_648) );
AND2x2_ASAP7_75t_L g662 ( .A(n_487), .B(n_536), .Y(n_662) );
AND2x2_ASAP7_75t_L g688 ( .A(n_487), .B(n_572), .Y(n_688) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g568 ( .A(n_488), .B(n_541), .Y(n_568) );
BUFx2_ASAP7_75t_L g702 ( .A(n_488), .Y(n_702) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI32xp33_ASAP7_75t_L g668 ( .A1(n_499), .A2(n_629), .A3(n_643), .B1(n_669), .B2(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
AND2x2_ASAP7_75t_L g609 ( .A(n_500), .B(n_553), .Y(n_609) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g591 ( .A(n_501), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_501), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g663 ( .A(n_501), .B(n_553), .Y(n_663) );
AND2x2_ASAP7_75t_L g674 ( .A(n_501), .B(n_566), .Y(n_674) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g575 ( .A(n_502), .B(n_554), .Y(n_575) );
AND2x2_ASAP7_75t_L g579 ( .A(n_502), .B(n_554), .Y(n_579) );
AND2x2_ASAP7_75t_L g614 ( .A(n_502), .B(n_565), .Y(n_614) );
AND2x2_ASAP7_75t_L g621 ( .A(n_502), .B(n_523), .Y(n_621) );
OAI211xp5_ASAP7_75t_L g626 ( .A1(n_502), .A2(n_572), .B(n_583), .C(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g680 ( .A(n_502), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_502), .B(n_513), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_511), .B(n_563), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_511), .B(n_579), .Y(n_669) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g574 ( .A(n_512), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_523), .Y(n_512) );
AND2x2_ASAP7_75t_L g566 ( .A(n_513), .B(n_524), .Y(n_566) );
OR2x2_ASAP7_75t_L g581 ( .A(n_513), .B(n_524), .Y(n_581) );
AND2x2_ASAP7_75t_L g604 ( .A(n_513), .B(n_565), .Y(n_604) );
INVx1_ASAP7_75t_L g608 ( .A(n_513), .Y(n_608) );
AND2x2_ASAP7_75t_L g627 ( .A(n_513), .B(n_564), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_513), .A2(n_592), .B1(n_638), .B2(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_513), .B(n_680), .Y(n_704) );
AND2x2_ASAP7_75t_L g719 ( .A(n_513), .B(n_579), .Y(n_719) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
AND2x2_ASAP7_75t_L g593 ( .A(n_514), .B(n_524), .Y(n_593) );
AND2x2_ASAP7_75t_L g595 ( .A(n_514), .B(n_553), .Y(n_595) );
AND3x2_ASAP7_75t_L g657 ( .A(n_514), .B(n_621), .C(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g692 ( .A(n_523), .B(n_564), .Y(n_692) );
INVx1_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g553 ( .A(n_524), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_524), .B(n_563), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_524), .B(n_604), .C(n_680), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_550), .B1(n_562), .B2(n_567), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_536), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g644 ( .A(n_536), .Y(n_644) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_539), .A2(n_661), .A3(n_662), .B(n_663), .Y(n_660) );
AND2x2_ASAP7_75t_L g685 ( .A(n_539), .B(n_572), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_539), .B(n_598), .Y(n_731) );
AND2x2_ASAP7_75t_L g640 ( .A(n_540), .B(n_572), .Y(n_640) );
AND2x2_ASAP7_75t_L g701 ( .A(n_540), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g571 ( .A(n_541), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g629 ( .A(n_541), .Y(n_629) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g650 ( .A(n_551), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_552), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AOI221x1_ASAP7_75t_SL g617 ( .A1(n_553), .A2(n_618), .B1(n_620), .B2(n_622), .C(n_624), .Y(n_617) );
INVx2_ASAP7_75t_L g565 ( .A(n_554), .Y(n_565) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_554), .Y(n_659) );
INVx1_ASAP7_75t_L g647 ( .A(n_562), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_563), .B(n_580), .Y(n_672) );
INVx1_ASAP7_75t_SL g735 ( .A(n_563), .Y(n_735) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g653 ( .A(n_566), .B(n_579), .Y(n_653) );
INVx1_ASAP7_75t_L g721 ( .A(n_567), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_567), .B(n_650), .Y(n_734) );
INVx2_ASAP7_75t_SL g573 ( .A(n_568), .Y(n_573) );
AND2x2_ASAP7_75t_L g616 ( .A(n_568), .B(n_572), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_568), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_568), .B(n_643), .Y(n_670) );
AOI21xp33_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_573), .B(n_574), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_571), .B(n_643), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_571), .B(n_598), .Y(n_739) );
OR2x2_ASAP7_75t_L g611 ( .A(n_572), .B(n_590), .Y(n_611) );
AND2x2_ASAP7_75t_L g710 ( .A(n_572), .B(n_701), .Y(n_710) );
OAI22xp5_ASAP7_75t_SL g585 ( .A1(n_573), .A2(n_586), .B1(n_591), .B2(n_594), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_573), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g633 ( .A(n_575), .B(n_581), .Y(n_633) );
INVx1_ASAP7_75t_L g697 ( .A(n_575), .Y(n_697) );
AOI311xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_582), .A3(n_584), .B(n_585), .C(n_596), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_580), .A2(n_712), .B1(n_724), .B2(n_727), .C(n_729), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_580), .B(n_735), .Y(n_737) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g634 ( .A(n_582), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g624 ( .A1(n_583), .A2(n_625), .B(n_626), .C(n_628), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_SL g693 ( .A1(n_587), .A2(n_589), .B(n_694), .C(n_695), .Y(n_693) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_588), .B(n_662), .Y(n_728) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_591), .A2(n_611), .B1(n_612), .B2(n_615), .C(n_617), .Y(n_610) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g613 ( .A(n_593), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g696 ( .A(n_593), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_597), .A2(n_655), .B(n_656), .C(n_660), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_598), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_598), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g620 ( .A(n_604), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_608), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g722 ( .A(n_611), .Y(n_722) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_614), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g649 ( .A(n_614), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g726 ( .A(n_614), .Y(n_726) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g667 ( .A(n_616), .B(n_643), .Y(n_667) );
INVx1_ASAP7_75t_SL g661 ( .A(n_623), .Y(n_661) );
INVx1_ASAP7_75t_L g638 ( .A(n_629), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_631), .B(n_648), .C(n_664), .Y(n_630) );
AOI322xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .A3(n_635), .B1(n_637), .B2(n_641), .C1(n_645), .C2(n_647), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_632), .A2(n_685), .B(n_686), .C(n_693), .Y(n_684) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_635), .A2(n_656), .B1(n_687), .B2(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g645 ( .A(n_643), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g682 ( .A(n_643), .B(n_683), .Y(n_682) );
AOI32xp33_ASAP7_75t_L g733 ( .A1(n_643), .A2(n_734), .A3(n_735), .B1(n_736), .B2(n_738), .Y(n_733) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g655 ( .A(n_646), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_646), .A2(n_699), .B1(n_703), .B2(n_705), .C(n_708), .Y(n_698) );
AND2x2_ASAP7_75t_L g712 ( .A(n_646), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g715 ( .A(n_650), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g725 ( .A(n_650), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g716 ( .A(n_659), .B(n_680), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_668), .C(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_681), .B(n_684), .C(n_698), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_692), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g707 ( .A(n_704), .Y(n_707) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B(n_714), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI211xp5_ASAP7_75t_SL g717 ( .A1(n_718), .A2(n_720), .B(n_723), .C(n_733), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule