module real_jpeg_33783_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_0),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_1),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_143),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_1),
.A2(n_143),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_3),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_5),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_5),
.A2(n_134),
.B1(n_218),
.B2(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_5),
.A2(n_134),
.B1(n_371),
.B2(n_375),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_5),
.A2(n_134),
.B1(n_417),
.B2(n_422),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_6),
.A2(n_146),
.B1(n_147),
.B2(n_153),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_6),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_6),
.A2(n_146),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_6),
.A2(n_146),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_6),
.A2(n_146),
.B1(n_259),
.B2(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_8),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_8),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_8),
.A2(n_175),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_8),
.A2(n_140),
.B1(n_175),
.B2(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_8),
.A2(n_175),
.B1(n_394),
.B2(n_397),
.Y(n_393)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_9),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_56),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_10),
.A2(n_56),
.B1(n_225),
.B2(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_10),
.A2(n_56),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_11),
.A2(n_71),
.B1(n_247),
.B2(n_252),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_13),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_14),
.A2(n_119),
.B(n_124),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_14),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_14),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_14),
.B(n_182),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_14),
.A2(n_75),
.B1(n_416),
.B2(n_433),
.Y(n_432)
);

OAI32xp33_ASAP7_75t_L g454 ( 
.A1(n_14),
.A2(n_157),
.A3(n_345),
.B1(n_455),
.B2(n_456),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_14),
.A2(n_153),
.B1(n_280),
.B2(n_315),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_15),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_16),
.A2(n_35),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_17),
.A2(n_259),
.B1(n_262),
.B2(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_17),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_287),
.Y(n_18)
);

OAI21xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_239),
.B(n_285),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_20),
.B(n_239),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_91),
.C(n_184),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_22),
.B(n_92),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_23),
.B(n_67),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B1(n_47),
.B2(n_57),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_24),
.A2(n_47),
.B1(n_57),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_24),
.A2(n_57),
.B1(n_139),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_24),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_24),
.A2(n_57),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_24),
.B(n_315),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_25),
.Y(n_245)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AO21x2_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_58),
.B(n_63),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_26)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_27),
.Y(n_263)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_28),
.Y(n_309)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_29),
.Y(n_236)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_34),
.A2(n_57),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B(n_41),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_38),
.Y(n_368)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_42),
.Y(n_142)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_46),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_46),
.Y(n_332)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_46),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_50),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_54),
.Y(n_409)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_55),
.Y(n_254)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_57),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_62),
.Y(n_251)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_62),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_63),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_75),
.B1(n_81),
.B2(n_88),
.Y(n_67)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_68),
.Y(n_228)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_69),
.Y(n_381)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_70),
.Y(n_237)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_70),
.Y(n_421)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_75),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_75),
.A2(n_81),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_75),
.A2(n_393),
.B1(n_399),
.B2(n_401),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_75),
.A2(n_416),
.B1(n_425),
.B2(n_429),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_78),
.Y(n_341)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_80),
.Y(n_261)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_80),
.Y(n_312)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_80),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_80),
.Y(n_398)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_80),
.Y(n_424)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_89),
.Y(n_313)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_90),
.Y(n_343)
);

INVx8_ASAP7_75t_L g429 ( 
.A(n_90),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_137),
.C(n_144),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_94),
.B(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_118),
.B1(n_129),
.B2(n_130),
.Y(n_94)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_95),
.A2(n_129),
.B1(n_203),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_95),
.A2(n_129),
.B1(n_203),
.B2(n_269),
.Y(n_282)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_101),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_101),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_101),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_103),
.Y(n_217)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

AOI22x1_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_113),
.Y(n_352)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_124),
.A2(n_213),
.B(n_221),
.Y(n_212)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_129),
.B(n_315),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_130),
.Y(n_199)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_144),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_156),
.B1(n_174),
.B2(n_181),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_145),
.A2(n_156),
.B1(n_181),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_152),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_174),
.B1(n_189),
.B2(n_195),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_156),
.A2(n_189),
.B1(n_195),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_156),
.A2(n_195),
.B1(n_300),
.B2(n_459),
.Y(n_458)
);

AO21x2_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_162),
.B(n_167),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g344 ( 
.A1(n_157),
.A2(n_345),
.B(n_351),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_184),
.B(n_291),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_211),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_196),
.B(n_210),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_187),
.B(n_211),
.C(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_198),
.Y(n_210)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_192),
.Y(n_280)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_193),
.Y(n_225)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

AOI22x1_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_226),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_212),
.A2(n_226),
.B1(n_227),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_222),
.C(n_224),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_234),
.B2(n_238),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_230),
.B(n_315),
.Y(n_436)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_232),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_233),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_234),
.A2(n_238),
.B1(n_307),
.B2(n_313),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_238),
.A2(n_307),
.B1(n_337),
.B2(n_342),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_238),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_283),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_265),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_255),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_245),
.A2(n_329),
.B1(n_369),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_254),
.Y(n_365)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_260),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_262),
.Y(n_437)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_277),
.B1(n_278),
.B2(n_281),
.Y(n_267)
);

INVx11_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_316),
.B(n_472),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_290),
.B(n_292),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.C(n_298),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_298),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.C(n_314),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_306),
.B1(n_314),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_346),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_352),
.C(n_353),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_SL g363 ( 
.A1(n_315),
.A2(n_364),
.B(n_366),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_356),
.B(n_471),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_320),
.B(n_322),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.C(n_333),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_323),
.A2(n_324),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_327),
.A2(n_333),
.B1(n_334),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_327),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_335),
.A2(n_336),
.B1(n_344),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_352),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

OAI21x1_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_463),
.B(n_470),
.Y(n_356)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_449),
.B(n_462),
.Y(n_357)
);

OAI21x1_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_412),
.B(n_448),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_391),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_360),
.B(n_391),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_378),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_361),
.A2(n_362),
.B1(n_378),
.B2(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_369),
.B1(n_370),
.B2(n_377),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_386),
.B1(n_387),
.B2(n_390),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_402),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_404),
.C(n_410),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_398),
.Y(n_428)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_410),
.B2(n_411),
.Y(n_402)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_403),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_439),
.B(n_447),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_431),
.B(n_438),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_430),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_415),
.B(n_430),
.Y(n_438)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_446),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_446),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_451),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_460),
.C(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_468),
.Y(n_470)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);


endmodule