module fake_aes_2680_n_41 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_16;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g14 ( .A(n_3), .B(n_0), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_9), .B(n_5), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_1), .B(n_6), .Y(n_18) );
OA21x2_ASAP7_75t_L g19 ( .A1(n_10), .A2(n_8), .B(n_4), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_1), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_14), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_20), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_17), .B(n_19), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx5_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
NAND2x1p5_ASAP7_75t_L g30 ( .A(n_29), .B(n_22), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_25), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g32 ( .A(n_31), .B(n_28), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_24), .Y(n_33) );
NAND3xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_18), .C(n_16), .Y(n_34) );
AOI221xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_21), .B1(n_30), .B2(n_14), .C(n_16), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_34), .B(n_2), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
HB1xp67_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
OAI22xp5_ASAP7_75t_SL g40 ( .A1(n_38), .A2(n_11), .B1(n_13), .B2(n_26), .Y(n_40) );
AOI22x1_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_39), .B1(n_15), .B2(n_26), .Y(n_41) );
endmodule