module fake_jpeg_31312_n_330 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_330);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_21),
.Y(n_46)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_51),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_26),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_9),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_24),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_66),
.Y(n_95)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_38),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_41),
.B1(n_37),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_84),
.B1(n_97),
.B2(n_38),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_39),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_8),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_55),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_37),
.B(n_41),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_101),
.B(n_109),
.C(n_27),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_37),
.B1(n_29),
.B2(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_85),
.B(n_96),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_94),
.B1(n_108),
.B2(n_68),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_25),
.B1(n_40),
.B2(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_42),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_25),
.B1(n_40),
.B2(n_27),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_31),
.B(n_28),
.C(n_23),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_31),
.B(n_28),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_47),
.A2(n_25),
.B1(n_39),
.B2(n_36),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_30),
.B1(n_61),
.B2(n_55),
.Y(n_113)
);

CKINVDCx9p33_ASAP7_75t_R g107 ( 
.A(n_45),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_107),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_42),
.B1(n_36),
.B2(n_32),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_54),
.B(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_38),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_122),
.B1(n_87),
.B2(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_127),
.B1(n_138),
.B2(n_72),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_30),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_118),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_61),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_52),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_125),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_52),
.B1(n_49),
.B2(n_69),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_78),
.B(n_73),
.C(n_109),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_124),
.B(n_14),
.C(n_1),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_12),
.B(n_1),
.C(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_49),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_53),
.C(n_38),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_38),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_0),
.B(n_104),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_11),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_0),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_91),
.Y(n_155)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_7),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_97),
.B1(n_111),
.B2(n_92),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_154),
.B1(n_158),
.B2(n_139),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_111),
.B1(n_92),
.B2(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_76),
.B1(n_90),
.B2(n_110),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_144),
.B(n_3),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_170),
.B1(n_129),
.B2(n_148),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_178),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_87),
.B1(n_110),
.B2(n_72),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_134),
.B(n_124),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_72),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_137),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_128),
.Y(n_204)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_130),
.B(n_149),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_119),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_191),
.B1(n_166),
.B2(n_178),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_193),
.B(n_195),
.C(n_211),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_129),
.B1(n_126),
.B2(n_114),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

OAI22x1_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_126),
.B1(n_145),
.B2(n_122),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_206),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_153),
.B(n_116),
.CI(n_143),
.CON(n_198),
.SN(n_198)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_198),
.B(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_145),
.C(n_131),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_166),
.C(n_165),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_203),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_205),
.B(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_144),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

AO21x2_ASAP7_75t_L g213 ( 
.A1(n_158),
.A2(n_150),
.B(n_140),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_179),
.B(n_157),
.Y(n_240)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_167),
.B1(n_154),
.B2(n_181),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_225),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_222),
.C(n_231),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_186),
.Y(n_221)
);

NAND4xp25_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_198),
.C(n_207),
.D(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_159),
.C(n_165),
.Y(n_222)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_176),
.A3(n_175),
.B1(n_160),
.B2(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_239),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_151),
.B1(n_155),
.B2(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_184),
.C(n_183),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_198),
.B(n_173),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_236),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_2),
.C(n_3),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_163),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_241),
.B(n_199),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_163),
.B(n_156),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_245),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_258),
.B1(n_185),
.B2(n_180),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_217),
.B(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_254),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_212),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_189),
.B(n_168),
.Y(n_274)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_256),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_191),
.A3(n_192),
.B1(n_213),
.B2(n_197),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_192),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_261),
.C(n_231),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_213),
.B1(n_190),
.B2(n_196),
.Y(n_258)
);

OAI322xp33_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_212),
.A3(n_193),
.B1(n_213),
.B2(n_208),
.C1(n_214),
.C2(n_210),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_249),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_193),
.CI(n_213),
.CON(n_260),
.SN(n_260)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_220),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_156),
.C(n_168),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_225),
.B1(n_229),
.B2(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_279),
.B(n_255),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_269),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_233),
.B(n_220),
.C(n_223),
.D(n_228),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_235),
.B1(n_226),
.B2(n_216),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_235),
.B1(n_219),
.B2(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_185),
.C(n_189),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_277),
.A2(n_262),
.B(n_260),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_161),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_4),
.B(n_7),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_286),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_261),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_252),
.B1(n_244),
.B2(n_253),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_254),
.B1(n_274),
.B2(n_265),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_269),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_263),
.B1(n_270),
.B2(n_257),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_298),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_267),
.C(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_300),
.C(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_290),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_264),
.B1(n_273),
.B2(n_272),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_291),
.B(n_282),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_247),
.C(n_268),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_247),
.C(n_271),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_283),
.B(n_293),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_308),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_309),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_283),
.B(n_292),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_265),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_292),
.B1(n_285),
.B2(n_260),
.Y(n_311)
);

AOI321xp33_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_295),
.A3(n_301),
.B1(n_300),
.B2(n_296),
.C(n_304),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_294),
.C(n_285),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_310),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_18),
.C(n_14),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_279),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_17),
.C(n_18),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_324),
.B(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_4),
.C(n_16),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_4),
.B(n_16),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_320),
.C(n_17),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);


endmodule