module fake_jpeg_21228_n_43 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_43);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NAND2x1_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_5),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_22),
.B(n_2),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_29),
.B1(n_20),
.B2(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_21),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_31),
.B1(n_29),
.B2(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_19),
.C(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_23),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_37),
.C(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_36),
.C(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_23),
.B1(n_5),
.B2(n_6),
.Y(n_42)
);

AOI221xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.C(n_34),
.Y(n_43)
);


endmodule