module fake_jpeg_1342_n_192 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_34),
.Y(n_84)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_0),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_11),
.Y(n_82)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_34),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_11),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_14),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_14),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_22),
.B1(n_21),
.B2(n_0),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_22),
.C(n_4),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_8),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_40),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_10),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_73),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_33),
.A2(n_12),
.B1(n_36),
.B2(n_34),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_50),
.B1(n_61),
.B2(n_86),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_93),
.B1(n_104),
.B2(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_55),
.B1(n_58),
.B2(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_111),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_59),
.B1(n_70),
.B2(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_71),
.B(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_127),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_122),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_85),
.B(n_84),
.C(n_64),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_113),
.B1(n_120),
.B2(n_130),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_79),
.B(n_81),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_79),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_60),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_126),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_70),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_64),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_111),
.C(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_96),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_91),
.B1(n_110),
.B2(n_95),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_139),
.B(n_118),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_95),
.B1(n_110),
.B2(n_100),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_149),
.Y(n_160)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_114),
.B1(n_126),
.B2(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_123),
.C(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_129),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_160),
.A2(n_135),
.B1(n_140),
.B2(n_141),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_167),
.B1(n_169),
.B2(n_155),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_170),
.B(n_155),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_140),
.B(n_147),
.C(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_160),
.B1(n_161),
.B2(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_173),
.B1(n_170),
.B2(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_150),
.C(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_176),
.C(n_164),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_143),
.CI(n_134),
.CON(n_173),
.SN(n_173)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_175),
.B(n_170),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_137),
.C(n_168),
.Y(n_176)
);

NOR2xp67_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_181),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_173),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_189),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_188),
.B1(n_183),
.B2(n_184),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_191),
.Y(n_192)
);


endmodule