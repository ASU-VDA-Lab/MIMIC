module fake_jpeg_75_n_545 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_545);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_51),
.Y(n_165)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_53),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_60),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g166 ( 
.A(n_61),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_13),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_48),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_75),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_14),
.Y(n_90)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_14),
.Y(n_93)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_98),
.A2(n_22),
.B(n_32),
.Y(n_170)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_22),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_27),
.B(n_36),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_50),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_109),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_51),
.A2(n_37),
.B1(n_47),
.B2(n_28),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_113),
.A2(n_144),
.B1(n_147),
.B2(n_26),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_32),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_54),
.A2(n_59),
.B1(n_100),
.B2(n_55),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_124),
.A2(n_150),
.B1(n_45),
.B2(n_17),
.Y(n_215)
);

OR2x4_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_22),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_139),
.C(n_35),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_71),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_94),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_37),
.B1(n_47),
.B2(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_44),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_145),
.B(n_152),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_70),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_39),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_90),
.B(n_22),
.Y(n_212)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_80),
.B1(n_64),
.B2(n_65),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_177),
.B1(n_192),
.B2(n_206),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_173),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_106),
.A2(n_164),
.B1(n_107),
.B2(n_151),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_179),
.Y(n_223)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

AO22x1_ASAP7_75t_SL g184 ( 
.A1(n_116),
.A2(n_76),
.B1(n_88),
.B2(n_63),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_212),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_195),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_136),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_213),
.Y(n_229)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_147),
.B1(n_126),
.B2(n_135),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_191),
.B(n_200),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_85),
.B1(n_81),
.B2(n_68),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_198),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_199),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_36),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_165),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_201),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_203),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_207),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_124),
.A2(n_96),
.B1(n_92),
.B2(n_26),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_211),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_35),
.B1(n_31),
.B2(n_48),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_215),
.B1(n_31),
.B2(n_46),
.Y(n_236)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_38),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_219),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_172),
.A2(n_144),
.B1(n_113),
.B2(n_87),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_232),
.B1(n_257),
.B2(n_136),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_114),
.C(n_117),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_224),
.C(n_237),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_236),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_89),
.B1(n_91),
.B2(n_162),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_46),
.B(n_16),
.C(n_19),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g277 ( 
.A(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_177),
.A2(n_184),
.B1(n_192),
.B2(n_173),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_215),
.B1(n_217),
.B2(n_211),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_258),
.A2(n_189),
.B1(n_230),
.B2(n_178),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_224),
.A2(n_184),
.B1(n_214),
.B2(n_173),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_265),
.B1(n_287),
.B2(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_174),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_264),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_223),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_267),
.Y(n_303)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_174),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_127),
.B1(n_121),
.B2(n_154),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_268),
.B1(n_280),
.B2(n_284),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_194),
.B1(n_162),
.B2(n_207),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_224),
.B(n_186),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_R g299 ( 
.A(n_269),
.B(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_271),
.B(n_230),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_171),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_273),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_188),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_205),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_285),
.C(n_221),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_176),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_225),
.A2(n_181),
.B1(n_183),
.B2(n_115),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_180),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_286),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_228),
.A2(n_121),
.B1(n_134),
.B2(n_132),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_138),
.C(n_137),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_223),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_236),
.A2(n_163),
.B1(n_143),
.B2(n_132),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_289),
.A2(n_298),
.B1(n_316),
.B2(n_220),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_229),
.B1(n_230),
.B2(n_236),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_290),
.A2(n_319),
.B1(n_284),
.B2(n_270),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_229),
.B(n_253),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_291),
.A2(n_293),
.B(n_294),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_230),
.B(n_253),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_229),
.B(n_245),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_313),
.C(n_315),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_266),
.A2(n_245),
.B1(n_233),
.B2(n_256),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_289),
.B1(n_287),
.B2(n_310),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_261),
.A2(n_256),
.B(n_233),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_308),
.B(n_311),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_264),
.A2(n_249),
.B(n_244),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_243),
.B(n_249),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_318),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_250),
.C(n_221),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_250),
.C(n_252),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_260),
.A2(n_238),
.B1(n_244),
.B2(n_203),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_252),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_317),
.B(n_312),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_239),
.C(n_241),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_238),
.B1(n_231),
.B2(n_254),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_292),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_323),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_298),
.B1(n_311),
.B2(n_302),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_300),
.A2(n_270),
.B1(n_286),
.B2(n_262),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_292),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_327),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_314),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_315),
.Y(n_359)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_290),
.A2(n_277),
.B1(n_268),
.B2(n_280),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_345),
.B1(n_346),
.B2(n_300),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_278),
.B(n_277),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_334),
.A2(n_341),
.B(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_303),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_338),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_295),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_343),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_293),
.A2(n_277),
.B(n_283),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_342),
.B(n_350),
.Y(n_357)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

A2O1A1O1Ixp25_ASAP7_75t_L g348 ( 
.A1(n_296),
.A2(n_269),
.B(n_285),
.C(n_282),
.D(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_263),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_349),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_320),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_351),
.B(n_353),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_312),
.B(n_222),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_313),
.Y(n_355)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_313),
.C(n_302),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_379),
.C(n_321),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_355),
.B(n_336),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_358),
.A2(n_333),
.B1(n_345),
.B2(n_329),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_361),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_331),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_317),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_364),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_317),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_350),
.B(n_315),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_367),
.B(n_374),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_370),
.B1(n_371),
.B2(n_381),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_304),
.B1(n_318),
.B2(n_308),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_322),
.A2(n_318),
.B1(n_299),
.B2(n_305),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_338),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_294),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_378),
.B(n_326),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_299),
.C(n_305),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_322),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_382),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_324),
.A2(n_299),
.B1(n_297),
.B2(n_276),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_251),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_347),
.A2(n_328),
.B1(n_327),
.B2(n_323),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_383),
.A2(n_321),
.B1(n_341),
.B2(n_349),
.Y(n_390)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_409),
.B1(n_255),
.B2(n_254),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_397),
.B1(n_410),
.B2(n_235),
.Y(n_437)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_384),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_392),
.B(n_407),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_401),
.Y(n_417)
);

BUFx4f_ASAP7_75t_SL g394 ( 
.A(n_385),
.Y(n_394)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_395),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_396),
.B(n_402),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_369),
.A2(n_335),
.B1(n_351),
.B2(n_353),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_399),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_359),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_362),
.B(n_334),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_404),
.Y(n_423)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_405),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_406),
.A2(n_409),
.B1(n_360),
.B2(n_391),
.Y(n_427)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_241),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_408),
.B(n_384),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_358),
.A2(n_332),
.B1(n_339),
.B2(n_337),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_383),
.A2(n_348),
.B1(n_276),
.B2(n_220),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_222),
.C(n_247),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_412),
.C(n_414),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_247),
.C(n_239),
.Y(n_412)
);

AO21x1_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_235),
.B(n_234),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_413),
.A2(n_376),
.B(n_381),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_247),
.C(n_234),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_420),
.A2(n_437),
.B1(n_218),
.B2(n_198),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_379),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_426),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_398),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_441),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_370),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_427),
.A2(n_428),
.B1(n_435),
.B2(n_187),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_406),
.A2(n_377),
.B1(n_360),
.B2(n_372),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_382),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_440),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_371),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_201),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_415),
.A2(n_377),
.B(n_366),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_432),
.A2(n_420),
.B(n_437),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_390),
.A2(n_375),
.B1(n_255),
.B2(n_254),
.Y(n_435)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_401),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_412),
.B(n_235),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_424),
.A2(n_394),
.B1(n_397),
.B2(n_413),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_442),
.A2(n_444),
.B1(n_445),
.B2(n_456),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_416),
.A2(n_394),
.B1(n_400),
.B2(n_410),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_389),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_458),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_414),
.C(n_389),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_451),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_396),
.C(n_402),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_423),
.A2(n_419),
.B(n_427),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_452),
.A2(n_457),
.B(n_462),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_421),
.Y(n_468)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_433),
.A2(n_143),
.B1(n_163),
.B2(n_154),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_428),
.A2(n_208),
.B(n_130),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_175),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_464),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_460),
.A2(n_438),
.B1(n_435),
.B2(n_422),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_439),
.B(n_179),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_463),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_423),
.A2(n_46),
.B(n_17),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_119),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_153),
.C(n_134),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_468),
.B(n_0),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_432),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_469),
.B(n_471),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_431),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_426),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_477),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_438),
.Y(n_476)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_439),
.Y(n_477)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_445),
.A2(n_38),
.B(n_16),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_479),
.A2(n_19),
.B(n_1),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_160),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_153),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_481),
.B(n_483),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_484),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_464),
.B(n_129),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_129),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_489),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_SL g487 ( 
.A(n_465),
.B(n_451),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_487),
.A2(n_493),
.B(n_502),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_474),
.A2(n_461),
.B1(n_458),
.B2(n_454),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_446),
.C(n_443),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_490),
.B(n_491),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_463),
.B1(n_443),
.B2(n_48),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_13),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_492),
.B(n_495),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_45),
.B(n_38),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_45),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_467),
.A2(n_19),
.B1(n_17),
.B2(n_2),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_2),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_501),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_1),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_499),
.B(n_466),
.Y(n_504)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_477),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_511),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_499),
.A2(n_466),
.B(n_467),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_509),
.A2(n_497),
.B(n_498),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_1),
.Y(n_510)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_510),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_1),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_2),
.C(n_3),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_514),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_2),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_516),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_3),
.C(n_4),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_5),
.C(n_6),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_517),
.B(n_5),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_508),
.A2(n_489),
.B1(n_486),
.B2(n_488),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_518),
.B(n_520),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_493),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_522),
.A2(n_505),
.B(n_513),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_523),
.B(n_7),
.Y(n_531)
);

OAI21xp33_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_516),
.B(n_517),
.Y(n_530)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_506),
.A2(n_7),
.B(n_8),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_SL g534 ( 
.A1(n_525),
.A2(n_522),
.B(n_528),
.C(n_515),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_529),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_531),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_519),
.Y(n_533)
);

A2O1A1O1Ixp25_ASAP7_75t_L g539 ( 
.A1(n_533),
.A2(n_534),
.B(n_535),
.C(n_526),
.D(n_9),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_527),
.B(n_510),
.C(n_503),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_532),
.Y(n_537)
);

OAI321xp33_ASAP7_75t_L g542 ( 
.A1(n_537),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_536),
.C(n_532),
.Y(n_542)
);

OAI321xp33_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_532),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_8),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_541),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_10),
.Y(n_541)
);

NOR3xp33_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_538),
.C(n_542),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_544),
.A2(n_11),
.B(n_12),
.Y(n_545)
);


endmodule