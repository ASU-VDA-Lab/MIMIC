module real_aes_18418_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1441;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1914;
wire n_1648;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_1951;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1671;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1931;
wire n_1691;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1960 ( .A(n_0), .Y(n_1960) );
OAI22xp5_ASAP7_75t_L g1923 ( .A1(n_1), .A2(n_85), .B1(n_722), .B2(n_1924), .Y(n_1923) );
INVxp67_ASAP7_75t_SL g1936 ( .A(n_1), .Y(n_1936) );
INVx1_ASAP7_75t_L g782 ( .A(n_2), .Y(n_782) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_2), .A2(n_372), .B1(n_807), .B2(n_809), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g775 ( .A1(n_3), .A2(n_199), .B1(n_595), .B2(n_718), .C(n_776), .Y(n_775) );
AOI222xp33_ASAP7_75t_L g820 ( .A1(n_3), .A2(n_131), .B1(n_335), .B2(n_442), .C1(n_821), .C2(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g388 ( .A(n_4), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_4), .B(n_398), .Y(n_470) );
AND2x2_ASAP7_75t_L g583 ( .A(n_4), .B(n_280), .Y(n_583) );
AND2x2_ASAP7_75t_L g605 ( .A(n_4), .B(n_544), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g1976 ( .A1(n_5), .A2(n_549), .B(n_1436), .C(n_1977), .Y(n_1976) );
INVx1_ASAP7_75t_L g1986 ( .A(n_5), .Y(n_1986) );
INVx1_ASAP7_75t_L g936 ( .A(n_6), .Y(n_936) );
INVx1_ASAP7_75t_L g1664 ( .A(n_7), .Y(n_1664) );
INVx1_ASAP7_75t_L g1300 ( .A(n_8), .Y(n_1300) );
INVx1_ASAP7_75t_L g1408 ( .A(n_9), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_10), .A2(n_174), .B1(n_970), .B2(n_1502), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_10), .A2(n_174), .B1(n_530), .B2(n_1289), .Y(n_1514) );
INVx1_ASAP7_75t_L g425 ( .A(n_11), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g1503 ( .A1(n_12), .A2(n_303), .B1(n_390), .B2(n_541), .Y(n_1503) );
OAI22xp33_ASAP7_75t_L g1509 ( .A1(n_12), .A2(n_303), .B1(n_896), .B2(n_1510), .Y(n_1509) );
OAI211xp5_ASAP7_75t_L g1661 ( .A1(n_13), .A2(n_766), .B(n_1662), .C(n_1663), .Y(n_1661) );
INVx1_ASAP7_75t_L g1675 ( .A(n_13), .Y(n_1675) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_14), .A2(n_87), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
AOI221xp5_ASAP7_75t_L g1317 ( .A1(n_14), .A2(n_23), .B1(n_1005), .B2(n_1318), .C(n_1320), .Y(n_1317) );
INVx1_ASAP7_75t_L g1904 ( .A(n_15), .Y(n_1904) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_16), .A2(n_34), .B1(n_828), .B2(n_1167), .Y(n_1195) );
INVx1_ASAP7_75t_L g1232 ( .A(n_16), .Y(n_1232) );
OAI211xp5_ASAP7_75t_L g1570 ( .A1(n_17), .A2(n_513), .B(n_1571), .C(n_1572), .Y(n_1570) );
INVx1_ASAP7_75t_L g1579 ( .A(n_17), .Y(n_1579) );
INVx1_ASAP7_75t_L g1595 ( .A(n_18), .Y(n_1595) );
INVx1_ASAP7_75t_L g1445 ( .A(n_19), .Y(n_1445) );
OAI211xp5_ASAP7_75t_L g1454 ( .A1(n_19), .A2(n_513), .B(n_732), .C(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1350 ( .A(n_20), .Y(n_1350) );
INVx1_ASAP7_75t_L g631 ( .A(n_21), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_22), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g1309 ( .A1(n_23), .A2(n_262), .B1(n_821), .B2(n_828), .Y(n_1309) );
INVx1_ASAP7_75t_L g1412 ( .A(n_24), .Y(n_1412) );
INVx2_ASAP7_75t_L g416 ( .A(n_25), .Y(n_416) );
INVx1_ASAP7_75t_L g1557 ( .A(n_26), .Y(n_1557) );
OAI22xp33_ASAP7_75t_L g526 ( .A1(n_27), .A2(n_250), .B1(n_527), .B2(n_530), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_27), .A2(n_250), .B1(n_566), .B2(n_568), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g1717 ( .A1(n_28), .A2(n_30), .B1(n_1688), .B2(n_1696), .Y(n_1717) );
OAI22xp33_ASAP7_75t_L g1614 ( .A1(n_29), .A2(n_313), .B1(n_390), .B2(n_1615), .Y(n_1614) );
OAI22xp5_ASAP7_75t_L g1622 ( .A1(n_29), .A2(n_313), .B1(n_1510), .B2(n_1623), .Y(n_1622) );
XNOR2xp5_ASAP7_75t_L g1897 ( .A(n_30), .B(n_1898), .Y(n_1897) );
AOI22xp33_ASAP7_75t_L g1945 ( .A1(n_30), .A2(n_1946), .B1(n_1949), .B2(n_1988), .Y(n_1945) );
INVx1_ASAP7_75t_L g1963 ( .A(n_31), .Y(n_1963) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_32), .A2(n_244), .B1(n_503), .B2(n_506), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_32), .A2(n_244), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_33), .A2(n_237), .B1(n_591), .B2(n_610), .C(n_611), .Y(n_609) );
INVxp67_ASAP7_75t_SL g637 ( .A(n_33), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g1214 ( .A1(n_34), .A2(n_52), .B1(n_617), .B2(n_1215), .C(n_1216), .Y(n_1214) );
INVx1_ASAP7_75t_L g1304 ( .A(n_35), .Y(n_1304) );
INVx1_ASAP7_75t_L g831 ( .A(n_36), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_37), .A2(n_318), .B1(n_527), .B2(n_896), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_37), .A2(n_346), .B1(n_568), .B2(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g1420 ( .A(n_38), .Y(n_1420) );
OA222x2_ASAP7_75t_L g1111 ( .A1(n_39), .A2(n_94), .B1(n_275), .B2(n_1112), .C1(n_1114), .C2(n_1118), .Y(n_1111) );
INVx1_ASAP7_75t_L g1165 ( .A(n_39), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_40), .Y(n_383) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_40), .B(n_381), .Y(n_1689) );
INVx1_ASAP7_75t_L g706 ( .A(n_41), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g1756 ( .A1(n_41), .A2(n_222), .B1(n_1696), .B2(n_1757), .Y(n_1756) );
XNOR2xp5_ASAP7_75t_L g770 ( .A(n_42), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g1483 ( .A(n_43), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_44), .A2(n_350), .B1(n_616), .B2(n_630), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g1269 ( .A(n_44), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_45), .A2(n_114), .B1(n_591), .B2(n_592), .C(n_595), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_45), .A2(n_121), .B1(n_658), .B2(n_663), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_46), .A2(n_238), .B1(n_1037), .B2(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1218 ( .A(n_46), .Y(n_1218) );
INVx1_ASAP7_75t_L g1602 ( .A(n_47), .Y(n_1602) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_48), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_49), .A2(n_299), .B1(n_541), .B2(n_1353), .Y(n_1352) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_49), .A2(n_205), .B1(n_896), .B2(n_1361), .Y(n_1360) );
XNOR2xp5_ASAP7_75t_L g1546 ( .A(n_50), .B(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1066 ( .A(n_51), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_52), .A2(n_342), .B1(n_828), .B2(n_1203), .Y(n_1202) );
INVxp67_ASAP7_75t_SL g1303 ( .A(n_53), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_53), .A2(n_196), .B1(n_791), .B2(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g525 ( .A(n_54), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g547 ( .A1(n_54), .A2(n_548), .B(n_549), .C(n_554), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g1364 ( .A1(n_55), .A2(n_151), .B1(n_1365), .B2(n_1366), .Y(n_1364) );
AOI22xp33_ASAP7_75t_SL g1394 ( .A1(n_55), .A2(n_279), .B1(n_663), .B2(n_1389), .Y(n_1394) );
INVx1_ASAP7_75t_L g1637 ( .A(n_56), .Y(n_1637) );
INVx1_ASAP7_75t_L g1073 ( .A(n_57), .Y(n_1073) );
INVxp67_ASAP7_75t_SL g1922 ( .A(n_58), .Y(n_1922) );
OAI22xp5_ASAP7_75t_L g1937 ( .A1(n_58), .A2(n_85), .B1(n_1938), .B2(n_1939), .Y(n_1937) );
OAI211xp5_ASAP7_75t_L g1616 ( .A1(n_59), .A2(n_973), .B(n_977), .C(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1626 ( .A(n_59), .Y(n_1626) );
CKINVDCx5p33_ASAP7_75t_R g1136 ( .A(n_60), .Y(n_1136) );
INVx1_ASAP7_75t_L g620 ( .A(n_61), .Y(n_620) );
INVx1_ASAP7_75t_L g1313 ( .A(n_62), .Y(n_1313) );
INVx1_ASAP7_75t_L g930 ( .A(n_63), .Y(n_930) );
INVx1_ASAP7_75t_L g628 ( .A(n_64), .Y(n_628) );
OAI322xp33_ASAP7_75t_L g635 ( .A1(n_64), .A2(n_408), .A3(n_636), .B1(n_643), .B2(n_651), .C1(n_665), .C2(n_667), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g1257 ( .A1(n_65), .A2(n_286), .B1(n_616), .B2(n_1258), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_65), .A2(n_269), .B1(n_663), .B2(n_1158), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g1770 ( .A1(n_66), .A2(n_236), .B1(n_1688), .B2(n_1693), .Y(n_1770) );
OAI22xp33_ASAP7_75t_L g1666 ( .A1(n_67), .A2(n_166), .B1(n_1452), .B2(n_1628), .Y(n_1666) );
OAI22xp5_ASAP7_75t_L g1676 ( .A1(n_67), .A2(n_166), .B1(n_892), .B2(n_1447), .Y(n_1676) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_68), .Y(n_1302) );
INVx1_ASAP7_75t_L g1335 ( .A(n_69), .Y(n_1335) );
AOI22xp5_ASAP7_75t_L g1703 ( .A1(n_69), .A2(n_363), .B1(n_1696), .B2(n_1704), .Y(n_1703) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_70), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_71), .A2(n_86), .B1(n_1199), .B2(n_1201), .Y(n_1198) );
INVx1_ASAP7_75t_L g1217 ( .A(n_71), .Y(n_1217) );
OAI22xp33_ASAP7_75t_SL g1249 ( .A1(n_72), .A2(n_277), .B1(n_951), .B2(n_1135), .Y(n_1249) );
INVx1_ASAP7_75t_L g1284 ( .A(n_72), .Y(n_1284) );
INVx1_ASAP7_75t_L g1486 ( .A(n_73), .Y(n_1486) );
INVx1_ASAP7_75t_L g744 ( .A(n_74), .Y(n_744) );
INVx1_ASAP7_75t_L g1519 ( .A(n_75), .Y(n_1519) );
AOI21xp33_ASAP7_75t_L g1016 ( .A1(n_76), .A2(n_610), .B(n_1017), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1044 ( .A1(n_76), .A2(n_295), .B1(n_1037), .B2(n_1045), .C(n_1046), .Y(n_1044) );
INVx1_ASAP7_75t_L g713 ( .A(n_77), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_78), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_79), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g1771 ( .A1(n_80), .A2(n_339), .B1(n_1696), .B2(n_1757), .Y(n_1771) );
INVx1_ASAP7_75t_L g1598 ( .A(n_81), .Y(n_1598) );
OAI22xp33_ASAP7_75t_L g878 ( .A1(n_82), .A2(n_141), .B1(n_390), .B2(n_879), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_82), .A2(n_141), .B1(n_768), .B2(n_896), .Y(n_895) );
OAI222xp33_ASAP7_75t_L g984 ( .A1(n_83), .A2(n_92), .B1(n_101), .B2(n_698), .C1(n_985), .C2(n_990), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g1724 ( .A1(n_84), .A2(n_150), .B1(n_1688), .B2(n_1693), .Y(n_1724) );
INVx1_ASAP7_75t_L g1236 ( .A(n_86), .Y(n_1236) );
INVx1_ASAP7_75t_L g1334 ( .A(n_87), .Y(n_1334) );
INVx1_ASAP7_75t_L g1926 ( .A(n_88), .Y(n_1926) );
INVx1_ASAP7_75t_L g933 ( .A(n_89), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_90), .A2(n_93), .B1(n_566), .B2(n_1062), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1100 ( .A1(n_90), .A2(n_93), .B1(n_530), .B2(n_1101), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_91), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_94), .A2(n_215), .B1(n_1152), .B2(n_1154), .C(n_1156), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_95), .A2(n_326), .B1(n_478), .B2(n_791), .Y(n_1225) );
INVx1_ASAP7_75t_L g1238 ( .A(n_95), .Y(n_1238) );
INVx1_ASAP7_75t_L g1126 ( .A(n_96), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_96), .A2(n_163), .B1(n_1038), .B2(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1927 ( .A(n_97), .Y(n_1927) );
INVx1_ASAP7_75t_L g1079 ( .A(n_98), .Y(n_1079) );
XOR2x2_ASAP7_75t_L g1458 ( .A(n_99), .B(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1918 ( .A(n_100), .Y(n_1918) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_101), .A2(n_371), .B1(n_1027), .B2(n_1031), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1620 ( .A1(n_102), .A2(n_195), .B1(n_1447), .B2(n_1466), .Y(n_1620) );
OAI22xp33_ASAP7_75t_L g1627 ( .A1(n_102), .A2(n_195), .B1(n_904), .B2(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g463 ( .A(n_103), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g510 ( .A1(n_104), .A2(n_511), .B(n_513), .C(n_517), .Y(n_510) );
INVx1_ASAP7_75t_L g564 ( .A(n_104), .Y(n_564) );
INVx1_ASAP7_75t_L g449 ( .A(n_105), .Y(n_449) );
INVx1_ASAP7_75t_L g1956 ( .A(n_106), .Y(n_1956) );
INVx1_ASAP7_75t_L g1978 ( .A(n_107), .Y(n_1978) );
AOI22xp5_ASAP7_75t_L g1711 ( .A1(n_108), .A2(n_369), .B1(n_1688), .B2(n_1693), .Y(n_1711) );
INVx1_ASAP7_75t_L g1463 ( .A(n_109), .Y(n_1463) );
XOR2x2_ASAP7_75t_L g912 ( .A(n_110), .B(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_111), .A2(n_187), .B1(n_601), .B2(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1040 ( .A(n_111), .Y(n_1040) );
XNOR2xp5_ASAP7_75t_L g1632 ( .A(n_112), .B(n_1633), .Y(n_1632) );
CKINVDCx5p33_ASAP7_75t_R g1312 ( .A(n_113), .Y(n_1312) );
INVx1_ASAP7_75t_L g648 ( .A(n_114), .Y(n_648) );
INVx1_ASAP7_75t_L g522 ( .A(n_115), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_116), .A2(n_347), .B1(n_1199), .B2(n_1307), .Y(n_1306) );
AOI221xp5_ASAP7_75t_L g1331 ( .A1(n_116), .A2(n_234), .B1(n_616), .B2(n_617), .C(n_1332), .Y(n_1331) );
OAI211xp5_ASAP7_75t_L g1504 ( .A1(n_117), .A2(n_549), .B(n_957), .C(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1513 ( .A(n_117), .Y(n_1513) );
INVx1_ASAP7_75t_L g1641 ( .A(n_118), .Y(n_1641) );
AOI22xp5_ASAP7_75t_SL g1712 ( .A1(n_119), .A2(n_248), .B1(n_1696), .B2(n_1704), .Y(n_1712) );
INVx1_ASAP7_75t_L g1239 ( .A(n_120), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_121), .A2(n_364), .B1(n_614), .B2(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g1905 ( .A(n_122), .Y(n_1905) );
AOI22xp33_ASAP7_75t_L g1933 ( .A1(n_122), .A2(n_316), .B1(n_779), .B2(n_1005), .Y(n_1933) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_123), .A2(n_173), .B1(n_541), .B2(n_724), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_123), .A2(n_173), .B1(n_1093), .B2(n_1095), .Y(n_1092) );
OAI22xp33_ASAP7_75t_L g1438 ( .A1(n_124), .A2(n_129), .B1(n_879), .B2(n_1439), .Y(n_1438) );
OAI22xp33_ASAP7_75t_L g1449 ( .A1(n_124), .A2(n_129), .B1(n_1093), .B2(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1618 ( .A(n_125), .Y(n_1618) );
OAI22xp5_ASAP7_75t_L g1575 ( .A1(n_126), .A2(n_203), .B1(n_530), .B2(n_768), .Y(n_1575) );
OAI22xp5_ASAP7_75t_L g1580 ( .A1(n_126), .A2(n_242), .B1(n_1447), .B2(n_1581), .Y(n_1580) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_127), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_127), .A2(n_199), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g381 ( .A(n_128), .Y(n_381) );
INVx1_ASAP7_75t_L g1914 ( .A(n_130), .Y(n_1914) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_131), .A2(n_341), .B1(n_614), .B2(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_132), .A2(n_340), .B1(n_541), .B2(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_132), .A2(n_340), .B1(n_503), .B2(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g717 ( .A(n_133), .Y(n_717) );
INVx1_ASAP7_75t_L g1554 ( .A(n_134), .Y(n_1554) );
INVx1_ASAP7_75t_L g917 ( .A(n_135), .Y(n_917) );
OAI211xp5_ASAP7_75t_L g1461 ( .A1(n_136), .A2(n_493), .B(n_549), .C(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1473 ( .A(n_136), .Y(n_1473) );
INVx1_ASAP7_75t_L g1507 ( .A(n_137), .Y(n_1507) );
OAI211xp5_ASAP7_75t_L g1511 ( .A1(n_137), .A2(n_511), .B(n_766), .C(n_1512), .Y(n_1511) );
AOI22xp5_ASAP7_75t_L g1708 ( .A1(n_138), .A2(n_349), .B1(n_1693), .B2(n_1704), .Y(n_1708) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_139), .A2(n_179), .B1(n_1127), .B2(n_1128), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_139), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1967 ( .A(n_140), .Y(n_1967) );
CKINVDCx5p33_ASAP7_75t_R g1210 ( .A(n_142), .Y(n_1210) );
INVx1_ASAP7_75t_L g1964 ( .A(n_143), .Y(n_1964) );
INVx1_ASAP7_75t_L g1966 ( .A(n_144), .Y(n_1966) );
XOR2xp5_ASAP7_75t_L g1950 ( .A(n_145), .B(n_1951), .Y(n_1950) );
OAI211xp5_ASAP7_75t_SL g772 ( .A1(n_146), .A2(n_773), .B(n_774), .C(n_780), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_146), .A2(n_361), .B1(n_698), .B2(n_805), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g1980 ( .A1(n_147), .A2(n_160), .B1(n_567), .B2(n_1345), .Y(n_1980) );
OAI22xp33_ASAP7_75t_L g1987 ( .A1(n_147), .A2(n_160), .B1(n_527), .B2(n_1357), .Y(n_1987) );
INVx1_ASAP7_75t_L g1599 ( .A(n_148), .Y(n_1599) );
INVx1_ASAP7_75t_L g1489 ( .A(n_149), .Y(n_1489) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_151), .A2(n_256), .B1(n_1385), .B2(n_1387), .Y(n_1384) );
INVx1_ASAP7_75t_L g1902 ( .A(n_152), .Y(n_1902) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_153), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_154), .A2(n_321), .B1(n_1345), .B2(n_1447), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1451 ( .A1(n_154), .A2(n_321), .B1(n_1101), .B2(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1444 ( .A(n_155), .Y(n_1444) );
INVx1_ASAP7_75t_L g1979 ( .A(n_156), .Y(n_1979) );
OAI211xp5_ASAP7_75t_L g1984 ( .A1(n_156), .A2(n_513), .B(n_1471), .C(n_1985), .Y(n_1984) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_157), .A2(n_346), .B1(n_506), .B2(n_530), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g968 ( .A1(n_157), .A2(n_318), .B1(n_390), .B2(n_879), .Y(n_968) );
INVx1_ASAP7_75t_L g1957 ( .A(n_158), .Y(n_1957) );
INVx1_ASAP7_75t_L g1402 ( .A(n_159), .Y(n_1402) );
INVx1_ASAP7_75t_L g446 ( .A(n_161), .Y(n_446) );
INVx1_ASAP7_75t_L g720 ( .A(n_162), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_163), .A2(n_201), .B1(n_1029), .B2(n_1138), .Y(n_1137) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_164), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_164), .A2(n_307), .B1(n_614), .B2(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_165), .A2(n_357), .B1(n_1447), .B2(n_1466), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_165), .A2(n_357), .B1(n_1289), .B2(n_1357), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_167), .A2(n_215), .B1(n_581), .B2(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1166 ( .A(n_167), .Y(n_1166) );
OAI211xp5_ASAP7_75t_L g880 ( .A1(n_168), .A2(n_549), .B(n_881), .C(n_885), .Y(n_880) );
INVx1_ASAP7_75t_L g902 ( .A(n_168), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g1467 ( .A1(n_169), .A2(n_207), .B1(n_879), .B2(n_1439), .Y(n_1467) );
OAI22xp33_ASAP7_75t_L g1474 ( .A1(n_169), .A2(n_207), .B1(n_505), .B2(n_1450), .Y(n_1474) );
OAI22xp33_ASAP7_75t_L g1981 ( .A1(n_170), .A2(n_270), .B1(n_1439), .B2(n_1615), .Y(n_1981) );
OAI22xp33_ASAP7_75t_L g1983 ( .A1(n_170), .A2(n_270), .B1(n_505), .B2(n_1095), .Y(n_1983) );
INVx1_ASAP7_75t_L g1076 ( .A(n_171), .Y(n_1076) );
INVx1_ASAP7_75t_L g1561 ( .A(n_172), .Y(n_1561) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_175), .A2(n_352), .B1(n_493), .B2(n_1262), .C(n_1264), .Y(n_1261) );
INVx1_ASAP7_75t_L g1281 ( .A(n_175), .Y(n_1281) );
INVx1_ASAP7_75t_L g1251 ( .A(n_176), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_176), .A2(n_286), .B1(n_1158), .B2(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1648 ( .A(n_177), .Y(n_1648) );
CKINVDCx5p33_ASAP7_75t_R g1255 ( .A(n_178), .Y(n_1255) );
INVx1_ASAP7_75t_L g1283 ( .A(n_179), .Y(n_1283) );
INVx1_ASAP7_75t_L g1644 ( .A(n_180), .Y(n_1644) );
INVx1_ASAP7_75t_L g1349 ( .A(n_181), .Y(n_1349) );
OAI211xp5_ASAP7_75t_L g1358 ( .A1(n_181), .A2(n_766), .B(n_962), .C(n_1359), .Y(n_1358) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_182), .A2(n_513), .B(n_962), .C(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g976 ( .A(n_182), .Y(n_976) );
INVx1_ASAP7_75t_L g1574 ( .A(n_183), .Y(n_1574) );
OAI211xp5_ASAP7_75t_SL g1577 ( .A1(n_183), .A2(n_549), .B(n_973), .C(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1415 ( .A(n_184), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g1569 ( .A1(n_185), .A2(n_242), .B1(n_527), .B2(n_896), .Y(n_1569) );
OAI22xp33_ASAP7_75t_L g1582 ( .A1(n_185), .A2(n_203), .B1(n_390), .B2(n_879), .Y(n_1582) );
INVx1_ASAP7_75t_L g1506 ( .A(n_186), .Y(n_1506) );
INVxp67_ASAP7_75t_SL g1047 ( .A(n_187), .Y(n_1047) );
INVx1_ASAP7_75t_L g741 ( .A(n_188), .Y(n_741) );
INVx1_ASAP7_75t_L g1645 ( .A(n_189), .Y(n_1645) );
OAI22xp33_ASAP7_75t_L g1658 ( .A1(n_190), .A2(n_362), .B1(n_768), .B2(n_1659), .Y(n_1658) );
OAI22xp33_ASAP7_75t_L g1669 ( .A1(n_190), .A2(n_362), .B1(n_390), .B2(n_879), .Y(n_1669) );
INVx1_ASAP7_75t_L g1604 ( .A(n_191), .Y(n_1604) );
OAI211xp5_ASAP7_75t_L g1440 ( .A1(n_192), .A2(n_1088), .B(n_1441), .C(n_1443), .Y(n_1440) );
INVx1_ASAP7_75t_L g1456 ( .A(n_192), .Y(n_1456) );
INVx1_ASAP7_75t_L g1639 ( .A(n_193), .Y(n_1639) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_194), .A2(n_335), .B1(n_610), .B2(n_611), .C(n_798), .Y(n_797) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_194), .Y(n_825) );
INVxp67_ASAP7_75t_SL g1315 ( .A(n_196), .Y(n_1315) );
CKINVDCx5p33_ASAP7_75t_R g1134 ( .A(n_197), .Y(n_1134) );
INVx1_ASAP7_75t_L g1242 ( .A(n_198), .Y(n_1242) );
INVx1_ASAP7_75t_L g1753 ( .A(n_200), .Y(n_1753) );
INVx1_ASAP7_75t_L g1178 ( .A(n_201), .Y(n_1178) );
XNOR2xp5_ASAP7_75t_L g1589 ( .A(n_202), .B(n_1590), .Y(n_1589) );
AOI22xp5_ASAP7_75t_SL g1723 ( .A1(n_202), .A2(n_211), .B1(n_1696), .B2(n_1704), .Y(n_1723) );
INVx1_ASAP7_75t_L g1485 ( .A(n_204), .Y(n_1485) );
INVx1_ASAP7_75t_L g1347 ( .A(n_205), .Y(n_1347) );
INVx1_ASAP7_75t_L g1464 ( .A(n_206), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1470 ( .A1(n_206), .A2(n_513), .B(n_1471), .C(n_1472), .Y(n_1470) );
INVx1_ASAP7_75t_L g1015 ( .A(n_208), .Y(n_1015) );
AOI221x1_ASAP7_75t_SL g1035 ( .A1(n_208), .A2(n_288), .B1(n_1036), .B2(n_1037), .C(n_1039), .Y(n_1035) );
INVx1_ASAP7_75t_L g1407 ( .A(n_209), .Y(n_1407) );
AOI221x1_ASAP7_75t_SL g1120 ( .A1(n_210), .A2(n_283), .B1(n_1121), .B2(n_1124), .C(n_1125), .Y(n_1120) );
AOI21xp33_ASAP7_75t_L g1180 ( .A1(n_210), .A2(n_448), .B(n_1181), .Y(n_1180) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_212), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_212), .A2(n_217), .B1(n_597), .B2(n_630), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g1022 ( .A1(n_213), .A2(n_1023), .B(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g1048 ( .A(n_213), .Y(n_1048) );
INVx2_ASAP7_75t_L g1691 ( .A(n_214), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_214), .B(n_1692), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_214), .B(n_324), .Y(n_1699) );
AOI22xp5_ASAP7_75t_SL g1716 ( .A1(n_216), .A2(n_282), .B1(n_1693), .B2(n_1698), .Y(n_1716) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_217), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_218), .A2(n_315), .B1(n_597), .B2(n_601), .Y(n_596) );
INVx1_ASAP7_75t_L g656 ( .A(n_218), .Y(n_656) );
INVx1_ASAP7_75t_L g719 ( .A(n_219), .Y(n_719) );
INVx1_ASAP7_75t_L g1351 ( .A(n_220), .Y(n_1351) );
INVx1_ASAP7_75t_L g1058 ( .A(n_221), .Y(n_1058) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_223), .A2(n_348), .B1(n_1696), .B2(n_1698), .Y(n_1695) );
INVx1_ASAP7_75t_L g964 ( .A(n_224), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g1702 ( .A1(n_225), .A2(n_285), .B1(n_1688), .B2(n_1693), .Y(n_1702) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_226), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_227), .A2(n_359), .B1(n_1368), .B2(n_1369), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_227), .A2(n_233), .B1(n_1392), .B2(n_1393), .Y(n_1391) );
OAI211xp5_ASAP7_75t_L g1056 ( .A1(n_228), .A2(n_548), .B(n_977), .C(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1099 ( .A(n_228), .Y(n_1099) );
XOR2x2_ASAP7_75t_L g1497 ( .A(n_229), .B(n_1498), .Y(n_1497) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_230), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1594 ( .A(n_231), .Y(n_1594) );
AOI22xp5_ASAP7_75t_L g1709 ( .A1(n_232), .A2(n_306), .B1(n_1688), .B2(n_1696), .Y(n_1709) );
AOI22xp33_ASAP7_75t_SL g1382 ( .A1(n_233), .A2(n_354), .B1(n_779), .B2(n_1368), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_234), .A2(n_329), .B1(n_1036), .B2(n_1201), .Y(n_1295) );
INVx1_ASAP7_75t_L g937 ( .A(n_235), .Y(n_937) );
INVx1_ASAP7_75t_L g654 ( .A(n_237), .Y(n_654) );
INVx1_ASAP7_75t_L g1234 ( .A(n_238), .Y(n_1234) );
INVx2_ASAP7_75t_L g415 ( .A(n_239), .Y(n_415) );
INVx1_ASAP7_75t_L g458 ( .A(n_239), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_239), .B(n_416), .Y(n_586) );
INVx1_ASAP7_75t_L g1642 ( .A(n_240), .Y(n_1642) );
INVx1_ASAP7_75t_L g1421 ( .A(n_241), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_243), .A2(n_252), .B1(n_891), .B2(n_892), .Y(n_890) );
OAI22xp33_ASAP7_75t_L g903 ( .A1(n_243), .A2(n_252), .B1(n_527), .B2(n_904), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_245), .B(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_245), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_246), .Y(n_849) );
INVx1_ASAP7_75t_L g1573 ( .A(n_247), .Y(n_1573) );
INVx1_ASAP7_75t_L g982 ( .A(n_248), .Y(n_982) );
INVx1_ASAP7_75t_L g1413 ( .A(n_249), .Y(n_1413) );
INVx1_ASAP7_75t_L g1560 ( .A(n_251), .Y(n_1560) );
BUFx3_ASAP7_75t_L g422 ( .A(n_253), .Y(n_422) );
INVx1_ASAP7_75t_L g587 ( .A(n_254), .Y(n_587) );
INVx1_ASAP7_75t_L g731 ( .A(n_255), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_256), .A2(n_279), .B1(n_1377), .B2(n_1378), .Y(n_1376) );
INVx1_ASAP7_75t_L g1601 ( .A(n_257), .Y(n_1601) );
AOI22xp5_ASAP7_75t_L g1687 ( .A1(n_258), .A2(n_302), .B1(n_1688), .B2(n_1693), .Y(n_1687) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_259), .Y(n_672) );
OAI22xp5_ASAP7_75t_SL g1000 ( .A1(n_260), .A2(n_308), .B1(n_584), .B2(n_675), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_260), .Y(n_1010) );
INVx1_ASAP7_75t_L g1907 ( .A(n_261), .Y(n_1907) );
INVx1_ASAP7_75t_L g1333 ( .A(n_262), .Y(n_1333) );
INVx1_ASAP7_75t_L g1479 ( .A(n_263), .Y(n_1479) );
INVx1_ASAP7_75t_L g606 ( .A(n_264), .Y(n_606) );
INVx1_ASAP7_75t_L g1619 ( .A(n_265), .Y(n_1619) );
OAI211xp5_ASAP7_75t_SL g1624 ( .A1(n_265), .A2(n_513), .B(n_1043), .C(n_1625), .Y(n_1624) );
XOR2xp5_ASAP7_75t_L g404 ( .A(n_266), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g434 ( .A(n_267), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_268), .Y(n_845) );
AOI21xp33_ASAP7_75t_L g1252 ( .A1(n_269), .A2(n_1023), .B(n_1024), .Y(n_1252) );
INVx1_ASAP7_75t_L g926 ( .A(n_271), .Y(n_926) );
INVx1_ASAP7_75t_L g1071 ( .A(n_272), .Y(n_1071) );
INVx1_ASAP7_75t_L g1522 ( .A(n_273), .Y(n_1522) );
INVx1_ASAP7_75t_L g1558 ( .A(n_274), .Y(n_1558) );
INVx1_ASAP7_75t_L g1157 ( .A(n_275), .Y(n_1157) );
INVx1_ASAP7_75t_L g735 ( .A(n_276), .Y(n_735) );
INVx1_ASAP7_75t_L g1287 ( .A(n_277), .Y(n_1287) );
INVx1_ASAP7_75t_L g1913 ( .A(n_278), .Y(n_1913) );
AOI22xp33_ASAP7_75t_L g1930 ( .A1(n_278), .A2(n_327), .B1(n_779), .B2(n_1931), .Y(n_1930) );
BUFx3_ASAP7_75t_L g398 ( .A(n_280), .Y(n_398) );
INVx1_ASAP7_75t_L g544 ( .A(n_280), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_281), .Y(n_769) );
INVx1_ASAP7_75t_L g1177 ( .A(n_283), .Y(n_1177) );
INVx1_ASAP7_75t_L g1551 ( .A(n_284), .Y(n_1551) );
INVx1_ASAP7_75t_L g1109 ( .A(n_287), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_288), .A2(n_295), .B1(n_601), .B2(n_1019), .Y(n_1025) );
INVx1_ASAP7_75t_L g1552 ( .A(n_289), .Y(n_1552) );
INVx1_ASAP7_75t_L g1961 ( .A(n_290), .Y(n_1961) );
INVx1_ASAP7_75t_L g1530 ( .A(n_291), .Y(n_1530) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_292), .A2(n_360), .B1(n_784), .B2(n_787), .C(n_788), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_292), .A2(n_360), .B1(n_813), .B2(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g1059 ( .A(n_293), .Y(n_1059) );
OAI211xp5_ASAP7_75t_L g1096 ( .A1(n_293), .A2(n_766), .B(n_846), .C(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g920 ( .A(n_294), .Y(n_920) );
INVx1_ASAP7_75t_L g1482 ( .A(n_296), .Y(n_1482) );
INVx1_ASAP7_75t_L g440 ( .A(n_297), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_298), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g1355 ( .A1(n_299), .A2(n_374), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
INVx1_ASAP7_75t_L g1077 ( .A(n_300), .Y(n_1077) );
INVx1_ASAP7_75t_L g1527 ( .A(n_301), .Y(n_1527) );
INVx1_ASAP7_75t_L g418 ( .A(n_304), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g1212 ( .A(n_305), .Y(n_1212) );
INVx1_ASAP7_75t_L g740 ( .A(n_307), .Y(n_740) );
INVx1_ASAP7_75t_L g1004 ( .A(n_308), .Y(n_1004) );
INVx1_ASAP7_75t_L g1524 ( .A(n_309), .Y(n_1524) );
INVx1_ASAP7_75t_L g424 ( .A(n_310), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_310), .Y(n_431) );
INVx1_ASAP7_75t_L g1665 ( .A(n_311), .Y(n_1665) );
OAI211xp5_ASAP7_75t_L g1670 ( .A1(n_311), .A2(n_1671), .B(n_1673), .C(n_1674), .Y(n_1670) );
INVx1_ASAP7_75t_L g1533 ( .A(n_312), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_314), .Y(n_887) );
INVxp67_ASAP7_75t_SL g641 ( .A(n_315), .Y(n_641) );
INVx1_ASAP7_75t_L g1909 ( .A(n_316), .Y(n_1909) );
INVx1_ASAP7_75t_L g922 ( .A(n_317), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_319), .Y(n_848) );
INVx1_ASAP7_75t_L g1021 ( .A(n_320), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_322), .A2(n_1053), .B1(n_1054), .B2(n_1102), .Y(n_1052) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_322), .Y(n_1102) );
CKINVDCx5p33_ASAP7_75t_R g1207 ( .A(n_323), .Y(n_1207) );
INVx1_ASAP7_75t_L g1692 ( .A(n_324), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_324), .B(n_1691), .Y(n_1697) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_325), .Y(n_859) );
INVx1_ASAP7_75t_L g1191 ( .A(n_326), .Y(n_1191) );
INVx1_ASAP7_75t_L g1901 ( .A(n_327), .Y(n_1901) );
INVx1_ASAP7_75t_L g1478 ( .A(n_328), .Y(n_1478) );
INVx1_ASAP7_75t_L g1322 ( .A(n_329), .Y(n_1322) );
INVx1_ASAP7_75t_L g1260 ( .A(n_330), .Y(n_1260) );
INVx1_ASAP7_75t_L g1917 ( .A(n_331), .Y(n_1917) );
INVx1_ASAP7_75t_L g889 ( .A(n_332), .Y(n_889) );
OAI211xp5_ASAP7_75t_L g898 ( .A1(n_332), .A2(n_513), .B(n_899), .C(n_901), .Y(n_898) );
INVx1_ASAP7_75t_L g1647 ( .A(n_333), .Y(n_1647) );
INVx1_ASAP7_75t_L g1755 ( .A(n_334), .Y(n_1755) );
INVx1_ASAP7_75t_L g1532 ( .A(n_336), .Y(n_1532) );
INVx1_ASAP7_75t_L g460 ( .A(n_337), .Y(n_460) );
INVx1_ASAP7_75t_L g1555 ( .A(n_338), .Y(n_1555) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_339), .A2(n_1339), .B1(n_1395), .B2(n_1396), .Y(n_1338) );
INVxp67_ASAP7_75t_SL g1396 ( .A(n_339), .Y(n_1396) );
INVx1_ASAP7_75t_L g826 ( .A(n_341), .Y(n_826) );
AOI211xp5_ASAP7_75t_SL g1229 ( .A1(n_342), .A2(n_1230), .B(n_1231), .C(n_1233), .Y(n_1229) );
INVx1_ASAP7_75t_L g1417 ( .A(n_343), .Y(n_1417) );
AOI21xp5_ASAP7_75t_SL g1256 ( .A1(n_344), .A2(n_611), .B(n_1023), .Y(n_1256) );
INVx1_ASAP7_75t_L g1268 ( .A(n_344), .Y(n_1268) );
INVx1_ASAP7_75t_L g1605 ( .A(n_345), .Y(n_1605) );
INVx1_ASAP7_75t_L g1321 ( .A(n_347), .Y(n_1321) );
INVxp67_ASAP7_75t_L g1273 ( .A(n_350), .Y(n_1273) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_351), .Y(n_842) );
INVxp67_ASAP7_75t_SL g1286 ( .A(n_352), .Y(n_1286) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g1388 ( .A1(n_354), .A2(n_359), .B1(n_1307), .B2(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1069 ( .A(n_355), .Y(n_1069) );
INVx1_ASAP7_75t_L g1080 ( .A(n_356), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g1148 ( .A(n_358), .Y(n_1148) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_364), .Y(n_644) );
INVx1_ASAP7_75t_L g1488 ( .A(n_365), .Y(n_1488) );
INVx1_ASAP7_75t_L g1525 ( .A(n_366), .Y(n_1525) );
INVx1_ASAP7_75t_L g965 ( .A(n_367), .Y(n_965) );
OAI211xp5_ASAP7_75t_L g972 ( .A1(n_367), .A2(n_973), .B(n_974), .C(n_977), .Y(n_972) );
INVx1_ASAP7_75t_L g413 ( .A(n_368), .Y(n_413) );
INVx1_ASAP7_75t_L g457 ( .A(n_368), .Y(n_457) );
INVx2_ASAP7_75t_L g469 ( .A(n_368), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_370), .Y(n_1149) );
INVx1_ASAP7_75t_L g999 ( .A(n_371), .Y(n_999) );
INVx1_ASAP7_75t_L g781 ( .A(n_372), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_373), .Y(n_1193) );
INVx1_ASAP7_75t_L g1343 ( .A(n_374), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_399), .B(n_1677), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_384), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g1944 ( .A(n_378), .B(n_387), .Y(n_1944) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g1948 ( .A(n_380), .B(n_383), .Y(n_1948) );
INVx1_ASAP7_75t_L g1991 ( .A(n_380), .Y(n_1991) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g1994 ( .A(n_383), .B(n_1991), .Y(n_1994) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g573 ( .A(n_387), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g499 ( .A(n_388), .B(n_398), .Y(n_499) );
AND2x4_ASAP7_75t_L g612 ( .A(n_388), .B(n_397), .Y(n_612) );
INVx1_ASAP7_75t_L g540 ( .A(n_389), .Y(n_540) );
INVx1_ASAP7_75t_L g724 ( .A(n_389), .Y(n_724) );
INVxp67_ASAP7_75t_SL g1353 ( .A(n_389), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1916 ( .A1(n_389), .A2(n_542), .B1(n_1917), .B2(n_1918), .Y(n_1916) );
AND2x4_ASAP7_75t_SL g1943 ( .A(n_389), .B(n_1944), .Y(n_1943) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_396), .Y(n_390) );
OR2x6_ASAP7_75t_L g567 ( .A(n_391), .B(n_543), .Y(n_567) );
INVx1_ASAP7_75t_L g956 ( .A(n_391), .Y(n_956) );
BUFx4f_ASAP7_75t_L g1430 ( .A(n_391), .Y(n_1430) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx4f_ASAP7_75t_L g474 ( .A(n_392), .Y(n_474) );
INVx3_ASAP7_75t_L g791 ( .A(n_392), .Y(n_791) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g480 ( .A(n_394), .Y(n_480) );
INVx2_ASAP7_75t_L g485 ( .A(n_394), .Y(n_485) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_394), .B(n_395), .Y(n_489) );
AND2x2_ASAP7_75t_L g545 ( .A(n_394), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g553 ( .A(n_394), .B(n_395), .Y(n_553) );
INVx1_ASAP7_75t_L g563 ( .A(n_394), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_395), .B(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g484 ( .A(n_395), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g546 ( .A(n_395), .Y(n_546) );
BUFx2_ASAP7_75t_L g558 ( .A(n_395), .Y(n_558) );
INVx1_ASAP7_75t_L g600 ( .A(n_395), .Y(n_600) );
AND2x2_ASAP7_75t_L g602 ( .A(n_395), .B(n_480), .Y(n_602) );
OR2x6_ASAP7_75t_L g1439 ( .A(n_396), .B(n_791), .Y(n_1439) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g551 ( .A(n_397), .Y(n_551) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g557 ( .A(n_398), .Y(n_557) );
AND2x4_ASAP7_75t_L g561 ( .A(n_398), .B(n_562), .Y(n_561) );
XNOR2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_907), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_402), .B1(n_835), .B2(n_836), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AO22x2_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_707), .B1(n_833), .B2(n_834), .Y(n_402) );
INVx1_ASAP7_75t_L g833 ( .A(n_403), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_576), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_501), .C(n_538), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_464), .Y(n_406) );
OAI33xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_417), .A3(n_433), .B1(n_445), .B2(n_451), .B3(n_459), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g727 ( .A1(n_408), .A2(n_728), .A3(n_734), .B1(n_739), .B2(n_742), .B3(n_743), .Y(n_727) );
OAI33xp33_ASAP7_75t_L g915 ( .A1(n_408), .A2(n_665), .A3(n_916), .B1(n_921), .B2(n_928), .B3(n_934), .Y(n_915) );
OAI33xp33_ASAP7_75t_L g1064 ( .A1(n_408), .A2(n_451), .A3(n_1065), .B1(n_1070), .B2(n_1074), .B3(n_1078), .Y(n_1064) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_408), .A2(n_1266), .B1(n_1271), .B2(n_1276), .Y(n_1265) );
OAI33xp33_ASAP7_75t_L g1635 ( .A1(n_408), .A2(n_742), .A3(n_1636), .B1(n_1640), .B2(n_1643), .B3(n_1646), .Y(n_1635) );
OAI33xp33_ASAP7_75t_L g1899 ( .A1(n_408), .A2(n_1900), .A3(n_1903), .B1(n_1906), .B2(n_1910), .B3(n_1912), .Y(n_1899) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx4f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g816 ( .A(n_410), .Y(n_816) );
BUFx8_ASAP7_75t_L g840 ( .A(n_410), .Y(n_840) );
BUFx4f_ASAP7_75t_L g1535 ( .A(n_410), .Y(n_1535) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g498 ( .A(n_411), .Y(n_498) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_411), .Y(n_537) );
OR2x2_ASAP7_75t_L g585 ( .A(n_411), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_SL g1433 ( .A(n_411), .B(n_499), .Y(n_1433) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g575 ( .A(n_412), .Y(n_575) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g1181 ( .A(n_414), .Y(n_1181) );
NAND2xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_416), .Y(n_414) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_415), .Y(n_535) );
INVx1_ASAP7_75t_L g685 ( .A(n_415), .Y(n_685) );
AND3x4_ASAP7_75t_L g1050 ( .A(n_415), .B(n_520), .C(n_634), .Y(n_1050) );
INVx3_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
BUFx3_ASAP7_75t_L g520 ( .A(n_416), .Y(n_520) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_425), .B2(n_426), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_418), .A2(n_460), .B1(n_472), .B2(n_475), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_419), .A2(n_460), .B1(n_461), .B2(n_463), .Y(n_459) );
OR2x6_ASAP7_75t_L g807 ( .A(n_419), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_419), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g1563 ( .A1(n_419), .A2(n_649), .B1(n_1551), .B2(n_1557), .Y(n_1563) );
OAI22xp33_ASAP7_75t_L g1567 ( .A1(n_419), .A2(n_962), .B1(n_1552), .B2(n_1558), .Y(n_1567) );
OAI22xp33_ASAP7_75t_L g1912 ( .A1(n_419), .A2(n_649), .B1(n_1913), .B2(n_1914), .Y(n_1912) );
INVx2_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g1042 ( .A(n_420), .Y(n_1042) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x4_ASAP7_75t_L g505 ( .A(n_421), .B(n_455), .Y(n_505) );
OR2x4_ASAP7_75t_L g529 ( .A(n_421), .B(n_508), .Y(n_529) );
BUFx3_ASAP7_75t_L g647 ( .A(n_421), .Y(n_647) );
BUFx3_ASAP7_75t_L g730 ( .A(n_421), .Y(n_730) );
BUFx4f_ASAP7_75t_L g919 ( .A(n_421), .Y(n_919) );
OR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_422), .Y(n_432) );
INVx2_ASAP7_75t_L g439 ( .A(n_422), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_422), .B(n_431), .Y(n_444) );
AND2x4_ASAP7_75t_L g515 ( .A(n_422), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g662 ( .A(n_423), .Y(n_662) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g438 ( .A(n_424), .Y(n_438) );
OAI22xp33_ASAP7_75t_SL g490 ( .A1(n_425), .A2(n_463), .B1(n_491), .B2(n_492), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_426), .A2(n_919), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
OAI211xp5_ASAP7_75t_L g1179 ( .A1(n_426), .A2(n_1134), .B(n_1180), .C(n_1182), .Y(n_1179) );
OAI22xp33_ASAP7_75t_L g1491 ( .A1(n_426), .A2(n_1042), .B1(n_1478), .B2(n_1485), .Y(n_1491) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g962 ( .A(n_427), .Y(n_962) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
INVx4_ASAP7_75t_L g512 ( .A(n_428), .Y(n_512) );
OR2x2_ASAP7_75t_L g584 ( .A(n_428), .B(n_585), .Y(n_584) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g650 ( .A(n_429), .Y(n_650) );
BUFx2_ASAP7_75t_L g862 ( .A(n_429), .Y(n_862) );
NAND2x1p5_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
BUFx2_ASAP7_75t_L g524 ( .A(n_430), .Y(n_524) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g516 ( .A(n_431), .Y(n_516) );
BUFx2_ASAP7_75t_L g521 ( .A(n_432), .Y(n_521) );
INVx2_ASAP7_75t_L g687 ( .A(n_432), .Y(n_687) );
AND2x4_ASAP7_75t_L g1038 ( .A(n_432), .B(n_693), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_440), .B2(n_441), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_446), .B1(n_482), .B2(n_486), .Y(n_481) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g669 ( .A(n_436), .Y(n_669) );
INVx1_ASAP7_75t_L g822 ( .A(n_436), .Y(n_822) );
BUFx2_ASAP7_75t_L g1386 ( .A(n_436), .Y(n_1386) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx8_ASAP7_75t_L g448 ( .A(n_437), .Y(n_448) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_437), .Y(n_509) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_437), .Y(n_640) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x4_ASAP7_75t_L g661 ( .A(n_439), .B(n_662), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_440), .A2(n_449), .B1(n_472), .B2(n_475), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_441), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_441), .A2(n_935), .B1(n_936), .B2(n_937), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g1600 ( .A1(n_441), .A2(n_745), .B1(n_1601), .B2(n_1602), .Y(n_1600) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g450 ( .A(n_442), .Y(n_450) );
CKINVDCx8_ASAP7_75t_R g642 ( .A(n_442), .Y(n_642) );
INVx1_ASAP7_75t_L g655 ( .A(n_442), .Y(n_655) );
INVx3_ASAP7_75t_L g1418 ( .A(n_442), .Y(n_1418) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g676 ( .A(n_443), .Y(n_676) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g532 ( .A(n_444), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_449), .B2(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g1045 ( .A(n_447), .Y(n_1045) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g810 ( .A(n_448), .B(n_705), .Y(n_810) );
INVx3_ASAP7_75t_L g1075 ( .A(n_448), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1416 ( .A(n_448), .Y(n_1416) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_450), .A2(n_824), .B1(n_825), .B2(n_826), .C(n_827), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_450), .A2(n_1071), .B1(n_1072), .B2(n_1073), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_450), .A2(n_1075), .B1(n_1076), .B2(n_1077), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_450), .A2(n_929), .B1(n_1524), .B2(n_1532), .Y(n_1539) );
OAI22xp5_ASAP7_75t_L g1903 ( .A1(n_450), .A2(n_1565), .B1(n_1904), .B2(n_1905), .Y(n_1903) );
OAI22xp5_ASAP7_75t_SL g815 ( .A1(n_451), .A2(n_816), .B1(n_817), .B2(n_823), .Y(n_815) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g1911 ( .A(n_453), .Y(n_1911) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g666 ( .A(n_454), .Y(n_666) );
NAND3x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .C(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g508 ( .A(n_455), .Y(n_508) );
AND2x4_ASAP7_75t_L g514 ( .A(n_455), .B(n_515), .Y(n_514) );
OR2x6_ASAP7_75t_L g531 ( .A(n_455), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g684 ( .A(n_455), .B(n_685), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g1175 ( .A(n_455), .B(n_458), .Y(n_1175) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g678 ( .A(n_457), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_457), .B(n_605), .Y(n_1117) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_461), .A2(n_730), .B1(n_740), .B2(n_741), .Y(n_739) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g932 ( .A(n_462), .Y(n_932) );
HB1xp67_ASAP7_75t_L g1596 ( .A(n_462), .Y(n_1596) );
OAI22xp33_ASAP7_75t_L g1900 ( .A1(n_462), .A2(n_1544), .B1(n_1901), .B2(n_1902), .Y(n_1900) );
OAI22xp33_ASAP7_75t_L g1965 ( .A1(n_462), .A2(n_1042), .B1(n_1966), .B2(n_1967), .Y(n_1965) );
OAI33xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_471), .A3(n_481), .B1(n_490), .B2(n_494), .B3(n_500), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_465), .A2(n_748), .B1(n_751), .B2(n_753), .Y(n_747) );
OAI33xp33_ASAP7_75t_L g864 ( .A1(n_465), .A2(n_753), .A3(n_865), .B1(n_868), .B2(n_871), .B3(n_875), .Y(n_864) );
OAI33xp33_ASAP7_75t_L g1606 ( .A1(n_465), .A2(n_958), .A3(n_1607), .B1(n_1609), .B2(n_1610), .B3(n_1612), .Y(n_1606) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g939 ( .A(n_467), .Y(n_939) );
INVx1_ASAP7_75t_L g1082 ( .A(n_467), .Y(n_1082) );
INVx4_ASAP7_75t_L g1374 ( .A(n_467), .Y(n_1374) );
INVx2_ASAP7_75t_L g1480 ( .A(n_467), .Y(n_1480) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g801 ( .A(n_468), .Y(n_801) );
OR2x6_ASAP7_75t_L g1205 ( .A(n_468), .B(n_1175), .Y(n_1205) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g634 ( .A(n_469), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_469), .B(n_583), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_472), .A2(n_917), .B1(n_936), .B2(n_941), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g1550 ( .A1(n_472), .A2(n_941), .B1(n_1551), .B2(n_1552), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1559 ( .A1(n_472), .A2(n_475), .B1(n_1560), .B2(n_1561), .Y(n_1559) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g1086 ( .A(n_474), .Y(n_1086) );
INVx4_ASAP7_75t_L g1235 ( .A(n_474), .Y(n_1235) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g795 ( .A(n_477), .Y(n_795) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_477), .Y(n_867) );
INVx2_ASAP7_75t_L g876 ( .A(n_477), .Y(n_876) );
INVx2_ASAP7_75t_SL g943 ( .A(n_477), .Y(n_943) );
INVx2_ASAP7_75t_L g1129 ( .A(n_477), .Y(n_1129) );
INVx2_ASAP7_75t_L g1326 ( .A(n_477), .Y(n_1326) );
INVx1_ASAP7_75t_L g1651 ( .A(n_477), .Y(n_1651) );
INVx8_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_557), .Y(n_571) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_478), .Y(n_1431) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI221xp5_ASAP7_75t_SL g748 ( .A1(n_482), .A2(n_548), .B1(n_735), .B2(n_744), .C(n_749), .Y(n_748) );
OAI221xp5_ASAP7_75t_SL g751 ( .A1(n_482), .A2(n_548), .B1(n_731), .B2(n_741), .C(n_752), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_482), .A2(n_612), .B1(n_874), .B2(n_1217), .C(n_1218), .Y(n_1216) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g491 ( .A(n_483), .Y(n_491) );
BUFx2_ASAP7_75t_L g873 ( .A(n_483), .Y(n_873) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g870 ( .A(n_484), .Y(n_870) );
BUFx2_ASAP7_75t_L g947 ( .A(n_484), .Y(n_947) );
BUFx3_ASAP7_75t_L g951 ( .A(n_484), .Y(n_951) );
BUFx2_ASAP7_75t_L g1425 ( .A(n_484), .Y(n_1425) );
AND2x2_ASAP7_75t_L g599 ( .A(n_485), .B(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_485), .Y(n_1012) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g874 ( .A(n_487), .Y(n_874) );
INVx1_ASAP7_75t_L g957 ( .A(n_487), .Y(n_957) );
INVx1_ASAP7_75t_L g1007 ( .A(n_487), .Y(n_1007) );
INVx2_ASAP7_75t_L g1436 ( .A(n_487), .Y(n_1436) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_488), .Y(n_493) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
BUFx4f_ASAP7_75t_L g1088 ( .A(n_488), .Y(n_1088) );
BUFx4f_ASAP7_75t_L g1135 ( .A(n_488), .Y(n_1135) );
OR2x6_ASAP7_75t_L g1139 ( .A(n_488), .B(n_1140), .Y(n_1139) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_488), .A2(n_499), .B1(n_951), .B2(n_1333), .C(n_1334), .Y(n_1332) );
BUFx4f_ASAP7_75t_L g1426 ( .A(n_488), .Y(n_1426) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g884 ( .A(n_489), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_491), .A2(n_1071), .B1(n_1076), .B2(n_1088), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_491), .A2(n_1069), .B1(n_1080), .B2(n_1088), .Y(n_1089) );
OAI221xp5_ASAP7_75t_L g1320 ( .A1(n_491), .A2(n_612), .B1(n_874), .B2(n_1321), .C(n_1322), .Y(n_1320) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_491), .A2(n_1088), .B1(n_1524), .B2(n_1525), .Y(n_1523) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_491), .A2(n_1527), .B1(n_1528), .B2(n_1530), .Y(n_1526) );
OAI221xp5_ASAP7_75t_L g1929 ( .A1(n_491), .A2(n_883), .B1(n_1904), .B2(n_1907), .C(n_1930), .Y(n_1929) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g868 ( .A1(n_493), .A2(n_848), .B1(n_854), .B2(n_869), .Y(n_868) );
OAI33xp33_ASAP7_75t_L g1081 ( .A1(n_494), .A2(n_1082), .A3(n_1083), .B1(n_1087), .B2(n_1089), .B3(n_1090), .Y(n_1081) );
OAI33xp33_ASAP7_75t_L g1517 ( .A1(n_494), .A2(n_1480), .A3(n_1518), .B1(n_1523), .B2(n_1526), .B3(n_1531), .Y(n_1517) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI33xp33_ASAP7_75t_L g1549 ( .A1(n_496), .A2(n_1374), .A3(n_1550), .B1(n_1553), .B2(n_1556), .B3(n_1559), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
AND2x4_ASAP7_75t_L g754 ( .A(n_497), .B(n_499), .Y(n_754) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_SL g595 ( .A(n_499), .Y(n_595) );
INVx4_ASAP7_75t_L g1024 ( .A(n_499), .Y(n_1024) );
OAI21xp33_ASAP7_75t_L g1231 ( .A1(n_499), .A2(n_951), .B(n_1232), .Y(n_1231) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_510), .A3(n_526), .B(n_533), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g897 ( .A(n_505), .Y(n_897) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_505), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1623 ( .A(n_505), .Y(n_1623) );
INVx1_ASAP7_75t_L g1660 ( .A(n_505), .Y(n_1660) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g768 ( .A(n_507), .Y(n_768) );
INVx2_ASAP7_75t_L g1095 ( .A(n_507), .Y(n_1095) );
INVxp67_ASAP7_75t_L g1356 ( .A(n_507), .Y(n_1356) );
INVx1_ASAP7_75t_L g1450 ( .A(n_507), .Y(n_1450) );
INVx1_ASAP7_75t_L g1510 ( .A(n_507), .Y(n_1510) );
AOI22xp33_ASAP7_75t_L g1940 ( .A1(n_507), .A2(n_1094), .B1(n_1917), .B2(n_1918), .Y(n_1940) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_509), .Y(n_653) );
INVx2_ASAP7_75t_L g736 ( .A(n_509), .Y(n_736) );
INVx1_ASAP7_75t_L g745 ( .A(n_509), .Y(n_745) );
BUFx6f_ASAP7_75t_L g1197 ( .A(n_509), .Y(n_1197) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g900 ( .A(n_512), .Y(n_900) );
INVx2_ASAP7_75t_L g1043 ( .A(n_512), .Y(n_1043) );
INVx2_ASAP7_75t_L g1173 ( .A(n_512), .Y(n_1173) );
CKINVDCx8_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
CKINVDCx8_ASAP7_75t_R g766 ( .A(n_514), .Y(n_766) );
OAI31xp33_ASAP7_75t_L g1277 ( .A1(n_514), .A2(n_1278), .A3(n_1288), .B(n_1290), .Y(n_1277) );
AOI211xp5_ASAP7_75t_L g1935 ( .A1(n_514), .A2(n_829), .B(n_1936), .C(n_1937), .Y(n_1935) );
INVx2_ASAP7_75t_L g664 ( .A(n_515), .Y(n_664) );
BUFx2_ASAP7_75t_L g695 ( .A(n_515), .Y(n_695) );
BUFx2_ASAP7_75t_L g763 ( .A(n_515), .Y(n_763) );
BUFx2_ASAP7_75t_L g821 ( .A(n_515), .Y(n_821) );
BUFx3_ASAP7_75t_L g829 ( .A(n_515), .Y(n_829) );
BUFx2_ASAP7_75t_L g1167 ( .A(n_515), .Y(n_1167) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_515), .Y(n_1275) );
INVx1_ASAP7_75t_L g693 ( .A(n_516), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_522), .B1(n_523), .B2(n_525), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_518), .A2(n_523), .B1(n_887), .B2(n_902), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_518), .A2(n_523), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g1285 ( .A1(n_518), .A2(n_523), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
AOI22xp33_ASAP7_75t_SL g1455 ( .A1(n_518), .A2(n_523), .B1(n_1444), .B2(n_1456), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_518), .A2(n_523), .B1(n_1463), .B2(n_1473), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_518), .A2(n_523), .B1(n_1573), .B2(n_1574), .Y(n_1572) );
INVx1_ASAP7_75t_L g1938 ( .A(n_518), .Y(n_1938) );
AOI22xp33_ASAP7_75t_L g1985 ( .A1(n_518), .A2(n_523), .B1(n_1978), .B2(n_1986), .Y(n_1985) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
AND2x4_ASAP7_75t_L g523 ( .A(n_519), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g759 ( .A(n_519), .B(n_521), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g1278 ( .A1(n_519), .A2(n_1279), .B(n_1282), .C(n_1285), .Y(n_1278) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_522), .A2(n_555), .B1(n_559), .B2(n_564), .Y(n_554) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_523), .Y(n_760) );
INVx1_ASAP7_75t_L g1939 ( .A(n_523), .Y(n_1939) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_528), .A2(n_713), .B1(n_715), .B2(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g1101 ( .A(n_528), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1941 ( .A1(n_528), .A2(n_765), .B1(n_1926), .B2(n_1927), .Y(n_1941) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_529), .Y(n_1289) );
BUFx3_ASAP7_75t_L g1361 ( .A(n_529), .Y(n_1361) );
BUFx2_ASAP7_75t_L g1628 ( .A(n_529), .Y(n_1628) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g765 ( .A(n_531), .Y(n_765) );
INVx1_ASAP7_75t_L g905 ( .A(n_531), .Y(n_905) );
INVx1_ASAP7_75t_L g1453 ( .A(n_531), .Y(n_1453) );
BUFx3_ASAP7_75t_L g738 ( .A(n_532), .Y(n_738) );
INVx1_ASAP7_75t_L g852 ( .A(n_532), .Y(n_852) );
OAI21xp33_ASAP7_75t_L g755 ( .A1(n_533), .A2(n_756), .B(n_767), .Y(n_755) );
OAI31xp33_ASAP7_75t_SL g959 ( .A1(n_533), .A2(n_960), .A3(n_961), .B(n_966), .Y(n_959) );
OAI31xp33_ASAP7_75t_L g1091 ( .A1(n_533), .A2(n_1092), .A3(n_1096), .B(n_1100), .Y(n_1091) );
OAI31xp33_ASAP7_75t_L g1621 ( .A1(n_533), .A2(n_1622), .A3(n_1624), .B(n_1627), .Y(n_1621) );
AND2x2_ASAP7_75t_SL g533 ( .A(n_534), .B(n_536), .Y(n_533) );
AND2x4_ASAP7_75t_L g906 ( .A(n_534), .B(n_536), .Y(n_906) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_534), .B(n_536), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_534), .B(n_536), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_534), .B(n_536), .Y(n_1667) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI31xp33_ASAP7_75t_SL g538 ( .A1(n_539), .A2(n_547), .A3(n_565), .B(n_572), .Y(n_538) );
INVx3_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g879 ( .A(n_542), .Y(n_879) );
INVx4_ASAP7_75t_L g1615 ( .A(n_542), .Y(n_1615) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
BUFx3_ASAP7_75t_L g610 ( .A(n_545), .Y(n_610) );
INVx2_ASAP7_75t_L g777 ( .A(n_545), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_548), .A2(n_922), .B1(n_930), .B2(n_945), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_548), .A2(n_945), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_549), .B(n_712), .C(n_716), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g1341 ( .A(n_549), .B(n_1342), .C(n_1348), .Y(n_1341) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g977 ( .A(n_550), .Y(n_977) );
INVx1_ASAP7_75t_L g1673 ( .A(n_550), .Y(n_1673) );
AOI211xp5_ASAP7_75t_L g1919 ( .A1(n_550), .A2(n_1920), .B(n_1922), .C(n_1923), .Y(n_1919) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_551), .B(n_1371), .Y(n_1442) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_552), .Y(n_591) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_552), .B(n_605), .Y(n_604) );
AND2x6_ASAP7_75t_L g607 ( .A(n_552), .B(n_583), .Y(n_607) );
BUFx3_ASAP7_75t_L g718 ( .A(n_552), .Y(n_718) );
BUFx3_ASAP7_75t_L g798 ( .A(n_552), .Y(n_798) );
BUFx3_ASAP7_75t_L g1230 ( .A(n_552), .Y(n_1230) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g1372 ( .A(n_553), .Y(n_1372) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_555), .A2(n_717), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_721), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_555), .A2(n_964), .B1(n_975), .B2(n_976), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_555), .A2(n_975), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_555), .A2(n_975), .B1(n_1506), .B2(n_1507), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1578 ( .A1(n_555), .A2(n_975), .B1(n_1573), .B2(n_1579), .Y(n_1578) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_556), .A2(n_561), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
INVx1_ASAP7_75t_L g1924 ( .A(n_556), .Y(n_1924) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g714 ( .A(n_557), .B(n_616), .Y(n_714) );
AND2x2_ASAP7_75t_L g886 ( .A(n_557), .B(n_558), .Y(n_886) );
INVx1_ASAP7_75t_L g624 ( .A(n_558), .Y(n_624) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_558), .Y(n_1009) );
INVx1_ASAP7_75t_L g1146 ( .A(n_558), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_558), .A2(n_1011), .B1(n_1189), .B2(n_1210), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_559), .A2(n_886), .B1(n_1664), .B2(n_1675), .Y(n_1674) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g722 ( .A(n_561), .Y(n_722) );
BUFx3_ASAP7_75t_L g975 ( .A(n_561), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_562), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_L g891 ( .A(n_567), .Y(n_891) );
INVx1_ASAP7_75t_L g971 ( .A(n_567), .Y(n_971) );
BUFx6f_ASAP7_75t_L g1447 ( .A(n_567), .Y(n_1447) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_569), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g1581 ( .A(n_570), .Y(n_1581) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g893 ( .A(n_571), .Y(n_893) );
INVx1_ASAP7_75t_L g1346 ( .A(n_571), .Y(n_1346) );
OAI31xp33_ASAP7_75t_L g877 ( .A1(n_572), .A2(n_878), .A3(n_880), .B(n_890), .Y(n_877) );
OAI31xp33_ASAP7_75t_L g1613 ( .A1(n_572), .A2(n_1614), .A3(n_1616), .B(n_1620), .Y(n_1613) );
OAI31xp33_ASAP7_75t_L g1668 ( .A1(n_572), .A2(n_1669), .A3(n_1670), .B(n_1676), .Y(n_1668) );
BUFx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g725 ( .A(n_573), .Y(n_725) );
BUFx2_ASAP7_75t_SL g978 ( .A(n_573), .Y(n_978) );
OAI31xp33_ASAP7_75t_L g1055 ( .A1(n_573), .A2(n_1056), .A3(n_1060), .B(n_1061), .Y(n_1055) );
INVx1_ASAP7_75t_L g1499 ( .A(n_573), .Y(n_1499) );
OAI31xp33_ASAP7_75t_L g1975 ( .A1(n_573), .A2(n_1976), .A3(n_1980), .B(n_1981), .Y(n_1975) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g581 ( .A(n_575), .B(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g700 ( .A(n_575), .Y(n_700) );
INVx1_ASAP7_75t_L g989 ( .A(n_575), .Y(n_989) );
XNOR2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_706), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_578), .B(n_671), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_587), .B1(n_588), .B2(n_632), .C(n_635), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
AND2x4_ASAP7_75t_L g805 ( .A(n_581), .B(n_584), .Y(n_805) );
INVx1_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_583), .B(n_599), .Y(n_679) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_583), .Y(n_1013) );
INVx2_ASAP7_75t_L g1188 ( .A(n_584), .Y(n_1188) );
INVx1_ASAP7_75t_L g670 ( .A(n_585), .Y(n_670) );
OR2x2_ASAP7_75t_L g675 ( .A(n_585), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g705 ( .A(n_585), .Y(n_705) );
INVx1_ASAP7_75t_L g1170 ( .A(n_586), .Y(n_1170) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_608), .C(n_626), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_596), .B1(n_603), .B2(n_606), .C(n_607), .Y(n_589) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_591), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1222 ( .A1(n_591), .A2(n_1207), .B1(n_1212), .B2(n_1223), .C(n_1225), .Y(n_1222) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_591), .A2(n_1223), .B1(n_1300), .B2(n_1313), .C(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1921 ( .A(n_591), .Y(n_1921) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g627 ( .A(n_594), .B(n_605), .Y(n_627) );
AND2x2_ASAP7_75t_L g994 ( .A(n_594), .B(n_605), .Y(n_994) );
BUFx6f_ASAP7_75t_L g1023 ( .A(n_594), .Y(n_1023) );
INVx2_ASAP7_75t_L g1224 ( .A(n_594), .Y(n_1224) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g1019 ( .A(n_598), .Y(n_1019) );
INVx2_ASAP7_75t_L g1138 ( .A(n_598), .Y(n_1138) );
INVx1_ASAP7_75t_L g1368 ( .A(n_598), .Y(n_1368) );
INVx2_ASAP7_75t_L g1931 ( .A(n_598), .Y(n_1931) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_599), .Y(n_616) );
AND2x2_ASAP7_75t_L g619 ( .A(n_599), .B(n_605), .Y(n_619) );
BUFx3_ASAP7_75t_L g1366 ( .A(n_601), .Y(n_1366) );
BUFx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx3_ASAP7_75t_L g617 ( .A(n_602), .Y(n_617) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_602), .Y(n_630) );
INVx2_ASAP7_75t_L g1030 ( .A(n_602), .Y(n_1030) );
BUFx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g786 ( .A(n_604), .Y(n_786) );
AND2x4_ASAP7_75t_L g629 ( .A(n_605), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_605), .B(n_1029), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_605), .Y(n_1221) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_606), .A2(n_682), .B1(n_688), .B2(n_689), .C(n_694), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_607), .A2(n_775), .B(n_778), .Y(n_774) );
AOI221xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_613), .B1(n_618), .B2(n_620), .C(n_621), .Y(n_608) );
BUFx2_ASAP7_75t_L g1365 ( .A(n_610), .Y(n_1365) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g1017 ( .A(n_612), .Y(n_1017) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g1215 ( .A(n_615), .Y(n_1215) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_616), .Y(n_1005) );
A2O1A1Ixp33_ASAP7_75t_L g1226 ( .A1(n_616), .A2(n_1013), .B(n_1193), .C(n_1227), .Y(n_1226) );
A2O1A1Ixp33_ASAP7_75t_L g1327 ( .A1(n_616), .A2(n_1304), .B(n_1328), .C(n_1330), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_618), .A2(n_627), .B1(n_781), .B2(n_782), .Y(n_780) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g988 ( .A(n_619), .B(n_989), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_620), .B(n_702), .Y(n_701) );
BUFx2_ASAP7_75t_L g787 ( .A(n_622), .Y(n_787) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g1263 ( .A(n_624), .Y(n_1263) );
INVx1_ASAP7_75t_L g1330 ( .A(n_625), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_629), .B2(n_631), .Y(n_626) );
INVx3_ASAP7_75t_L g773 ( .A(n_629), .Y(n_773) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_630), .Y(n_750) );
BUFx2_ASAP7_75t_L g779 ( .A(n_630), .Y(n_779) );
INVx1_ASAP7_75t_L g1319 ( .A(n_630), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_631), .B(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_633), .Y(n_1033) );
OAI31xp33_ASAP7_75t_L g1213 ( .A1(n_633), .A2(n_1214), .A3(n_1219), .B(n_1229), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1245 ( .A(n_633), .Y(n_1245) );
OAI31xp33_ASAP7_75t_L g1316 ( .A1(n_633), .A2(n_1317), .A3(n_1323), .B(n_1331), .Y(n_1316) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_641), .B2(n_642), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_638), .A2(n_642), .B1(n_854), .B2(n_855), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g1646 ( .A1(n_638), .A2(n_738), .B1(n_1647), .B2(n_1648), .Y(n_1646) );
BUFx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx8_ASAP7_75t_L g1036 ( .A(n_639), .Y(n_1036) );
INVx5_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g925 ( .A(n_640), .Y(n_925) );
INVx2_ASAP7_75t_SL g1200 ( .A(n_640), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_640), .A2(n_828), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g1542 ( .A(n_640), .Y(n_1542) );
INVx2_ASAP7_75t_SL g1565 ( .A(n_640), .Y(n_1565) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_642), .A2(n_652), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1266 ( .A1(n_642), .A2(n_1267), .B1(n_1268), .B2(n_1269), .C(n_1270), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_642), .A2(n_1255), .B1(n_1272), .B2(n_1273), .C(n_1274), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g1597 ( .A1(n_642), .A2(n_1565), .B1(n_1598), .B2(n_1599), .Y(n_1597) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_648), .B2(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g844 ( .A(n_647), .Y(n_844) );
INVx1_ASAP7_75t_L g858 ( .A(n_647), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_649), .A2(n_917), .B1(n_918), .B2(n_920), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g1543 ( .A1(n_649), .A2(n_1522), .B1(n_1530), .B2(n_1544), .Y(n_1543) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g733 ( .A(n_650), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g1494 ( .A1(n_650), .A2(n_1042), .B1(n_1479), .B2(n_1486), .Y(n_1494) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_SL g1267 ( .A(n_653), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_655), .A2(n_1386), .B1(n_1412), .B2(n_1413), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_655), .A2(n_1386), .B1(n_1482), .B2(n_1488), .Y(n_1492) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g819 ( .A(n_660), .Y(n_819) );
BUFx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g699 ( .A(n_661), .B(n_684), .Y(n_699) );
INVx8_ASAP7_75t_L g704 ( .A(n_661), .Y(n_704) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_661), .Y(n_1163) );
BUFx3_ASAP7_75t_L g1297 ( .A(n_661), .Y(n_1297) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1203 ( .A(n_664), .Y(n_1203) );
INVx1_ASAP7_75t_L g1298 ( .A(n_664), .Y(n_1298) );
OAI33xp33_ASAP7_75t_L g1534 ( .A1(n_665), .A2(n_1535), .A3(n_1536), .B1(n_1539), .B2(n_1540), .B3(n_1543), .Y(n_1534) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_666), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_666), .A2(n_694), .B1(n_1035), .B2(n_1044), .C(n_1049), .Y(n_1034) );
INVx2_ASAP7_75t_L g1276 ( .A(n_666), .Y(n_1276) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_666), .B(n_1391), .C(n_1394), .Y(n_1390) );
NAND2x1_ASAP7_75t_L g991 ( .A(n_667), .B(n_992), .Y(n_991) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g1272 ( .A(n_669), .Y(n_1272) );
INVxp67_ASAP7_75t_L g808 ( .A(n_670), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_680), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_673), .A2(n_831), .B(n_832), .Y(n_830) );
INVx8_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g1192 ( .A(n_675), .Y(n_1192) );
BUFx3_ASAP7_75t_L g1908 ( .A(n_676), .Y(n_1908) );
INVx1_ASAP7_75t_L g1113 ( .A(n_677), .Y(n_1113) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
AND2x4_ASAP7_75t_L g683 ( .A(n_678), .B(n_684), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_696), .C(n_701), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g1209 ( .A1(n_682), .A2(n_694), .B1(n_1210), .B2(n_1211), .C(n_1212), .Y(n_1209) );
AOI221xp5_ASAP7_75t_L g1311 ( .A1(n_682), .A2(n_694), .B1(n_1211), .B2(n_1312), .C(n_1313), .Y(n_1311) );
AND2x4_ASAP7_75t_SL g682 ( .A(n_683), .B(n_686), .Y(n_682) );
AND2x4_ASAP7_75t_L g689 ( .A(n_683), .B(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g694 ( .A(n_683), .B(n_695), .Y(n_694) );
NAND2x1_ASAP7_75t_L g813 ( .A(n_683), .B(n_686), .Y(n_813) );
AND2x4_ASAP7_75t_SL g1211 ( .A(n_683), .B(n_690), .Y(n_1211) );
AND2x6_ASAP7_75t_L g1153 ( .A(n_684), .B(n_686), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_684), .B(n_692), .Y(n_1155) );
INVx1_ASAP7_75t_L g1160 ( .A(n_684), .Y(n_1160) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g814 ( .A(n_689), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_689), .A2(n_997), .B1(n_998), .B2(n_999), .C(n_1000), .Y(n_996) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_694), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_697), .B(n_1238), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_697), .B(n_1315), .Y(n_1314) );
INVx5_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x6_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
AND2x4_ASAP7_75t_L g1190 ( .A(n_703), .B(n_705), .Y(n_1190) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx8_ASAP7_75t_L g828 ( .A(n_704), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g1158 ( .A(n_704), .Y(n_1158) );
INVx3_ASAP7_75t_L g1183 ( .A(n_704), .Y(n_1183) );
INVx1_ASAP7_75t_L g834 ( .A(n_707), .Y(n_834) );
XNOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_770), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_769), .Y(n_708) );
NAND3x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_726), .C(n_755), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_723), .B(n_725), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g1342 ( .A1(n_714), .A2(n_1343), .B1(n_1344), .B2(n_1347), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1925 ( .A1(n_714), .A2(n_1344), .B1(n_1926), .B2(n_1927), .Y(n_1925) );
AOI222xp33_ASAP7_75t_L g757 ( .A1(n_717), .A2(n_719), .B1(n_720), .B2(n_758), .C1(n_760), .C2(n_761), .Y(n_757) );
AOI222xp33_ASAP7_75t_L g1348 ( .A1(n_718), .A2(n_721), .B1(n_886), .B2(n_1349), .C1(n_1350), .C2(n_1351), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_721), .A2(n_886), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1977 ( .A1(n_721), .A2(n_886), .B1(n_1978), .B2(n_1979), .Y(n_1977) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g888 ( .A(n_722), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g1340 ( .A1(n_725), .A2(n_1341), .B(n_1352), .Y(n_1340) );
OAI31xp33_ASAP7_75t_L g1437 ( .A1(n_725), .A2(n_1438), .A3(n_1440), .B(n_1446), .Y(n_1437) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_747), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g1172 ( .A1(n_730), .A2(n_1130), .B1(n_1136), .B2(n_1173), .C(n_1174), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g1419 ( .A1(n_730), .A2(n_1420), .B1(n_1421), .B2(n_1422), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g1593 ( .A1(n_730), .A2(n_1594), .B1(n_1595), .B2(n_1596), .Y(n_1593) );
OAI22xp33_ASAP7_75t_L g1643 ( .A1(n_730), .A2(n_846), .B1(n_1644), .B2(n_1645), .Y(n_1643) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g846 ( .A(n_733), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1564 ( .A1(n_738), .A2(n_1554), .B1(n_1560), .B2(n_1565), .Y(n_1564) );
OAI33xp33_ASAP7_75t_L g839 ( .A1(n_742), .A2(n_840), .A3(n_841), .B1(n_847), .B2(n_853), .B3(n_856), .Y(n_839) );
OAI33xp33_ASAP7_75t_L g1592 ( .A1(n_742), .A2(n_1535), .A3(n_1593), .B1(n_1597), .B2(n_1600), .B3(n_1603), .Y(n_1592) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_745), .A2(n_848), .B1(n_849), .B2(n_850), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g1132 ( .A1(n_753), .A2(n_1133), .B(n_1139), .Y(n_1132) );
OAI22xp5_ASAP7_75t_SL g1928 ( .A1(n_753), .A2(n_939), .B1(n_1929), .B2(n_1932), .Y(n_1928) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g958 ( .A(n_754), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g1375 ( .A(n_754), .B(n_1376), .C(n_1382), .Y(n_1375) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_764), .C(n_766), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g1663 ( .A1(n_758), .A2(n_760), .B1(n_1664), .B2(n_1665), .Y(n_1663) );
BUFx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx3_ASAP7_75t_L g1098 ( .A(n_759), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_760), .A2(n_1058), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_760), .A2(n_1098), .B1(n_1350), .B2(n_1351), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_760), .A2(n_1098), .B1(n_1506), .B2(n_1513), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1625 ( .A1(n_760), .A2(n_1098), .B1(n_1618), .B2(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g1357 ( .A(n_765), .Y(n_1357) );
O2A1O1Ixp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_783), .B(n_799), .C(n_802), .Y(n_771) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g1123 ( .A(n_777), .Y(n_1123) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g1031 ( .A(n_785), .Y(n_1031) );
INVx4_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_792), .B1(n_793), .B2(n_796), .C(n_797), .Y(n_788) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_789), .A2(n_842), .B1(n_859), .B2(n_866), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_789), .A2(n_849), .B1(n_855), .B2(n_876), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g1971 ( .A1(n_789), .A2(n_795), .B1(n_1956), .B2(n_1966), .Y(n_1971) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
BUFx3_ASAP7_75t_L g1127 ( .A(n_791), .Y(n_1127) );
BUFx6f_ASAP7_75t_L g1428 ( .A(n_791), .Y(n_1428) );
BUFx3_ASAP7_75t_L g1656 ( .A(n_791), .Y(n_1656) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_792), .A2(n_818), .B(n_820), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_793), .A2(n_1066), .B1(n_1079), .B2(n_1084), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_793), .A2(n_1073), .B1(n_1077), .B2(n_1084), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1518 ( .A1(n_793), .A2(n_1519), .B1(n_1520), .B2(n_1522), .Y(n_1518) );
OAI22xp5_ASAP7_75t_L g1531 ( .A1(n_793), .A2(n_1520), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_795), .A2(n_1234), .B1(n_1235), .B2(n_1236), .Y(n_1233) );
OAI22xp33_ASAP7_75t_L g1427 ( .A1(n_795), .A2(n_1407), .B1(n_1420), .B2(n_1428), .Y(n_1427) );
OAI22xp33_ASAP7_75t_L g1477 ( .A1(n_795), .A2(n_1428), .B1(n_1478), .B2(n_1479), .Y(n_1477) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI31xp67_ASAP7_75t_L g1150 ( .A1(n_800), .A2(n_1151), .A3(n_1161), .B(n_1171), .Y(n_1150) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_811), .C(n_830), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_807), .B(n_987), .Y(n_986) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_810), .B(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_810), .B(n_1300), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_815), .Y(n_811) );
INVx2_ASAP7_75t_L g997 ( .A(n_813), .Y(n_997) );
OAI33xp33_ASAP7_75t_L g1405 ( .A1(n_816), .A2(n_1205), .A3(n_1406), .B1(n_1411), .B2(n_1414), .B3(n_1419), .Y(n_1405) );
OAI33xp33_ASAP7_75t_L g1490 ( .A1(n_816), .A2(n_1205), .A3(n_1491), .B1(n_1492), .B2(n_1493), .B3(n_1494), .Y(n_1490) );
OAI33xp33_ASAP7_75t_L g1954 ( .A1(n_816), .A2(n_1205), .A3(n_1955), .B1(n_1959), .B2(n_1962), .B3(n_1965), .Y(n_1954) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g824 ( .A(n_822), .Y(n_824) );
INVx1_ASAP7_75t_L g929 ( .A(n_822), .Y(n_929) );
A2O1A1Ixp33_ASAP7_75t_L g1156 ( .A1(n_829), .A2(n_1157), .B(n_1158), .C(n_1159), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_829), .A2(n_1260), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_877), .C(n_894), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_864), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_845), .B2(n_846), .Y(n_841) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_845), .A2(n_863), .B1(n_872), .B2(n_874), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_846), .A2(n_1067), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1536 ( .A1(n_846), .A2(n_1519), .B1(n_1527), .B2(n_1537), .Y(n_1536) );
OAI22xp5_ASAP7_75t_L g1640 ( .A1(n_846), .A2(n_1042), .B1(n_1641), .B2(n_1642), .Y(n_1640) );
OAI22xp33_ASAP7_75t_SL g1636 ( .A1(n_850), .A2(n_1637), .B1(n_1638), .B2(n_1639), .Y(n_1636) );
INVx3_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g927 ( .A(n_852), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_859), .B1(n_860), .B2(n_863), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
HB1xp67_ASAP7_75t_L g1571 ( .A(n_860), .Y(n_1571) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_861), .Y(n_860) );
INVxp67_ASAP7_75t_SL g1422 ( .A(n_861), .Y(n_1422) );
INVx1_ASAP7_75t_L g1662 ( .A(n_861), .Y(n_1662) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g1410 ( .A(n_862), .Y(n_1410) );
OAI22xp33_ASAP7_75t_L g1487 ( .A1(n_866), .A2(n_1430), .B1(n_1488), .B2(n_1489), .Y(n_1487) );
INVx5_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx6_ASAP7_75t_L g1608 ( .A(n_867), .Y(n_1608) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_869), .A2(n_1134), .B1(n_1135), .B2(n_1136), .C(n_1137), .Y(n_1133) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1609 ( .A1(n_872), .A2(n_1528), .B1(n_1598), .B2(n_1601), .Y(n_1609) );
OAI22xp5_ASAP7_75t_L g1610 ( .A1(n_872), .A2(n_1595), .B1(n_1605), .B2(n_1611), .Y(n_1610) );
INVx4_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI211xp5_ASAP7_75t_L g1020 ( .A1(n_874), .A2(n_1021), .B(n_1022), .C(n_1025), .Y(n_1020) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
BUFx2_ASAP7_75t_L g973 ( .A(n_883), .Y(n_973) );
OAI221xp5_ASAP7_75t_L g1932 ( .A1(n_883), .A2(n_949), .B1(n_1902), .B2(n_1914), .C(n_1933), .Y(n_1932) );
OAI22xp5_ASAP7_75t_L g1972 ( .A1(n_883), .A2(n_1425), .B1(n_1960), .B2(n_1963), .Y(n_1972) );
OAI22xp5_ASAP7_75t_L g1973 ( .A1(n_883), .A2(n_1425), .B1(n_1957), .B2(n_1967), .Y(n_1973) );
BUFx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_884), .B(n_1117), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_884), .B(n_1228), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_884), .B(n_1329), .Y(n_1328) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_884), .Y(n_1529) );
BUFx2_ASAP7_75t_SL g1611 ( .A(n_884), .Y(n_1611) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_886), .A2(n_888), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g1062 ( .A(n_893), .Y(n_1062) );
INVx2_ASAP7_75t_L g1466 ( .A(n_893), .Y(n_1466) );
OAI31xp33_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_898), .A3(n_903), .B(n_906), .Y(n_894) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI31xp33_ASAP7_75t_L g1354 ( .A1(n_906), .A2(n_1355), .A3(n_1358), .B(n_1360), .Y(n_1354) );
CKINVDCx14_ASAP7_75t_R g1515 ( .A(n_906), .Y(n_1515) );
OAI31xp33_ASAP7_75t_L g1568 ( .A1(n_906), .A2(n_1569), .A3(n_1570), .B(n_1575), .Y(n_1568) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .B1(n_1585), .B2(n_1586), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_1397), .Y(n_909) );
XNOR2x1_ASAP7_75t_L g910 ( .A(n_911), .B(n_1104), .Y(n_910) );
XNOR2xp5_ASAP7_75t_L g911 ( .A(n_912), .B(n_979), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_959), .C(n_967), .Y(n_913) );
NOR2xp33_ASAP7_75t_SL g914 ( .A(n_915), .B(n_938), .Y(n_914) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_919), .Y(n_935) );
INVx1_ASAP7_75t_L g1538 ( .A(n_919), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_920), .A2(n_937), .B1(n_941), .B2(n_949), .Y(n_948) );
OAI22xp33_ASAP7_75t_SL g921 ( .A1(n_922), .A2(n_923), .B1(n_926), .B2(n_927), .Y(n_921) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_924), .A2(n_1148), .B1(n_1149), .B2(n_1163), .Y(n_1162) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
OAI22xp33_ASAP7_75t_L g952 ( .A1(n_926), .A2(n_933), .B1(n_953), .B2(n_957), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_927), .A2(n_1072), .B1(n_1555), .B2(n_1561), .Y(n_1566) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_931), .B2(n_933), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_931), .A2(n_1066), .B1(n_1067), .B2(n_1069), .Y(n_1065) );
INVx2_ASAP7_75t_SL g931 ( .A(n_932), .Y(n_931) );
OAI33xp33_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_940), .A3(n_944), .B1(n_948), .B2(n_952), .B3(n_958), .Y(n_938) );
OAI33xp33_ASAP7_75t_L g1423 ( .A1(n_939), .A2(n_1424), .A3(n_1427), .B1(n_1429), .B2(n_1432), .B3(n_1434), .Y(n_1423) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx4_ASAP7_75t_L g1435 ( .A(n_946), .Y(n_1435) );
INVx2_ASAP7_75t_L g1654 ( .A(n_946), .Y(n_1654) );
INVx4_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_949), .A2(n_1528), .B1(n_1557), .B2(n_1558), .Y(n_1556) );
INVx3_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_957), .A2(n_1015), .B(n_1016), .C(n_1018), .Y(n_1014) );
OAI33xp33_ASAP7_75t_L g1649 ( .A1(n_958), .A2(n_1082), .A3(n_1650), .B1(n_1652), .B2(n_1653), .B3(n_1655), .Y(n_1649) );
OAI22xp33_ASAP7_75t_L g1603 ( .A1(n_962), .A2(n_1041), .B1(n_1604), .B2(n_1605), .Y(n_1603) );
OAI31xp33_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .A3(n_972), .B(n_978), .Y(n_967) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OAI31xp33_ASAP7_75t_L g1460 ( .A1(n_978), .A2(n_1461), .A3(n_1465), .B(n_1467), .Y(n_1460) );
OAI31xp33_ASAP7_75t_L g1576 ( .A1(n_978), .A2(n_1577), .A3(n_1580), .B(n_1582), .Y(n_1576) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AO22x2_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1051), .B1(n_1052), .B2(n_1103), .Y(n_980) );
INVx1_ASAP7_75t_SL g1103 ( .A(n_981), .Y(n_1103) );
XNOR2x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
NOR2x1_ASAP7_75t_L g983 ( .A(n_984), .B(n_995), .Y(n_983) );
INVxp67_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx3_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g1147 ( .A1(n_988), .A2(n_993), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
AND2x4_ASAP7_75t_L g993 ( .A(n_989), .B(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
NAND3xp33_ASAP7_75t_SL g995 ( .A(n_996), .B(n_1001), .C(n_1034), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_998), .A2(n_1009), .B1(n_1010), .B2(n_1011), .Y(n_1008) );
OAI21xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1026), .B(n_1032), .Y(n_1001) );
NAND3xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1014), .C(n_1020), .Y(n_1002) );
A2O1A1Ixp33_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B(n_1006), .C(n_1013), .Y(n_1003) );
A2O1A1Ixp33_ASAP7_75t_SL g1259 ( .A1(n_1005), .A2(n_1013), .B(n_1260), .C(n_1261), .Y(n_1259) );
NAND2xp5_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
OAI22xp5_ASAP7_75t_SL g1481 ( .A1(n_1007), .A2(n_1425), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
AOI22xp5_ASAP7_75t_L g1329 ( .A1(n_1009), .A2(n_1011), .B1(n_1302), .B2(n_1312), .Y(n_1329) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1011), .Y(n_1264) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1021), .A2(n_1040), .B1(n_1041), .B2(n_1043), .Y(n_1039) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_1029), .B(n_1116), .Y(n_1115) );
INVx3_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1030), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1036), .Y(n_1072) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1036), .Y(n_1638) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_1037), .A2(n_1165), .B1(n_1166), .B2(n_1167), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
BUFx3_ASAP7_75t_L g1201 ( .A(n_1038), .Y(n_1201) );
BUFx12f_ASAP7_75t_L g1280 ( .A(n_1038), .Y(n_1280) );
INVx5_ASAP7_75t_L g1308 ( .A(n_1038), .Y(n_1308) );
OAI22xp33_ASAP7_75t_L g1406 ( .A1(n_1041), .A2(n_1407), .B1(n_1408), .B2(n_1409), .Y(n_1406) );
OAI22xp33_ASAP7_75t_L g1955 ( .A1(n_1041), .A2(n_1956), .B1(n_1957), .B2(n_1958), .Y(n_1955) );
BUFx4f_ASAP7_75t_SL g1041 ( .A(n_1042), .Y(n_1041) );
NAND3xp33_ASAP7_75t_L g1383 ( .A(n_1049), .B(n_1384), .C(n_1388), .Y(n_1383) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
AOI33xp33_ASAP7_75t_L g1194 ( .A1(n_1050), .A2(n_1195), .A3(n_1196), .B1(n_1198), .B2(n_1202), .B3(n_1204), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1294 ( .A(n_1050), .B(n_1295), .C(n_1296), .Y(n_1294) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
NAND3xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1063), .C(n_1091), .Y(n_1054) );
NOR2xp33_ASAP7_75t_SL g1063 ( .A(n_1064), .B(n_1081), .Y(n_1063) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1068), .Y(n_1544) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1075), .Y(n_1392) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1082), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1607 ( .A1(n_1084), .A2(n_1594), .B1(n_1604), .B2(n_1608), .Y(n_1607) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_1086), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1612 ( .A1(n_1086), .A2(n_1599), .B1(n_1602), .B2(n_1608), .Y(n_1612) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_1094), .Y(n_1093) );
XNOR2x1_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1337), .Y(n_1104) );
OA22x2_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .B1(n_1240), .B2(n_1336), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
XOR2xp5_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1184), .Y(n_1107) );
XNOR2x1_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
NAND4xp75_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1119), .C(n_1147), .D(n_1150), .Y(n_1110) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
AOI211x1_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1131), .B(n_1132), .C(n_1143), .Y(n_1119) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1377 ( .A(n_1123), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_1126), .A2(n_1127), .B1(n_1128), .B2(n_1130), .Y(n_1125) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1127), .Y(n_1521) );
BUFx6f_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
OAI211xp5_ASAP7_75t_SL g1250 ( .A1(n_1135), .A2(n_1251), .B(n_1252), .C(n_1253), .Y(n_1250) );
OAI211xp5_ASAP7_75t_SL g1254 ( .A1(n_1135), .A2(n_1255), .B(n_1256), .C(n_1257), .Y(n_1254) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NAND2x2_ASAP7_75t_L g1144 ( .A(n_1141), .B(n_1145), .Y(n_1144) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx2_ASAP7_75t_SL g1145 ( .A(n_1146), .Y(n_1145) );
INVx4_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_1162), .A2(n_1164), .B(n_1168), .Y(n_1161) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
OAI21xp5_ASAP7_75t_SL g1171 ( .A1(n_1172), .A2(n_1176), .B(n_1179), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1471 ( .A(n_1173), .Y(n_1471) );
INVx3_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
XNOR2x1_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1239), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1208), .Y(n_1185) );
NAND3xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1194), .C(n_1206), .Y(n_1186) );
AOI222xp33_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1189), .B1(n_1190), .B2(n_1191), .C1(n_1192), .C2(n_1193), .Y(n_1187) );
AOI222xp33_ASAP7_75t_L g1301 ( .A1(n_1188), .A2(n_1190), .B1(n_1192), .B2(n_1302), .C1(n_1303), .C2(n_1304), .Y(n_1301) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NAND3xp33_ASAP7_75t_L g1305 ( .A(n_1204), .B(n_1306), .C(n_1309), .Y(n_1305) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NAND3xp33_ASAP7_75t_SL g1208 ( .A(n_1209), .B(n_1213), .C(n_1237), .Y(n_1208) );
OAI21xp33_ASAP7_75t_L g1219 ( .A1(n_1220), .A2(n_1222), .B(n_1226), .Y(n_1219) );
OAI21xp5_ASAP7_75t_SL g1323 ( .A1(n_1220), .A2(n_1324), .B(n_1327), .Y(n_1323) );
INVxp67_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OAI21xp5_ASAP7_75t_L g1247 ( .A1(n_1221), .A2(n_1248), .B(n_1249), .Y(n_1247) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
XNOR2xp5_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1291), .Y(n_1240) );
XOR2xp5_ASAP7_75t_L g1336 ( .A(n_1241), .B(n_1291), .Y(n_1336) );
XNOR2x1_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1243), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1277), .Y(n_1243) );
AOI21xp5_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1246), .B(n_1265), .Y(n_1244) );
NAND4xp25_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1250), .C(n_1254), .D(n_1259), .Y(n_1246) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1387 ( .A(n_1275), .Y(n_1387) );
OAI33xp33_ASAP7_75t_L g1562 ( .A1(n_1276), .A2(n_1535), .A3(n_1563), .B1(n_1564), .B2(n_1566), .B3(n_1567), .Y(n_1562) );
XNOR2x1_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1335), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1310), .Y(n_1292) );
NAND4xp25_ASAP7_75t_SL g1293 ( .A(n_1294), .B(n_1299), .C(n_1301), .D(n_1305), .Y(n_1293) );
BUFx3_ASAP7_75t_L g1389 ( .A(n_1297), .Y(n_1389) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1308), .Y(n_1393) );
NAND3xp33_ASAP7_75t_SL g1310 ( .A(n_1311), .B(n_1314), .C(n_1316), .Y(n_1310) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1339), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1354), .C(n_1362), .Y(n_1339) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1344), .Y(n_1502) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx2_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
AND4x1_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1375), .C(n_1383), .D(n_1390), .Y(n_1362) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1367), .C(n_1373), .Y(n_1363) );
INVx2_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
BUFx2_ASAP7_75t_L g1381 ( .A(n_1372), .Y(n_1381) );
INVx2_ASAP7_75t_SL g1373 ( .A(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_SL g1970 ( .A(n_1374), .Y(n_1970) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g1959 ( .A1(n_1386), .A2(n_1418), .B1(n_1960), .B2(n_1961), .Y(n_1959) );
OAI22xp5_ASAP7_75t_L g1962 ( .A1(n_1386), .A2(n_1908), .B1(n_1963), .B2(n_1964), .Y(n_1962) );
XNOR2xp5_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1496), .Y(n_1397) );
AOI22xp5_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .B1(n_1458), .B2(n_1495), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
HB1xp67_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
XNOR2xp5_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1403), .Y(n_1401) );
AND3x1_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1437), .C(n_1448), .Y(n_1403) );
NOR2xp33_ASAP7_75t_SL g1404 ( .A(n_1405), .B(n_1423), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_1408), .A2(n_1421), .B1(n_1435), .B2(n_1436), .Y(n_1434) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1958 ( .A(n_1410), .Y(n_1958) );
OAI22xp5_ASAP7_75t_L g1424 ( .A1(n_1412), .A2(n_1415), .B1(n_1425), .B2(n_1426), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_1413), .A2(n_1417), .B1(n_1430), .B2(n_1431), .Y(n_1429) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1416), .B1(n_1417), .B2(n_1418), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g1493 ( .A1(n_1416), .A2(n_1418), .B1(n_1483), .B2(n_1489), .Y(n_1493) );
OAI22xp5_ASAP7_75t_L g1906 ( .A1(n_1416), .A2(n_1907), .B1(n_1908), .B2(n_1909), .Y(n_1906) );
OAI22xp5_ASAP7_75t_L g1540 ( .A1(n_1418), .A2(n_1525), .B1(n_1533), .B2(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1426), .Y(n_1672) );
OAI22xp33_ASAP7_75t_L g1650 ( .A1(n_1430), .A2(n_1641), .B1(n_1644), .B2(n_1651), .Y(n_1650) );
OAI22xp5_ASAP7_75t_L g1974 ( .A1(n_1430), .A2(n_1431), .B1(n_1961), .B2(n_1964), .Y(n_1974) );
OAI33xp33_ASAP7_75t_L g1476 ( .A1(n_1432), .A2(n_1477), .A3(n_1480), .B1(n_1481), .B2(n_1484), .B3(n_1487), .Y(n_1476) );
OAI33xp33_ASAP7_75t_L g1968 ( .A1(n_1432), .A2(n_1969), .A3(n_1971), .B1(n_1972), .B2(n_1973), .B3(n_1974), .Y(n_1968) );
INVx2_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
OAI22xp5_ASAP7_75t_L g1484 ( .A1(n_1435), .A2(n_1436), .B1(n_1485), .B2(n_1486), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g1652 ( .A1(n_1435), .A2(n_1528), .B1(n_1637), .B2(n_1647), .Y(n_1652) );
INVx2_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
OAI31xp33_ASAP7_75t_SL g1448 ( .A1(n_1449), .A2(n_1451), .A3(n_1454), .B(n_1457), .Y(n_1448) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OAI31xp33_ASAP7_75t_L g1468 ( .A1(n_1457), .A2(n_1469), .A3(n_1470), .B(n_1474), .Y(n_1468) );
OAI31xp33_ASAP7_75t_L g1982 ( .A1(n_1457), .A2(n_1983), .A3(n_1984), .B(n_1987), .Y(n_1982) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1458), .Y(n_1495) );
NAND3xp33_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1468), .C(n_1475), .Y(n_1459) );
NOR2xp33_ASAP7_75t_SL g1475 ( .A(n_1476), .B(n_1490), .Y(n_1475) );
OAI22xp5_ASAP7_75t_L g1496 ( .A1(n_1497), .A2(n_1545), .B1(n_1583), .B2(n_1584), .Y(n_1496) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1497), .Y(n_1583) );
OAI221xp5_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1500), .B1(n_1508), .B2(n_1515), .C(n_1516), .Y(n_1498) );
AOI31xp33_ASAP7_75t_SL g1915 ( .A1(n_1499), .A2(n_1916), .A3(n_1919), .B(n_1925), .Y(n_1915) );
NOR3xp33_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1503), .C(n_1504), .Y(n_1500) );
NOR3xp33_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1511), .C(n_1514), .Y(n_1508) );
AOI31xp33_ASAP7_75t_L g1934 ( .A1(n_1515), .A2(n_1935), .A3(n_1940), .B(n_1941), .Y(n_1934) );
NOR2xp33_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1534), .Y(n_1516) );
INVx2_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx5_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx2_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1545), .Y(n_1584) );
BUFx2_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NAND3xp33_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1568), .C(n_1576), .Y(n_1547) );
NOR2xp33_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1562), .Y(n_1548) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
XOR2xp5_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1629), .Y(n_1586) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
BUFx2_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
AND3x1_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1613), .C(n_1621), .Y(n_1590) );
NOR2xp33_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1606), .Y(n_1591) );
OAI22xp5_ASAP7_75t_L g1655 ( .A1(n_1608), .A2(n_1639), .B1(n_1648), .B2(n_1656), .Y(n_1655) );
OAI22xp5_ASAP7_75t_L g1653 ( .A1(n_1611), .A2(n_1642), .B1(n_1645), .B2(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
NAND3xp33_ASAP7_75t_L g1633 ( .A(n_1634), .B(n_1657), .C(n_1668), .Y(n_1633) );
NOR2xp33_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1649), .Y(n_1634) );
OAI31xp33_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1661), .A3(n_1666), .B(n_1667), .Y(n_1657) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
OAI221xp5_ASAP7_75t_L g1677 ( .A1(n_1678), .A2(n_1893), .B1(n_1895), .B2(n_1942), .C(n_1945), .Y(n_1677) );
NOR3xp33_ASAP7_75t_L g1678 ( .A(n_1679), .B(n_1873), .C(n_1887), .Y(n_1678) );
OAI221xp5_ASAP7_75t_L g1679 ( .A1(n_1680), .A2(n_1772), .B1(n_1794), .B2(n_1830), .C(n_1831), .Y(n_1679) );
OAI21xp5_ASAP7_75t_SL g1680 ( .A1(n_1681), .A2(n_1718), .B(n_1766), .Y(n_1680) );
OAI22xp5_ASAP7_75t_L g1889 ( .A1(n_1681), .A2(n_1745), .B1(n_1818), .B2(n_1890), .Y(n_1889) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
NAND2xp5_ASAP7_75t_SL g1682 ( .A(n_1683), .B(n_1713), .Y(n_1682) );
AOI211xp5_ASAP7_75t_L g1881 ( .A1(n_1683), .A2(n_1759), .B(n_1882), .C(n_1883), .Y(n_1881) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
OR2x2_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1700), .Y(n_1684) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1685), .B(n_1738), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1685), .B(n_1761), .Y(n_1777) );
CKINVDCx5p33_ASAP7_75t_R g1785 ( .A(n_1685), .Y(n_1785) );
NAND2xp5_ASAP7_75t_L g1796 ( .A(n_1685), .B(n_1797), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1685), .B(n_1817), .Y(n_1816) );
OAI21xp5_ASAP7_75t_SL g1886 ( .A1(n_1685), .A2(n_1817), .B(n_1883), .Y(n_1886) );
INVx4_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
OR2x2_ASAP7_75t_L g1765 ( .A(n_1686), .B(n_1729), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1686), .B(n_1774), .Y(n_1773) );
INVx4_ASAP7_75t_L g1782 ( .A(n_1686), .Y(n_1782) );
NOR2xp33_ASAP7_75t_L g1788 ( .A(n_1686), .B(n_1731), .Y(n_1788) );
NOR2xp33_ASAP7_75t_L g1792 ( .A(n_1686), .B(n_1793), .Y(n_1792) );
AOI322xp5_ASAP7_75t_L g1798 ( .A1(n_1686), .A2(n_1799), .A3(n_1801), .B1(n_1803), .B2(n_1805), .C1(n_1806), .C2(n_1808), .Y(n_1798) );
AND2x2_ASAP7_75t_L g1805 ( .A(n_1686), .B(n_1734), .Y(n_1805) );
NAND2xp5_ASAP7_75t_SL g1825 ( .A(n_1686), .B(n_1729), .Y(n_1825) );
NAND2xp5_ASAP7_75t_L g1872 ( .A(n_1686), .B(n_1713), .Y(n_1872) );
AND2x4_ASAP7_75t_SL g1686 ( .A(n_1687), .B(n_1695), .Y(n_1686) );
AND2x4_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
AND2x6_ASAP7_75t_L g1693 ( .A(n_1689), .B(n_1694), .Y(n_1693) );
AND2x6_ASAP7_75t_L g1696 ( .A(n_1689), .B(n_1697), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1689), .B(n_1699), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1689), .B(n_1699), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1752 ( .A(n_1689), .B(n_1690), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1689), .B(n_1699), .Y(n_1757) );
HB1xp67_ASAP7_75t_L g1992 ( .A(n_1690), .Y(n_1992) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1692), .Y(n_1690) );
INVx2_ASAP7_75t_L g1754 ( .A(n_1693), .Y(n_1754) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1700), .Y(n_1882) );
OR2x2_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1705), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1701), .B(n_1734), .Y(n_1733) );
OR2x2_ASAP7_75t_L g1742 ( .A(n_1701), .B(n_1743), .Y(n_1742) );
OR2x2_ASAP7_75t_L g1842 ( .A(n_1701), .B(n_1707), .Y(n_1842) );
NAND2xp5_ASAP7_75t_L g1876 ( .A(n_1701), .B(n_1788), .Y(n_1876) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1703), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1702), .B(n_1703), .Y(n_1729) );
OR2x2_ASAP7_75t_L g1778 ( .A(n_1705), .B(n_1728), .Y(n_1778) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1705), .Y(n_1810) );
OR2x2_ASAP7_75t_L g1824 ( .A(n_1705), .B(n_1825), .Y(n_1824) );
NAND2xp5_ASAP7_75t_L g1858 ( .A(n_1705), .B(n_1859), .Y(n_1858) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1710), .Y(n_1705) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
OR2x2_ASAP7_75t_L g1731 ( .A(n_1707), .B(n_1710), .Y(n_1731) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1707), .B(n_1735), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1707), .B(n_1710), .Y(n_1738) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1707), .Y(n_1802) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1707), .B(n_1729), .Y(n_1829) );
NAND3xp33_ASAP7_75t_L g1833 ( .A(n_1707), .B(n_1749), .C(n_1769), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1709), .Y(n_1707) );
INVx2_ASAP7_75t_L g1735 ( .A(n_1710), .Y(n_1735) );
OR2x2_ASAP7_75t_L g1869 ( .A(n_1710), .B(n_1729), .Y(n_1869) );
NAND2x1p5_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1712), .Y(n_1710) );
AOI221xp5_ASAP7_75t_L g1772 ( .A1(n_1713), .A2(n_1745), .B1(n_1773), .B2(n_1775), .C(n_1786), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1891 ( .A(n_1713), .B(n_1784), .Y(n_1891) );
INVx2_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1714), .B(n_1721), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1828 ( .A(n_1714), .B(n_1782), .Y(n_1828) );
OAI322xp33_ASAP7_75t_L g1843 ( .A1(n_1714), .A2(n_1726), .A3(n_1766), .B1(n_1844), .B2(n_1847), .C1(n_1848), .C2(n_1851), .Y(n_1843) );
OR2x2_ASAP7_75t_L g1855 ( .A(n_1714), .B(n_1768), .Y(n_1855) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
OR2x2_ASAP7_75t_L g1740 ( .A(n_1715), .B(n_1721), .Y(n_1740) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1715), .Y(n_1762) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1717), .Y(n_1715) );
OAI211xp5_ASAP7_75t_L g1718 ( .A1(n_1719), .A2(n_1725), .B(n_1736), .C(n_1758), .Y(n_1718) );
NOR2xp33_ASAP7_75t_L g1823 ( .A(n_1719), .B(n_1824), .Y(n_1823) );
OAI21xp5_ASAP7_75t_L g1892 ( .A1(n_1719), .A2(n_1740), .B(n_1806), .Y(n_1892) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
AOI21xp5_ASAP7_75t_L g1791 ( .A1(n_1720), .A2(n_1748), .B(n_1792), .Y(n_1791) );
NAND2xp5_ASAP7_75t_L g1822 ( .A(n_1720), .B(n_1763), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1835 ( .A(n_1720), .B(n_1836), .Y(n_1835) );
INVx2_ASAP7_75t_L g1745 ( .A(n_1721), .Y(n_1745) );
OAI21xp33_ASAP7_75t_L g1746 ( .A1(n_1721), .A2(n_1747), .B(n_1748), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1808 ( .A(n_1721), .B(n_1769), .Y(n_1808) );
OR2x2_ASAP7_75t_L g1818 ( .A(n_1721), .B(n_1762), .Y(n_1818) );
OR2x2_ASAP7_75t_L g1847 ( .A(n_1721), .B(n_1769), .Y(n_1847) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1721), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1885 ( .A(n_1721), .B(n_1768), .Y(n_1885) );
INVx2_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1790 ( .A(n_1722), .B(n_1762), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1724), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1732), .Y(n_1725) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1784 ( .A(n_1727), .B(n_1785), .Y(n_1784) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1728), .B(n_1730), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1728), .B(n_1734), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1728), .B(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1729), .B(n_1738), .Y(n_1737) );
OR2x2_ASAP7_75t_L g1793 ( .A(n_1729), .B(n_1735), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1729), .B(n_1802), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1864 ( .A(n_1729), .B(n_1735), .Y(n_1864) );
NAND2xp5_ASAP7_75t_L g1815 ( .A(n_1730), .B(n_1816), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1845 ( .A(n_1730), .B(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
OR2x2_ASAP7_75t_L g1764 ( .A(n_1731), .B(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
NAND2xp5_ASAP7_75t_L g1851 ( .A(n_1734), .B(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1734), .Y(n_1859) );
OAI211xp5_ASAP7_75t_L g1867 ( .A1(n_1734), .A2(n_1868), .B(n_1870), .C(n_1871), .Y(n_1867) );
NAND3xp33_ASAP7_75t_L g1880 ( .A(n_1734), .B(n_1767), .C(n_1777), .Y(n_1880) );
AOI221xp5_ASAP7_75t_L g1736 ( .A1(n_1737), .A2(n_1739), .B1(n_1741), .B2(n_1744), .C(n_1746), .Y(n_1736) );
NAND2x1_ASAP7_75t_L g1807 ( .A(n_1737), .B(n_1782), .Y(n_1807) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1738), .Y(n_1743) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
OR2x2_ASAP7_75t_L g1812 ( .A(n_1740), .B(n_1813), .Y(n_1812) );
OAI21xp33_ASAP7_75t_L g1840 ( .A1(n_1741), .A2(n_1811), .B(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
NOR2x1_ASAP7_75t_L g1781 ( .A(n_1743), .B(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1748), .Y(n_1830) );
OAI321xp33_ASAP7_75t_L g1861 ( .A1(n_1748), .A2(n_1847), .A3(n_1862), .B1(n_1863), .B2(n_1866), .C(n_1867), .Y(n_1861) );
OAI221xp5_ASAP7_75t_L g1873 ( .A1(n_1748), .A2(n_1874), .B1(n_1881), .B2(n_1884), .C(n_1886), .Y(n_1873) );
INVx2_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1750), .B(n_1767), .Y(n_1766) );
NOR2xp33_ASAP7_75t_SL g1870 ( .A(n_1750), .B(n_1769), .Y(n_1870) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
OAI221xp5_ASAP7_75t_L g1751 ( .A1(n_1752), .A2(n_1753), .B1(n_1754), .B2(n_1755), .C(n_1756), .Y(n_1751) );
CKINVDCx5p33_ASAP7_75t_R g1894 ( .A(n_1752), .Y(n_1894) );
INVxp67_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1763), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1779 ( .A(n_1760), .B(n_1780), .Y(n_1779) );
NAND2xp5_ASAP7_75t_L g1844 ( .A(n_1760), .B(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
OR2x2_ASAP7_75t_L g1800 ( .A(n_1761), .B(n_1768), .Y(n_1800) );
NOR3xp33_ASAP7_75t_L g1838 ( .A(n_1761), .B(n_1824), .C(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
AOI221xp5_ASAP7_75t_L g1853 ( .A1(n_1764), .A2(n_1799), .B1(n_1851), .B2(n_1854), .C(n_1856), .Y(n_1853) );
INVx1_ASAP7_75t_L g1852 ( .A(n_1765), .Y(n_1852) );
AOI31xp33_ASAP7_75t_L g1856 ( .A1(n_1767), .A2(n_1846), .A3(n_1857), .B(n_1860), .Y(n_1856) );
NOR2xp33_ASAP7_75t_L g1883 ( .A(n_1767), .B(n_1778), .Y(n_1883) );
CKINVDCx14_ASAP7_75t_R g1767 ( .A(n_1768), .Y(n_1767) );
OR2x2_ASAP7_75t_L g1804 ( .A(n_1768), .B(n_1790), .Y(n_1804) );
OR2x2_ASAP7_75t_L g1821 ( .A(n_1768), .B(n_1818), .Y(n_1821) );
OAI21xp5_ASAP7_75t_L g1863 ( .A1(n_1768), .A2(n_1864), .B(n_1865), .Y(n_1863) );
INVx3_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1769), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1769), .B(n_1850), .Y(n_1849) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1770), .B(n_1771), .Y(n_1769) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1774), .Y(n_1789) );
OAI211xp5_ASAP7_75t_L g1775 ( .A1(n_1776), .A2(n_1778), .B(n_1779), .C(n_1783), .Y(n_1775) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1778), .Y(n_1797) );
O2A1O1Ixp33_ASAP7_75t_SL g1887 ( .A1(n_1778), .A2(n_1888), .B(n_1889), .C(n_1892), .Y(n_1887) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1781), .Y(n_1820) );
O2A1O1Ixp33_ASAP7_75t_L g1874 ( .A1(n_1781), .A2(n_1799), .B(n_1875), .C(n_1877), .Y(n_1874) );
CKINVDCx5p33_ASAP7_75t_R g1836 ( .A(n_1782), .Y(n_1836) );
NOR2xp33_ASAP7_75t_L g1841 ( .A(n_1782), .B(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
OR2x2_ASAP7_75t_L g1878 ( .A(n_1785), .B(n_1829), .Y(n_1878) );
A2O1A1Ixp33_ASAP7_75t_L g1786 ( .A1(n_1787), .A2(n_1789), .B(n_1790), .C(n_1791), .Y(n_1786) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
OAI211xp5_ASAP7_75t_SL g1795 ( .A1(n_1790), .A2(n_1796), .B(n_1798), .C(n_1809), .Y(n_1795) );
CKINVDCx5p33_ASAP7_75t_R g1860 ( .A(n_1790), .Y(n_1860) );
NAND2xp5_ASAP7_75t_L g1879 ( .A(n_1792), .B(n_1808), .Y(n_1879) );
INVx1_ASAP7_75t_L g1865 ( .A(n_1793), .Y(n_1865) );
NOR5xp2_ASAP7_75t_L g1794 ( .A(n_1795), .B(n_1814), .C(n_1819), .D(n_1823), .E(n_1826), .Y(n_1794) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1805), .Y(n_1862) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1808), .Y(n_1839) );
NAND2xp5_ASAP7_75t_L g1809 ( .A(n_1810), .B(n_1811), .Y(n_1809) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1816), .Y(n_1866) );
CKINVDCx5p33_ASAP7_75t_R g1817 ( .A(n_1818), .Y(n_1817) );
OAI21xp33_ASAP7_75t_L g1819 ( .A1(n_1820), .A2(n_1821), .B(n_1822), .Y(n_1819) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1825), .Y(n_1846) );
NOR2xp33_ASAP7_75t_L g1826 ( .A(n_1827), .B(n_1829), .Y(n_1826) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
NOR4xp25_ASAP7_75t_L g1831 ( .A(n_1832), .B(n_1843), .C(n_1853), .D(n_1861), .Y(n_1831) );
OAI211xp5_ASAP7_75t_SL g1832 ( .A1(n_1833), .A2(n_1834), .B(n_1837), .C(n_1840), .Y(n_1832) );
INVxp67_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVxp67_ASAP7_75t_SL g1837 ( .A(n_1838), .Y(n_1837) );
OAI211xp5_ASAP7_75t_L g1877 ( .A1(n_1848), .A2(n_1878), .B(n_1879), .C(n_1880), .Y(n_1877) );
INVx1_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1870), .Y(n_1888) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1876), .Y(n_1875) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
INVxp67_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
CKINVDCx20_ASAP7_75t_R g1893 ( .A(n_1894), .Y(n_1893) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1896), .Y(n_1895) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
NOR4xp25_ASAP7_75t_L g1898 ( .A(n_1899), .B(n_1915), .C(n_1928), .D(n_1934), .Y(n_1898) );
INVx1_ASAP7_75t_L g1910 ( .A(n_1911), .Y(n_1910) );
INVx1_ASAP7_75t_L g1920 ( .A(n_1921), .Y(n_1920) );
INVx3_ASAP7_75t_L g1942 ( .A(n_1943), .Y(n_1942) );
HB1xp67_ASAP7_75t_L g1946 ( .A(n_1947), .Y(n_1946) );
BUFx3_ASAP7_75t_L g1947 ( .A(n_1948), .Y(n_1947) );
INVxp33_ASAP7_75t_SL g1949 ( .A(n_1950), .Y(n_1949) );
HB1xp67_ASAP7_75t_L g1951 ( .A(n_1952), .Y(n_1951) );
NAND3xp33_ASAP7_75t_L g1952 ( .A(n_1953), .B(n_1975), .C(n_1982), .Y(n_1952) );
NOR2xp33_ASAP7_75t_L g1953 ( .A(n_1954), .B(n_1968), .Y(n_1953) );
INVx1_ASAP7_75t_L g1969 ( .A(n_1970), .Y(n_1969) );
HB1xp67_ASAP7_75t_L g1988 ( .A(n_1989), .Y(n_1988) );
HB1xp67_ASAP7_75t_L g1989 ( .A(n_1990), .Y(n_1989) );
OAI21xp5_ASAP7_75t_L g1990 ( .A1(n_1991), .A2(n_1992), .B(n_1993), .Y(n_1990) );
INVx1_ASAP7_75t_L g1993 ( .A(n_1994), .Y(n_1993) );
endmodule