module fake_jpeg_6098_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVxp67_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_0),
.A2(n_6),
.B1(n_4),
.B2(n_3),
.Y(n_12)
);

NAND2xp33_ASAP7_75t_SL g13 ( 
.A(n_1),
.B(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

AO22x1_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_24),
.B1(n_14),
.B2(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_15),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_12),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_7),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.C(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_32),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_36),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_28),
.B(n_38),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_42),
.B(n_34),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_40),
.Y(n_47)
);

FAx1_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_44),
.CI(n_42),
.CON(n_50),
.SN(n_50)
);


endmodule