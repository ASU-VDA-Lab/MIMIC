module real_aes_15888_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_1588, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_1588;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_0), .A2(n_88), .B1(n_395), .B2(n_398), .Y(n_783) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_0), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_1), .A2(n_66), .B1(n_608), .B2(n_920), .Y(n_919) );
INVxp33_ASAP7_75t_SL g958 ( .A(n_1), .Y(n_958) );
CKINVDCx5p33_ASAP7_75t_R g1541 ( .A(n_2), .Y(n_1541) );
INVx1_ASAP7_75t_L g523 ( .A(n_3), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_3), .A2(n_149), .B1(n_542), .B2(n_546), .C(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g767 ( .A(n_4), .Y(n_767) );
INVx1_ASAP7_75t_L g1042 ( .A(n_5), .Y(n_1042) );
OAI221xp5_ASAP7_75t_SL g1073 ( .A1(n_5), .A2(n_89), .B1(n_335), .B2(n_717), .C(n_837), .Y(n_1073) );
INVx1_ASAP7_75t_L g1118 ( .A(n_6), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_6), .A2(n_117), .B1(n_648), .B2(n_656), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_7), .A2(n_68), .B1(n_459), .B2(n_572), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_7), .A2(n_36), .B1(n_395), .B2(n_398), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_8), .A2(n_244), .B1(n_654), .B2(n_657), .C(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g681 ( .A(n_8), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_9), .A2(n_197), .B1(n_713), .B2(n_715), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g754 ( .A(n_9), .Y(n_754) );
INVx1_ASAP7_75t_L g297 ( .A(n_10), .Y(n_297) );
AND2x2_ASAP7_75t_L g415 ( .A(n_10), .B(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_10), .B(n_307), .Y(n_426) );
AND2x2_ASAP7_75t_L g462 ( .A(n_10), .B(n_230), .Y(n_462) );
INVx1_ASAP7_75t_L g834 ( .A(n_11), .Y(n_834) );
OAI221xp5_ASAP7_75t_SL g891 ( .A1(n_11), .A2(n_269), .B1(n_892), .B2(n_896), .C(n_900), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_12), .A2(n_221), .B1(n_335), .B2(n_837), .C(n_1080), .Y(n_1108) );
OA222x2_ASAP7_75t_L g1139 ( .A1(n_12), .A2(n_49), .B1(n_226), .B2(n_537), .C1(n_796), .C2(n_946), .Y(n_1139) );
INVx1_ASAP7_75t_L g1160 ( .A(n_13), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_13), .A2(n_259), .B1(n_332), .B2(n_1171), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1196 ( .A1(n_14), .A2(n_127), .B1(n_386), .B2(n_501), .Y(n_1196) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_14), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_15), .B(n_1248), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_15), .B(n_113), .Y(n_1250) );
INVx2_ASAP7_75t_L g1254 ( .A(n_15), .Y(n_1254) );
OAI21xp5_ASAP7_75t_SL g1580 ( .A1(n_16), .A2(n_866), .B(n_1581), .Y(n_1580) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_17), .A2(n_232), .B1(n_386), .B2(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_17), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_18), .A2(n_355), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g812 ( .A(n_18), .Y(n_812) );
INVx1_ASAP7_75t_L g1539 ( .A(n_19), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_20), .A2(n_156), .B1(n_509), .B2(n_519), .Y(n_789) );
AOI32xp33_ASAP7_75t_L g800 ( .A1(n_20), .A2(n_801), .A3(n_802), .B1(n_804), .B2(n_1588), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_21), .A2(n_210), .B1(n_646), .B2(n_1510), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_21), .A2(n_237), .B1(n_355), .B2(n_1517), .Y(n_1516) );
AOI22xp5_ASAP7_75t_L g1259 ( .A1(n_22), .A2(n_188), .B1(n_1255), .B2(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1205 ( .A(n_23), .Y(n_1205) );
AND2x2_ASAP7_75t_L g781 ( .A(n_24), .B(n_782), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_24), .A2(n_156), .B1(n_587), .B2(n_821), .C(n_822), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g1291 ( .A1(n_25), .A2(n_176), .B1(n_1249), .B2(n_1255), .Y(n_1291) );
INVx1_ASAP7_75t_L g393 ( .A(n_26), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_27), .A2(n_73), .B1(n_357), .B2(n_703), .C(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g963 ( .A1(n_27), .A2(n_29), .B1(n_964), .B2(n_965), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_28), .Y(n_997) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_29), .A2(n_141), .B1(n_505), .B2(n_608), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_30), .A2(n_200), .B1(n_1245), .B2(n_1252), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1554 ( .A1(n_31), .A2(n_173), .B1(n_507), .B2(n_782), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1573 ( .A1(n_31), .A2(n_144), .B1(n_1570), .B2(n_1574), .Y(n_1573) );
AOI222xp33_ASAP7_75t_L g1212 ( .A1(n_32), .A2(n_181), .B1(n_217), .B2(n_363), .C1(n_383), .C2(n_1125), .Y(n_1212) );
INVx1_ASAP7_75t_L g1235 ( .A(n_32), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_33), .B(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_33), .A2(n_274), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g1149 ( .A(n_34), .Y(n_1149) );
INVx1_ASAP7_75t_L g926 ( .A(n_35), .Y(n_926) );
OA222x2_ASAP7_75t_L g945 ( .A1(n_35), .A2(n_171), .B1(n_275), .B2(n_537), .C1(n_946), .C2(n_948), .Y(n_945) );
OAI211xp5_ASAP7_75t_L g568 ( .A1(n_36), .A2(n_408), .B(n_569), .C(n_597), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_37), .A2(n_205), .B1(n_379), .B2(n_916), .C(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g961 ( .A(n_37), .Y(n_961) );
INVx1_ASAP7_75t_L g1545 ( .A(n_38), .Y(n_1545) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_39), .A2(n_703), .B(n_704), .C(n_707), .Y(n_702) );
INVx1_ASAP7_75t_L g748 ( .A(n_39), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g1265 ( .A1(n_40), .A2(n_119), .B1(n_1245), .B2(n_1252), .Y(n_1265) );
INVx1_ASAP7_75t_L g662 ( .A(n_41), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_42), .A2(n_74), .B1(n_677), .B2(n_849), .Y(n_848) );
INVxp67_ASAP7_75t_SL g902 ( .A(n_42), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g1272 ( .A1(n_43), .A2(n_206), .B1(n_1245), .B2(n_1255), .Y(n_1272) );
OAI21xp33_ASAP7_75t_L g1151 ( .A1(n_44), .A2(n_946), .B(n_1152), .Y(n_1151) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_44), .A2(n_55), .B1(n_674), .B2(n_1182), .C(n_1183), .Y(n_1181) );
AOI22xp5_ASAP7_75t_L g1290 ( .A1(n_45), .A2(n_108), .B1(n_1245), .B2(n_1252), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_46), .A2(n_124), .B1(n_504), .B2(n_508), .C(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g549 ( .A(n_46), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_47), .A2(n_79), .B1(n_542), .B2(n_1510), .Y(n_1509) );
AOI22xp33_ASAP7_75t_SL g1520 ( .A1(n_47), .A2(n_87), .B1(n_509), .B2(n_672), .Y(n_1520) );
INVx1_ASAP7_75t_L g325 ( .A(n_48), .Y(n_325) );
INVx1_ASAP7_75t_L g342 ( .A(n_48), .Y(n_342) );
INVx1_ASAP7_75t_L g1106 ( .A(n_49), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_50), .A2(n_158), .B1(n_482), .B2(n_964), .Y(n_1057) );
INVx1_ASAP7_75t_L g1078 ( .A(n_50), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_51), .A2(n_250), .B1(n_332), .B2(n_337), .C(n_343), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_51), .A2(n_134), .B1(n_459), .B2(n_572), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_52), .A2(n_98), .B1(n_518), .B2(n_520), .C(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g557 ( .A(n_52), .Y(n_557) );
INVx1_ASAP7_75t_L g1161 ( .A(n_53), .Y(n_1161) );
INVx1_ASAP7_75t_L g372 ( .A(n_54), .Y(n_372) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_55), .Y(n_1187) );
INVx1_ASAP7_75t_L g1467 ( .A(n_56), .Y(n_1467) );
OAI221xp5_ASAP7_75t_L g1488 ( .A1(n_56), .A2(n_109), .B1(n_717), .B2(n_1489), .C(n_1493), .Y(n_1488) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_57), .A2(n_164), .B1(n_1199), .B2(n_1201), .C(n_1203), .Y(n_1198) );
AOI221xp5_ASAP7_75t_L g1231 ( .A1(n_57), .A2(n_223), .B1(n_818), .B2(n_1232), .C(n_1234), .Y(n_1231) );
OAI221xp5_ASAP7_75t_L g1195 ( .A1(n_58), .A2(n_249), .B1(n_332), .B2(n_337), .C(n_343), .Y(n_1195) );
OAI21xp33_ASAP7_75t_SL g1223 ( .A1(n_58), .A2(n_470), .B(n_537), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_59), .A2(n_243), .B1(n_386), .B2(n_501), .Y(n_604) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_59), .Y(n_623) );
INVx1_ASAP7_75t_L g290 ( .A(n_60), .Y(n_290) );
INVx2_ASAP7_75t_L g328 ( .A(n_61), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_62), .A2(n_83), .B1(n_1252), .B2(n_1260), .Y(n_1273) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_63), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_63), .A2(n_343), .B(n_689), .C(n_690), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g1206 ( .A1(n_64), .A2(n_67), .B1(n_395), .B2(n_398), .Y(n_1206) );
INVxp67_ASAP7_75t_SL g1218 ( .A(n_64), .Y(n_1218) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_65), .A2(n_378), .B(n_379), .Y(n_377) );
INVxp67_ASAP7_75t_L g437 ( .A(n_65), .Y(n_437) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_66), .Y(n_962) );
INVx1_ASAP7_75t_L g1222 ( .A(n_67), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_68), .A2(n_129), .B1(n_332), .B2(n_337), .C(n_343), .Y(n_603) );
INVx1_ASAP7_75t_L g526 ( .A(n_69), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_70), .A2(n_247), .B1(n_363), .B2(n_851), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_70), .A2(n_215), .B1(n_821), .B2(n_822), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_71), .A2(n_183), .B1(n_657), .B2(n_954), .C(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1079 ( .A(n_71), .Y(n_1079) );
INVx1_ASAP7_75t_L g1194 ( .A(n_72), .Y(n_1194) );
OAI21xp33_ASAP7_75t_L g1219 ( .A1(n_72), .A2(n_796), .B(n_1220), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_73), .A2(n_205), .B1(n_953), .B2(n_954), .C(n_955), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_74), .A2(n_101), .B1(n_878), .B2(n_880), .C(n_882), .Y(n_877) );
INVx1_ASAP7_75t_L g639 ( .A(n_75), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g1112 ( .A(n_76), .Y(n_1112) );
INVx1_ASAP7_75t_L g1120 ( .A(n_77), .Y(n_1120) );
AOI221x1_ASAP7_75t_SL g1132 ( .A1(n_77), .A2(n_104), .B1(n_482), .B2(n_657), .C(n_1133), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g1279 ( .A1(n_78), .A2(n_136), .B1(n_1245), .B2(n_1252), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_79), .A2(n_191), .B1(n_509), .B2(n_917), .Y(n_1515) );
INVx1_ASAP7_75t_L g939 ( .A(n_80), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_80), .B(n_408), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_81), .A2(n_1533), .B1(n_1534), .B2(n_1535), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g1533 ( .A(n_81), .Y(n_1533) );
XOR2x2_ASAP7_75t_L g694 ( .A(n_82), .B(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g1548 ( .A1(n_84), .A2(n_95), .B1(n_1517), .B2(n_1549), .Y(n_1548) );
AOI221xp5_ASAP7_75t_L g1567 ( .A1(n_84), .A2(n_133), .B1(n_801), .B2(n_818), .C(n_882), .Y(n_1567) );
XOR2x1_ASAP7_75t_L g762 ( .A(n_85), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g592 ( .A(n_86), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g1512 ( .A1(n_87), .A2(n_191), .B1(n_875), .B2(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g764 ( .A(n_88), .Y(n_764) );
INVx1_ASAP7_75t_L g1051 ( .A(n_89), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_90), .A2(n_235), .B1(n_642), .B2(n_646), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g684 ( .A1(n_90), .A2(n_379), .B(n_518), .Y(n_684) );
INVx1_ASAP7_75t_L g1103 ( .A(n_91), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_91), .A2(n_221), .B1(n_457), .B2(n_466), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_92), .A2(n_184), .B1(n_395), .B2(n_398), .Y(n_394) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_92), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_93), .A2(n_135), .B1(n_1245), .B2(n_1252), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_94), .A2(n_134), .B1(n_395), .B2(n_398), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g723 ( .A1(n_94), .A2(n_408), .B(n_724), .C(n_727), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g1575 ( .A1(n_95), .A2(n_208), .B1(n_880), .B2(n_1576), .C(n_1577), .Y(n_1575) );
INVx1_ASAP7_75t_L g940 ( .A(n_96), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_96), .A2(n_186), .B1(n_459), .B2(n_572), .Y(n_966) );
OAI221xp5_ASAP7_75t_L g1039 ( .A1(n_97), .A2(n_278), .B1(n_734), .B2(n_957), .C(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1064 ( .A(n_97), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_98), .A2(n_194), .B1(n_542), .B2(n_546), .C(n_548), .Y(n_541) );
INVx1_ASAP7_75t_L g710 ( .A(n_99), .Y(n_710) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_100), .Y(n_292) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_100), .B(n_290), .Y(n_1246) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_101), .A2(n_167), .B1(n_679), .B2(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g720 ( .A(n_102), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_103), .Y(n_1000) );
INVx1_ASAP7_75t_L g1130 ( .A(n_104), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_105), .A2(n_165), .B1(n_851), .B2(n_923), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_105), .A2(n_107), .B1(n_965), .B2(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g625 ( .A(n_106), .Y(n_625) );
INVx1_ASAP7_75t_L g1001 ( .A(n_107), .Y(n_1001) );
INVx1_ASAP7_75t_L g1474 ( .A(n_109), .Y(n_1474) );
AOI22xp33_ASAP7_75t_SL g1264 ( .A1(n_110), .A2(n_123), .B1(n_1249), .B2(n_1255), .Y(n_1264) );
AOI22xp33_ASAP7_75t_SL g1157 ( .A1(n_111), .A2(n_185), .B1(n_644), .B2(n_817), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_111), .A2(n_174), .B1(n_379), .B2(n_703), .C(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g843 ( .A(n_112), .Y(n_843) );
INVx1_ASAP7_75t_L g1248 ( .A(n_113), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_113), .B(n_1254), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g784 ( .A1(n_114), .A2(n_274), .B1(n_683), .B2(n_785), .C(n_788), .Y(n_784) );
INVx1_ASAP7_75t_L g813 ( .A(n_114), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_115), .A2(n_970), .B1(n_971), .B2(n_1027), .Y(n_969) );
INVx1_ASAP7_75t_L g1027 ( .A(n_115), .Y(n_1027) );
INVx1_ASAP7_75t_L g718 ( .A(n_116), .Y(n_718) );
INVx1_ASAP7_75t_L g1126 ( .A(n_117), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_118), .A2(n_277), .B1(n_1245), .B2(n_1249), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_120), .A2(n_265), .B1(n_386), .B2(n_501), .Y(n_769) );
INVxp33_ASAP7_75t_L g824 ( .A(n_120), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_121), .A2(n_161), .B1(n_395), .B2(n_398), .Y(n_516) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_121), .Y(n_563) );
INVx1_ASAP7_75t_L g1046 ( .A(n_122), .Y(n_1046) );
OAI21xp33_ASAP7_75t_L g1071 ( .A1(n_122), .A2(n_864), .B(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g555 ( .A(n_124), .Y(n_555) );
INVx2_ASAP7_75t_L g330 ( .A(n_125), .Y(n_330) );
INVx1_ASAP7_75t_L g360 ( .A(n_125), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_125), .B(n_328), .Y(n_389) );
INVx1_ASAP7_75t_L g374 ( .A(n_126), .Y(n_374) );
INVxp67_ASAP7_75t_SL g1215 ( .A(n_127), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_128), .A2(n_238), .B1(n_1245), .B2(n_1252), .Y(n_1261) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_129), .Y(n_599) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_130), .A2(n_159), .B1(n_332), .B2(n_337), .C(n_343), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_130), .B(n_486), .Y(n_803) );
XOR2xp5_ASAP7_75t_L g1094 ( .A(n_131), .B(n_1095), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_132), .A2(n_150), .B1(n_586), .B2(n_594), .C(n_596), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_132), .A2(n_162), .B1(n_355), .B2(n_608), .C(n_617), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_133), .A2(n_144), .B1(n_849), .B2(n_1517), .C(n_1556), .Y(n_1555) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_136), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_136), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g1158 ( .A1(n_137), .A2(n_261), .B1(n_965), .B2(n_1061), .Y(n_1158) );
AOI221xp5_ASAP7_75t_L g1177 ( .A1(n_137), .A2(n_212), .B1(n_355), .B2(n_357), .C(n_703), .Y(n_1177) );
INVx1_ASAP7_75t_L g590 ( .A(n_138), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_138), .A2(n_280), .B1(n_607), .B2(n_608), .C(n_609), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g1122 ( .A(n_139), .Y(n_1122) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_140), .A2(n_195), .B1(n_332), .B2(n_337), .C(n_343), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_140), .A2(n_470), .B(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_SL g956 ( .A(n_141), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g1104 ( .A1(n_142), .A2(n_148), .B1(n_719), .B2(n_918), .Y(n_1104) );
INVx1_ASAP7_75t_L g1142 ( .A(n_142), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_143), .A2(n_190), .B1(n_1013), .B2(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1089 ( .A(n_143), .Y(n_1089) );
XOR2x2_ASAP7_75t_L g313 ( .A(n_145), .B(n_314), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g1277 ( .A1(n_146), .A2(n_254), .B1(n_1255), .B2(n_1278), .Y(n_1277) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_147), .A2(n_153), .B1(n_386), .B2(n_501), .Y(n_700) );
INVxp67_ASAP7_75t_SL g728 ( .A(n_147), .Y(n_728) );
INVx1_ASAP7_75t_L g1141 ( .A(n_148), .Y(n_1141) );
INVx1_ASAP7_75t_L g511 ( .A(n_149), .Y(n_511) );
INVx1_ASAP7_75t_L g612 ( .A(n_150), .Y(n_612) );
INVx1_ASAP7_75t_L g659 ( .A(n_151), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_151), .A2(n_219), .B1(n_509), .B2(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g1455 ( .A(n_152), .Y(n_1455) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_153), .Y(n_725) );
AOI221xp5_ASAP7_75t_SL g1055 ( .A1(n_154), .A2(n_175), .B1(n_657), .B2(n_954), .C(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1082 ( .A(n_154), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_155), .A2(n_211), .B1(n_1061), .B2(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_155), .A2(n_261), .B1(n_355), .B2(n_509), .Y(n_1174) );
BUFx3_ASAP7_75t_L g322 ( .A(n_157), .Y(n_322) );
INVx1_ASAP7_75t_L g1091 ( .A(n_158), .Y(n_1091) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_159), .Y(n_797) );
INVx1_ASAP7_75t_L g498 ( .A(n_160), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_161), .A2(n_195), .B1(n_466), .B2(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_162), .A2(n_203), .B1(n_583), .B2(n_586), .C(n_587), .Y(n_582) );
INVx1_ASAP7_75t_L g317 ( .A(n_163), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_164), .B(n_546), .Y(n_1225) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_165), .A2(n_239), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
INVx1_ASAP7_75t_L g706 ( .A(n_166), .Y(n_706) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_167), .Y(n_904) );
INVx1_ASAP7_75t_L g663 ( .A(n_168), .Y(n_663) );
INVx1_ASAP7_75t_L g1204 ( .A(n_169), .Y(n_1204) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_170), .Y(n_304) );
INVx1_ASAP7_75t_L g942 ( .A(n_171), .Y(n_942) );
INVx1_ASAP7_75t_L g1153 ( .A(n_172), .Y(n_1153) );
AOI22xp33_ASAP7_75t_SL g1568 ( .A1(n_173), .A2(n_267), .B1(n_1569), .B2(n_1570), .Y(n_1568) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_174), .A2(n_212), .B1(n_642), .B2(n_646), .Y(n_1166) );
INVx1_ASAP7_75t_L g1088 ( .A(n_175), .Y(n_1088) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_177), .A2(n_355), .B(n_357), .Y(n_354) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_177), .Y(n_431) );
OAI222xp33_ASAP7_75t_L g862 ( .A1(n_178), .A2(n_214), .B1(n_240), .B2(n_863), .C1(n_866), .C2(n_868), .Y(n_862) );
OAI211xp5_ASAP7_75t_L g872 ( .A1(n_178), .A2(n_873), .B(n_876), .C(n_885), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g1053 ( .A(n_179), .Y(n_1053) );
INVx1_ASAP7_75t_L g637 ( .A(n_180), .Y(n_637) );
INVx1_ASAP7_75t_L g1228 ( .A(n_181), .Y(n_1228) );
INVx1_ASAP7_75t_L g986 ( .A(n_182), .Y(n_986) );
OAI221xp5_ASAP7_75t_L g1014 ( .A1(n_182), .A2(n_537), .B1(n_1015), .B2(n_1021), .C(n_1022), .Y(n_1014) );
INVx1_ASAP7_75t_L g1092 ( .A(n_183), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_184), .A2(n_207), .B1(n_457), .B2(n_466), .C(n_470), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_185), .A2(n_211), .B1(n_509), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g925 ( .A(n_186), .Y(n_925) );
AOI22xp5_ASAP7_75t_SL g1269 ( .A1(n_187), .A2(n_266), .B1(n_1255), .B2(n_1260), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_189), .A2(n_193), .B1(n_1249), .B2(n_1255), .Y(n_1339) );
INVx1_ASAP7_75t_L g1085 ( .A(n_190), .Y(n_1085) );
INVx1_ASAP7_75t_L g391 ( .A(n_192), .Y(n_391) );
INVx1_ASAP7_75t_L g513 ( .A(n_194), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g977 ( .A(n_196), .Y(n_977) );
INVx1_ASAP7_75t_L g738 ( .A(n_197), .Y(n_738) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_198), .Y(n_303) );
INVx1_ASAP7_75t_L g366 ( .A(n_199), .Y(n_366) );
XNOR2x1_ASAP7_75t_L g494 ( .A(n_200), .B(n_495), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g1115 ( .A(n_201), .Y(n_1115) );
INVx1_ASAP7_75t_L g708 ( .A(n_202), .Y(n_708) );
INVx1_ASAP7_75t_L g610 ( .A(n_203), .Y(n_610) );
INVx1_ASAP7_75t_L g598 ( .A(n_204), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g331 ( .A1(n_207), .A2(n_236), .B1(n_332), .B2(n_337), .C(n_343), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g1557 ( .A1(n_208), .A2(n_267), .B1(n_508), .B2(n_1549), .Y(n_1557) );
INVx1_ASAP7_75t_L g773 ( .A(n_209), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g1521 ( .A1(n_210), .A2(n_268), .B1(n_355), .B2(n_703), .C(n_1522), .Y(n_1521) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_213), .A2(n_281), .B1(n_1476), .B2(n_1477), .Y(n_1475) );
OAI22xp5_ASAP7_75t_L g1496 ( .A1(n_213), .A2(n_281), .B1(n_1497), .B2(n_1498), .Y(n_1496) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_215), .A2(n_245), .B1(n_853), .B2(n_855), .Y(n_852) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_216), .A2(n_533), .B(n_667), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_216), .A2(n_233), .B1(n_386), .B2(n_501), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g1229 ( .A1(n_217), .A2(n_732), .B(n_801), .Y(n_1229) );
INVx1_ASAP7_75t_L g632 ( .A(n_218), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_219), .A2(n_256), .B1(n_482), .B2(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g698 ( .A(n_220), .Y(n_698) );
INVx1_ASAP7_75t_L g1561 ( .A(n_222), .Y(n_1561) );
AOI21xp33_ASAP7_75t_L g1207 ( .A1(n_223), .A2(n_1208), .B(n_1211), .Y(n_1207) );
INVx1_ASAP7_75t_L g973 ( .A(n_224), .Y(n_973) );
INVxp67_ASAP7_75t_SL g978 ( .A(n_225), .Y(n_978) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_225), .A2(n_343), .B1(n_386), .B2(n_994), .C(n_999), .Y(n_993) );
INVx1_ASAP7_75t_L g1101 ( .A(n_226), .Y(n_1101) );
INVx1_ASAP7_75t_L g693 ( .A(n_227), .Y(n_693) );
INVx1_ASAP7_75t_L g1458 ( .A(n_228), .Y(n_1458) );
INVx1_ASAP7_75t_L g1544 ( .A(n_229), .Y(n_1544) );
BUFx3_ASAP7_75t_L g307 ( .A(n_230), .Y(n_307) );
INVx1_ASAP7_75t_L g416 ( .A(n_230), .Y(n_416) );
INVx1_ASAP7_75t_L g967 ( .A(n_231), .Y(n_967) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_232), .Y(n_531) );
INVxp33_ASAP7_75t_L g665 ( .A(n_233), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g991 ( .A1(n_234), .A2(n_379), .B(n_853), .Y(n_991) );
INVx1_ASAP7_75t_L g1010 ( .A(n_234), .Y(n_1010) );
INVx1_ASAP7_75t_L g673 ( .A(n_235), .Y(n_673) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_236), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1507 ( .A1(n_237), .A2(n_268), .B1(n_822), .B2(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g998 ( .A(n_239), .Y(n_998) );
CKINVDCx5p33_ASAP7_75t_R g983 ( .A(n_241), .Y(n_983) );
INVx2_ASAP7_75t_L g404 ( .A(n_242), .Y(n_404) );
INVx1_ASAP7_75t_L g413 ( .A(n_242), .Y(n_413) );
INVx1_ASAP7_75t_L g476 ( .A(n_242), .Y(n_476) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_243), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_244), .A2(n_256), .B1(n_357), .B2(n_677), .C(n_679), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_245), .A2(n_247), .B1(n_546), .B2(n_801), .C(n_906), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_246), .A2(n_258), .B1(n_382), .B2(n_383), .Y(n_381) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_246), .Y(n_451) );
INVx1_ASAP7_75t_L g1564 ( .A(n_248), .Y(n_1564) );
INVx1_ASAP7_75t_L g1221 ( .A(n_249), .Y(n_1221) );
INVxp67_ASAP7_75t_SL g726 ( .A(n_250), .Y(n_726) );
INVx1_ASAP7_75t_L g839 ( .A(n_251), .Y(n_839) );
XOR2x2_ASAP7_75t_L g1190 ( .A(n_252), .B(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_253), .A2(n_260), .B1(n_1252), .B2(n_1255), .Y(n_1251) );
XNOR2xp5_ASAP7_75t_L g1451 ( .A(n_253), .B(n_1452), .Y(n_1451) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_253), .A2(n_1528), .B1(n_1531), .B2(n_1582), .Y(n_1527) );
CKINVDCx5p33_ASAP7_75t_R g988 ( .A(n_255), .Y(n_988) );
INVx1_ASAP7_75t_L g350 ( .A(n_257), .Y(n_350) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_258), .Y(n_428) );
INVx1_ASAP7_75t_L g1154 ( .A(n_259), .Y(n_1154) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_262), .B(n_1024), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_263), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1464 ( .A(n_264), .Y(n_1464) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_265), .Y(n_792) );
INVx1_ASAP7_75t_L g831 ( .A(n_269), .Y(n_831) );
XNOR2xp5_ASAP7_75t_L g826 ( .A(n_270), .B(n_827), .Y(n_826) );
NAND2xp33_ASAP7_75t_SL g579 ( .A(n_271), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g618 ( .A(n_271), .Y(n_618) );
INVxp67_ASAP7_75t_SL g1145 ( .A(n_272), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g1041 ( .A(n_273), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_275), .A2(n_279), .B1(n_933), .B2(n_934), .C(n_938), .Y(n_932) );
INVx1_ASAP7_75t_L g985 ( .A(n_276), .Y(n_985) );
INVx1_ASAP7_75t_L g1066 ( .A(n_278), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g950 ( .A(n_279), .Y(n_950) );
INVx1_ASAP7_75t_L g575 ( .A(n_280), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_308), .B(n_1237), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1526 ( .A(n_287), .B(n_296), .Y(n_1526) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1530 ( .A(n_289), .B(n_292), .Y(n_1530) );
INVx1_ASAP7_75t_L g1583 ( .A(n_289), .Y(n_1583) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g1586 ( .A(n_292), .B(n_1583), .Y(n_1586) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g1479 ( .A(n_296), .B(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g454 ( .A(n_297), .B(n_307), .Y(n_454) );
AND2x4_ASAP7_75t_L g907 ( .A(n_297), .B(n_306), .Y(n_907) );
AND2x4_ASAP7_75t_SL g1525 ( .A(n_298), .B(n_1526), .Y(n_1525) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_300), .B(n_305), .Y(n_299) );
INVxp67_ASAP7_75t_L g551 ( .A(n_300), .Y(n_551) );
BUFx4f_ASAP7_75t_L g556 ( .A(n_300), .Y(n_556) );
INVx1_ASAP7_75t_L g661 ( .A(n_300), .Y(n_661) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_300), .B(n_1460), .Y(n_1476) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g430 ( .A(n_301), .Y(n_430) );
BUFx4f_ASAP7_75t_L g742 ( .A(n_301), .Y(n_742) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g418 ( .A(n_303), .Y(n_418) );
INVx2_ASAP7_75t_L g435 ( .A(n_303), .Y(n_435) );
NAND2x1_ASAP7_75t_L g443 ( .A(n_303), .B(n_304), .Y(n_443) );
INVx1_ASAP7_75t_L g469 ( .A(n_303), .Y(n_469) );
AND2x2_ASAP7_75t_L g492 ( .A(n_303), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g545 ( .A(n_303), .B(n_304), .Y(n_545) );
INVx1_ASAP7_75t_L g419 ( .A(n_304), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_304), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g440 ( .A(n_304), .B(n_418), .Y(n_440) );
BUFx2_ASAP7_75t_L g465 ( .A(n_304), .Y(n_465) );
AND2x2_ASAP7_75t_L g484 ( .A(n_304), .B(n_435), .Y(n_484) );
INVx2_ASAP7_75t_L g493 ( .A(n_304), .Y(n_493) );
OR2x6_ASAP7_75t_L g1457 ( .A(n_305), .B(n_430), .Y(n_1457) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g1466 ( .A(n_306), .Y(n_1466) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g1468 ( .A(n_307), .B(n_468), .Y(n_1468) );
XOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_757), .Y(n_308) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_628), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_566), .B1(n_626), .B2(n_627), .Y(n_310) );
INVx1_ASAP7_75t_L g626 ( .A(n_311), .Y(n_626) );
OA22x2_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_494), .B1(n_564), .B2(n_565), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_SL g565 ( .A(n_313), .Y(n_565) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_420), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_384), .B(n_401), .C(n_405), .Y(n_315) );
AOI211xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_331), .C(n_348), .Y(n_316) );
AOI222xp33_ASAP7_75t_L g472 ( .A1(n_317), .A2(n_393), .B1(n_473), .B2(n_479), .C1(n_485), .C2(n_487), .Y(n_472) );
AOI211xp5_ASAP7_75t_L g497 ( .A1(n_318), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
AOI211xp5_ASAP7_75t_SL g602 ( .A1(n_318), .A2(n_598), .B(n_603), .C(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g689 ( .A(n_318), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g697 ( .A1(n_318), .A2(n_698), .B(n_699), .C(n_700), .Y(n_697) );
AOI211xp5_ASAP7_75t_SL g766 ( .A1(n_318), .A2(n_767), .B(n_768), .C(n_769), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_318), .A2(n_929), .B1(n_932), .B2(n_942), .Y(n_928) );
AOI211xp5_ASAP7_75t_SL g1193 ( .A1(n_318), .A2(n_1194), .B(n_1195), .C(n_1196), .Y(n_1193) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x6_ASAP7_75t_L g868 ( .A(n_319), .B(n_869), .Y(n_868) );
OR2x2_ASAP7_75t_L g975 ( .A(n_319), .B(n_869), .Y(n_975) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_320), .B(n_326), .Y(n_319) );
INVx8_ASAP7_75t_L g356 ( .A(n_320), .Y(n_356) );
BUFx3_ASAP7_75t_L g382 ( .A(n_320), .Y(n_382) );
AND2x2_ASAP7_75t_L g396 ( .A(n_320), .B(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g507 ( .A(n_320), .Y(n_507) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
AND2x4_ASAP7_75t_L g364 ( .A(n_321), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_322), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_322), .B(n_342), .Y(n_371) );
AND2x4_ASAP7_75t_L g400 ( .A(n_322), .B(n_341), .Y(n_400) );
OR2x2_ASAP7_75t_L g525 ( .A(n_322), .B(n_324), .Y(n_525) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g365 ( .A(n_325), .Y(n_365) );
AND2x6_ASAP7_75t_L g333 ( .A(n_326), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g338 ( .A(n_326), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g347 ( .A(n_326), .Y(n_347) );
AND2x4_ASAP7_75t_L g833 ( .A(n_326), .B(n_475), .Y(n_833) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_327), .B(n_360), .Y(n_359) );
NAND3x1_ASAP7_75t_L g857 ( .A(n_327), .B(n_360), .C(n_858), .Y(n_857) );
OR2x4_ASAP7_75t_L g1484 ( .A(n_327), .B(n_525), .Y(n_1484) );
INVx1_ASAP7_75t_L g1486 ( .A(n_327), .Y(n_1486) );
OR2x6_ASAP7_75t_L g1498 ( .A(n_327), .B(n_937), .Y(n_1498) );
AND2x4_ASAP7_75t_L g1499 ( .A(n_327), .B(n_400), .Y(n_1499) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_328), .B(n_330), .Y(n_380) );
BUFx3_ASAP7_75t_L g515 ( .A(n_328), .Y(n_515) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g514 ( .A(n_330), .B(n_515), .Y(n_514) );
AND3x4_ASAP7_75t_L g847 ( .A(n_330), .B(n_403), .C(n_515), .Y(n_847) );
HB1xp67_ASAP7_75t_L g1503 ( .A(n_330), .Y(n_1503) );
INVx4_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_333), .A2(n_338), .B1(n_637), .B2(n_663), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_333), .A2(n_338), .B1(n_925), .B2(n_926), .C(n_927), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_333), .A2(n_338), .B1(n_985), .B2(n_986), .Y(n_984) );
AND2x2_ASAP7_75t_L g832 ( .A(n_334), .B(n_833), .Y(n_832) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_336), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g383 ( .A(n_336), .B(n_340), .Y(n_383) );
BUFx2_ASAP7_75t_L g1495 ( .A(n_336), .Y(n_1495) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_338), .Y(n_1172) );
INVx1_ASAP7_75t_L g837 ( .A(n_339), .Y(n_837) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g346 ( .A(n_342), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_343), .Y(n_927) );
OR2x6_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
INVx1_ASAP7_75t_L g683 ( .A(n_344), .Y(n_683) );
INVx1_ASAP7_75t_L g1210 ( .A(n_344), .Y(n_1210) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_345), .Y(n_353) );
BUFx3_ASAP7_75t_L g717 ( .A(n_345), .Y(n_717) );
BUFx2_ASAP7_75t_L g1492 ( .A(n_346), .Y(n_1492) );
INVx1_ASAP7_75t_L g1109 ( .A(n_347), .Y(n_1109) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_361), .B(n_373), .Y(n_348) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B(n_354), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_350), .A2(n_374), .B1(n_445), .B2(n_446), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_351), .A2(n_514), .B1(n_1128), .B2(n_1129), .C(n_1130), .Y(n_1127) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g611 ( .A(n_352), .Y(n_611) );
INVx1_ASAP7_75t_L g1119 ( .A(n_352), .Y(n_1119) );
INVx2_ASAP7_75t_L g1202 ( .A(n_352), .Y(n_1202) );
INVx4_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g376 ( .A(n_353), .Y(n_376) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_353), .Y(n_778) );
OR2x2_ASAP7_75t_L g867 ( .A(n_353), .B(n_842), .Y(n_867) );
BUFx6f_ASAP7_75t_L g1080 ( .A(n_353), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_355), .A2(n_916), .B1(n_977), .B2(n_983), .Y(n_982) );
A2O1A1Ixp33_ASAP7_75t_L g1072 ( .A1(n_355), .A2(n_833), .B(n_1041), .C(n_1073), .Y(n_1072) );
INVx8_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g679 ( .A(n_356), .Y(n_679) );
INVx2_ASAP7_75t_L g849 ( .A(n_356), .Y(n_849) );
INVx3_ASAP7_75t_L g1107 ( .A(n_356), .Y(n_1107) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_358), .A2(n_375), .B1(n_523), .B2(n_524), .C(n_526), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_358), .A2(n_610), .B1(n_611), .B2(n_612), .C(n_613), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_358), .A2(n_717), .B1(n_718), .B2(n_719), .C(n_720), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_358), .B(n_789), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g994 ( .A1(n_358), .A2(n_613), .B1(n_995), .B2(n_997), .C(n_998), .Y(n_994) );
OAI221xp5_ASAP7_75t_L g1117 ( .A1(n_358), .A2(n_524), .B1(n_1118), .B2(n_1119), .C(n_1120), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_358), .B(n_1212), .Y(n_1211) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_359), .B(n_425), .Y(n_1093) );
OR2x6_ASAP7_75t_L g1519 ( .A(n_359), .B(n_425), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B1(n_367), .B2(n_372), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_362), .A2(n_514), .B1(n_592), .B2(n_611), .C(n_618), .Y(n_617) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g512 ( .A(n_363), .Y(n_512) );
INVx3_ASAP7_75t_L g705 ( .A(n_363), .Y(n_705) );
AND2x4_ASAP7_75t_L g844 ( .A(n_363), .B(n_841), .Y(n_844) );
INVx3_ASAP7_75t_L g854 ( .A(n_363), .Y(n_854) );
BUFx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_364), .Y(n_378) );
INVx2_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_364), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_366), .A2(n_437), .B1(n_438), .B2(n_441), .Y(n_436) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g864 ( .A(n_369), .B(n_842), .Y(n_864) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_370), .Y(n_675) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g937 ( .A(n_371), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_372), .A2(n_432), .B1(n_449), .B2(n_451), .Y(n_448) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_377), .C(n_381), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_375), .A2(n_511), .B1(n_512), .B2(n_513), .C(n_514), .Y(n_510) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g990 ( .A(n_376), .Y(n_990) );
INVx2_ASAP7_75t_SL g918 ( .A(n_378), .Y(n_918) );
INVx2_ASAP7_75t_SL g921 ( .A(n_378), .Y(n_921) );
INVx3_ASAP7_75t_L g933 ( .A(n_378), .Y(n_933) );
INVx5_ASAP7_75t_L g1083 ( .A(n_378), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_378), .Y(n_1114) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_380), .B(n_455), .Y(n_1076) );
BUFx2_ASAP7_75t_L g923 ( .A(n_382), .Y(n_923) );
AND2x4_ASAP7_75t_L g392 ( .A(n_383), .B(n_388), .Y(n_392) );
BUFx12f_ASAP7_75t_L g509 ( .A(n_383), .Y(n_509) );
INVx5_ASAP7_75t_L g521 ( .A(n_383), .Y(n_521) );
BUFx2_ASAP7_75t_L g608 ( .A(n_383), .Y(n_608) );
BUFx3_ASAP7_75t_L g715 ( .A(n_383), .Y(n_715) );
BUFx3_ASAP7_75t_L g782 ( .A(n_383), .Y(n_782) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_391), .B1(n_392), .B2(n_393), .C(n_394), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
OR2x6_ASAP7_75t_SL g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_388), .Y(n_931) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g397 ( .A(n_389), .Y(n_397) );
OR2x2_ASAP7_75t_L g842 ( .A(n_389), .B(n_455), .Y(n_842) );
INVx3_ASAP7_75t_L g672 ( .A(n_390), .Y(n_672) );
BUFx2_ASAP7_75t_L g1550 ( .A(n_390), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_391), .B(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g501 ( .A(n_392), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_392), .B(n_529), .Y(n_1026) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_396), .A2(n_399), .B1(n_632), .B2(n_639), .Y(n_687) );
AND2x2_ASAP7_75t_L g399 ( .A(n_397), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g678 ( .A(n_400), .Y(n_678) );
BUFx3_ASAP7_75t_L g703 ( .A(n_400), .Y(n_703) );
BUFx2_ASAP7_75t_L g861 ( .A(n_400), .Y(n_861) );
BUFx2_ASAP7_75t_L g916 ( .A(n_400), .Y(n_916) );
BUFx2_ASAP7_75t_L g941 ( .A(n_400), .Y(n_941) );
INVx1_ASAP7_75t_L g621 ( .A(n_401), .Y(n_621) );
INVx1_ASAP7_75t_L g1002 ( .A(n_401), .Y(n_1002) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_402), .Y(n_790) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g1167 ( .A1(n_403), .A2(n_1168), .B1(n_1185), .B2(n_1187), .Y(n_1167) );
INVx2_ASAP7_75t_SL g1213 ( .A(n_403), .Y(n_1213) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g425 ( .A(n_404), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_404), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_409), .B(n_563), .Y(n_562) );
AOI211x1_ASAP7_75t_L g631 ( .A1(n_409), .A2(n_632), .B(n_633), .C(n_666), .Y(n_631) );
AO211x2_ASAP7_75t_L g763 ( .A1(n_409), .A2(n_764), .B(n_765), .C(n_793), .Y(n_763) );
AOI222xp33_ASAP7_75t_L g972 ( .A1(n_409), .A2(n_489), .B1(n_973), .B2(n_974), .C1(n_977), .C2(n_978), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g1140 ( .A1(n_409), .A2(n_489), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_409), .B(n_1149), .Y(n_1148) );
AOI211xp5_ASAP7_75t_L g1217 ( .A1(n_409), .A2(n_1218), .B(n_1219), .C(n_1223), .Y(n_1217) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
AND2x4_ASAP7_75t_L g489 ( .A(n_410), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g466 ( .A(n_411), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g572 ( .A(n_411), .B(n_467), .Y(n_572) );
INVxp67_ASAP7_75t_L g869 ( .A(n_411), .Y(n_869) );
INVx1_ASAP7_75t_L g1480 ( .A(n_411), .Y(n_1480) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g887 ( .A(n_414), .Y(n_887) );
BUFx6f_ASAP7_75t_L g1563 ( .A(n_414), .Y(n_1563) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_415), .B(n_476), .Y(n_481) );
AND2x2_ASAP7_75t_L g490 ( .A(n_415), .B(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_L g874 ( .A(n_415), .B(n_875), .Y(n_874) );
AND2x4_ASAP7_75t_L g890 ( .A(n_415), .B(n_491), .Y(n_890) );
AND2x4_ASAP7_75t_SL g895 ( .A(n_415), .B(n_656), .Y(n_895) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_415), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1460 ( .A(n_416), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_417), .B(n_462), .Y(n_478) );
INVx3_ASAP7_75t_L g649 ( .A(n_417), .Y(n_649) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_417), .Y(n_964) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_472), .C(n_488), .Y(n_420) );
NOR2xp33_ASAP7_75t_SL g421 ( .A(n_422), .B(n_456), .Y(n_421) );
OAI33xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .A3(n_436), .B1(n_444), .B2(n_448), .B3(n_452), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_424), .Y(n_552) );
INVx4_ASAP7_75t_L g596 ( .A(n_424), .Y(n_596) );
INVx2_ASAP7_75t_L g652 ( .A(n_424), .Y(n_652) );
INVx2_ASAP7_75t_L g732 ( .A(n_424), .Y(n_732) );
AOI31xp33_ASAP7_75t_L g1156 ( .A1(n_424), .A2(n_570), .A3(n_1157), .B(n_1158), .Y(n_1156) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g529 ( .A(n_425), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_431), .B2(n_432), .Y(n_427) );
INVx2_ASAP7_75t_L g586 ( .A(n_429), .Y(n_586) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g450 ( .A(n_430), .Y(n_450) );
BUFx3_ASAP7_75t_L g752 ( .A(n_430), .Y(n_752) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_430), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_432), .A2(n_526), .B1(n_549), .B2(n_550), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_432), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_554) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx8_ASAP7_75t_L g578 ( .A(n_433), .Y(n_578) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_433), .B(n_1466), .Y(n_1477) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_438), .A2(n_903), .B1(n_1115), .B2(n_1128), .C(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g445 ( .A(n_440), .Y(n_445) );
BUFx3_ASAP7_75t_L g581 ( .A(n_440), .Y(n_581) );
BUFx2_ASAP7_75t_L g736 ( .A(n_440), .Y(n_736) );
INVx2_ASAP7_75t_L g747 ( .A(n_440), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_441), .A2(n_1112), .B1(n_1122), .B2(n_1134), .Y(n_1133) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g486 ( .A(n_442), .B(n_481), .Y(n_486) );
OR2x2_ASAP7_75t_L g537 ( .A(n_442), .B(n_481), .Y(n_537) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_443), .Y(n_447) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g470 ( .A(n_447), .B(n_471), .Y(n_470) );
INVx4_ASAP7_75t_L g585 ( .A(n_447), .Y(n_585) );
BUFx4f_ASAP7_75t_L g589 ( .A(n_447), .Y(n_589) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_447), .Y(n_737) );
BUFx4f_ASAP7_75t_L g1017 ( .A(n_447), .Y(n_1017) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g750 ( .A(n_453), .Y(n_750) );
AOI33xp33_ASAP7_75t_L g1506 ( .A1(n_453), .A2(n_805), .A3(n_1507), .B1(n_1509), .B2(n_1511), .B3(n_1512), .Y(n_1506) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x4_ASAP7_75t_L g558 ( .A(n_454), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_454), .B(n_559), .Y(n_587) );
INVx4_ASAP7_75t_L g882 ( .A(n_454), .Y(n_882) );
INVx4_ASAP7_75t_L g1059 ( .A(n_454), .Y(n_1059) );
INVx1_ASAP7_75t_L g560 ( .A(n_455), .Y(n_560) );
HB1xp67_ASAP7_75t_L g1505 ( .A(n_455), .Y(n_1505) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_459), .Y(n_539) );
INVx1_ASAP7_75t_L g636 ( .A(n_459), .Y(n_636) );
NAND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_463), .Y(n_459) );
INVx1_ASAP7_75t_L g471 ( .A(n_460), .Y(n_471) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_462), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g884 ( .A(n_462), .B(n_656), .Y(n_884) );
INVx1_ASAP7_75t_L g899 ( .A(n_462), .Y(n_899) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_462), .B(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g898 ( .A(n_465), .Y(n_898) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_465), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_465), .B(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1052 ( .A(n_467), .Y(n_1052) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_470), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g959 ( .A1(n_470), .A2(n_651), .B(n_960), .Y(n_959) );
OAI21xp5_ASAP7_75t_SL g1004 ( .A1(n_470), .A2(n_1005), .B(n_1008), .Y(n_1004) );
OAI21xp5_ASAP7_75t_L g1135 ( .A1(n_470), .A2(n_1021), .B(n_1136), .Y(n_1135) );
AOI222xp33_ASAP7_75t_L g540 ( .A1(n_473), .A2(n_541), .B1(n_552), .B2(n_553), .C1(n_558), .C2(n_561), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g597 ( .A1(n_473), .A2(n_479), .B1(n_485), .B2(n_598), .C1(n_599), .C2(n_600), .Y(n_597) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_473), .A2(n_570), .B(n_665), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g724 ( .A1(n_473), .A2(n_479), .B1(n_485), .B2(n_698), .C1(n_725), .C2(n_726), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g823 ( .A1(n_473), .A2(n_570), .B(n_824), .Y(n_823) );
AOI322xp5_ASAP7_75t_L g1224 ( .A1(n_473), .A2(n_558), .A3(n_1225), .B1(n_1226), .B2(n_1229), .C1(n_1230), .C2(n_1231), .Y(n_1224) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_477), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g865 ( .A(n_475), .B(n_478), .Y(n_865) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g858 ( .A(n_476), .Y(n_858) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI211xp5_ASAP7_75t_L g535 ( .A1(n_479), .A2(n_498), .B(n_536), .C(n_538), .Y(n_535) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_479), .A2(n_635), .B1(n_636), .B2(n_637), .C1(n_638), .C2(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g796 ( .A(n_479), .Y(n_796) );
INVxp67_ASAP7_75t_L g948 ( .A(n_479), .Y(n_948) );
INVx1_ASAP7_75t_L g976 ( .A(n_479), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_479), .A2(n_485), .B1(n_1153), .B2(n_1154), .Y(n_1152) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g1508 ( .A(n_483), .Y(n_1508) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g821 ( .A(n_484), .Y(n_821) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_484), .Y(n_875) );
BUFx3_ASAP7_75t_L g965 ( .A(n_484), .Y(n_965) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_485), .A2(n_558), .A3(n_641), .B1(n_647), .B2(n_650), .C1(n_653), .C2(n_663), .Y(n_640) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g533 ( .A(n_489), .Y(n_533) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_489), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_489), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_489), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g1186 ( .A(n_489), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_489), .B(n_1215), .Y(n_1214) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_491), .Y(n_547) );
INVx2_ASAP7_75t_L g810 ( .A(n_491), .Y(n_810) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g645 ( .A(n_492), .Y(n_645) );
BUFx3_ASAP7_75t_L g819 ( .A(n_492), .Y(n_819) );
AND2x4_ASAP7_75t_L g1459 ( .A(n_492), .B(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g564 ( .A(n_494), .Y(n_564) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_534), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_502), .B(n_527), .C(n_530), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_516), .C(n_517), .Y(n_502) );
BUFx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g1203 ( .A1(n_506), .A2(n_514), .B1(n_521), .B2(n_1204), .C(n_1205), .Y(n_1203) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
BUFx3_ASAP7_75t_L g686 ( .A(n_507), .Y(n_686) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_512), .A2(n_674), .B1(n_1000), .B2(n_1001), .Y(n_999) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_514), .A2(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g780 ( .A(n_514), .Y(n_780) );
INVx3_ASAP7_75t_L g1491 ( .A(n_515), .Y(n_1491) );
INVx2_ASAP7_75t_L g1129 ( .A(n_518), .Y(n_1129) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_519), .Y(n_607) );
INVx2_ASAP7_75t_L g714 ( .A(n_519), .Y(n_714) );
INVx2_ASAP7_75t_L g1182 ( .A(n_519), .Y(n_1182) );
INVx1_ASAP7_75t_L g1200 ( .A(n_519), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_519), .B(n_1486), .Y(n_1485) );
INVx2_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g851 ( .A(n_521), .Y(n_851) );
INVx2_ASAP7_75t_L g855 ( .A(n_521), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_524), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx4f_ASAP7_75t_L g615 ( .A(n_525), .Y(n_615) );
BUFx3_ASAP7_75t_L g719 ( .A(n_525), .Y(n_719) );
INVx2_ASAP7_75t_L g1125 ( .A(n_525), .Y(n_1125) );
OR2x4_ASAP7_75t_L g1497 ( .A(n_525), .B(n_1486), .Y(n_1497) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g722 ( .A(n_528), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g911 ( .A1(n_528), .A2(n_912), .B(n_943), .Y(n_911) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g692 ( .A(n_529), .Y(n_692) );
AOI21xp5_ASAP7_75t_SL g1037 ( .A1(n_529), .A2(n_1038), .B(n_1054), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .C(n_562), .Y(n_534) );
INVx1_ASAP7_75t_L g879 ( .A(n_542), .Y(n_879) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g646 ( .A(n_543), .Y(n_646) );
INVx1_ASAP7_75t_L g1473 ( .A(n_543), .Y(n_1473) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g1471 ( .A(n_544), .Y(n_1471) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_545), .Y(n_656) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI211x1_ASAP7_75t_L g1131 ( .A1(n_552), .A2(n_1132), .B(n_1135), .C(n_1138), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_556), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_556), .A2(n_814), .B1(n_1205), .B2(n_1228), .Y(n_1227) );
AOI211xp5_ASAP7_75t_L g951 ( .A1(n_558), .A2(n_952), .B(n_959), .C(n_966), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_558), .Y(n_1021) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_558), .B(n_1163), .C(n_1166), .Y(n_1162) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g627 ( .A(n_566), .Y(n_627) );
XOR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_625), .Y(n_566) );
NOR2x1_ASAP7_75t_SL g567 ( .A(n_568), .B(n_601), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .C(n_573), .Y(n_569) );
OR3x1_ASAP7_75t_L g729 ( .A(n_570), .B(n_730), .C(n_731), .Y(n_729) );
INVx2_ASAP7_75t_SL g638 ( .A(n_572), .Y(n_638) );
AND2x4_ASAP7_75t_L g866 ( .A(n_572), .B(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_588), .Y(n_573) );
OAI211xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_579), .C(n_582), .Y(n_574) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_577), .A2(n_659), .B1(n_660), .B2(n_662), .Y(n_658) );
INVx4_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g595 ( .A(n_578), .Y(n_595) );
INVx2_ASAP7_75t_L g743 ( .A(n_578), .Y(n_743) );
INVx2_ASAP7_75t_SL g753 ( .A(n_578), .Y(n_753) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_578), .Y(n_815) );
INVx3_ASAP7_75t_L g591 ( .A(n_580), .Y(n_591) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_584), .A2(n_591), .B1(n_961), .B2(n_962), .C(n_963), .Y(n_960) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g749 ( .A(n_585), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_591), .B2(n_592), .C(n_593), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_589), .A2(n_1000), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1008) );
INVxp33_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g805 ( .A(n_596), .Y(n_805) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_596), .Y(n_1007) );
A2O1A1Ixp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_605), .B(n_620), .C(n_622), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_616), .C(n_619), .Y(n_605) );
INVx1_ASAP7_75t_L g774 ( .A(n_607), .Y(n_774) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g1077 ( .A1(n_615), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1077) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_615), .A2(n_717), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_620), .A2(n_872), .B(n_891), .Y(n_871) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_624), .B(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_694), .B1(n_755), .B2(n_756), .Y(n_629) );
INVx1_ASAP7_75t_L g755 ( .A(n_630), .Y(n_755) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_693), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_640), .C(n_664), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g794 ( .A1(n_636), .A2(n_638), .B1(n_767), .B2(n_795), .C1(n_797), .C2(n_798), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_636), .A2(n_638), .B1(n_983), .B2(n_985), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g1159 ( .A1(n_636), .A2(n_638), .B1(n_1160), .B2(n_1161), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_636), .A2(n_638), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g657 ( .A(n_643), .Y(n_657) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g953 ( .A(n_645), .Y(n_953) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_SL g822 ( .A(n_649), .Y(n_822) );
INVx2_ASAP7_75t_L g1012 ( .A(n_649), .Y(n_1012) );
INVx1_ASAP7_75t_L g1513 ( .A(n_649), .Y(n_1513) );
INVx2_ASAP7_75t_L g1569 ( .A(n_649), .Y(n_1569) );
INVx1_ASAP7_75t_L g1574 ( .A(n_649), .Y(n_1574) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
BUFx3_ASAP7_75t_L g801 ( .A(n_656), .Y(n_801) );
BUFx3_ASAP7_75t_L g817 ( .A(n_656), .Y(n_817) );
BUFx3_ASAP7_75t_L g954 ( .A(n_656), .Y(n_954) );
BUFx6f_ASAP7_75t_L g1233 ( .A(n_656), .Y(n_1233) );
BUFx3_ASAP7_75t_L g1576 ( .A(n_656), .Y(n_1576) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_662), .A2(n_671), .B1(n_673), .B2(n_674), .C(n_676), .Y(n_670) );
OAI31xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .A3(n_688), .B(n_691), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_680), .C(n_687), .Y(n_669) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_672), .B(n_1068), .Y(n_1067) );
INVx2_ASAP7_75t_L g1087 ( .A(n_672), .Y(n_1087) );
CKINVDCx8_ASAP7_75t_R g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g709 ( .A(n_675), .Y(n_709) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g1102 ( .A(n_678), .Y(n_1102) );
INVx2_ASAP7_75t_L g1517 ( .A(n_678), .Y(n_1517) );
AND2x4_ASAP7_75t_L g840 ( .A(n_679), .B(n_841), .Y(n_840) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B(n_684), .C(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g1184 ( .A(n_689), .Y(n_1184) );
OAI21x1_ASAP7_75t_L g1096 ( .A1(n_691), .A2(n_1097), .B(n_1110), .Y(n_1096) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g756 ( .A(n_694), .Y(n_756) );
AOI211x1_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_721), .B(n_723), .C(n_729), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_701), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_711), .C(n_712), .Y(n_701) );
INVx1_ASAP7_75t_L g1179 ( .A(n_705), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_706), .A2(n_734), .B1(n_737), .B2(n_738), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_708), .A2(n_720), .B1(n_740), .B2(n_743), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_710), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_SL g1100 ( .A1(n_715), .A2(n_1101), .B1(n_1102), .B2(n_1103), .C(n_1104), .Y(n_1100) );
INVx2_ASAP7_75t_L g996 ( .A(n_717), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_718), .A2(n_745), .B1(n_748), .B2(n_749), .Y(n_744) );
INVx1_ASAP7_75t_L g787 ( .A(n_719), .Y(n_787) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g1558 ( .A1(n_722), .A2(n_1559), .B(n_1580), .Y(n_1558) );
OAI33xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .A3(n_739), .B1(n_744), .B2(n_750), .B3(n_751), .Y(n_731) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g1016 ( .A(n_735), .Y(n_1016) );
INVx4_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g901 ( .A(n_741), .Y(n_901) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_L g957 ( .A(n_742), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_743), .A2(n_752), .B1(n_1204), .B2(n_1235), .Y(n_1234) );
INVx4_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g1009 ( .A(n_747), .Y(n_1009) );
XNOR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_1029), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_908), .B2(n_1028), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OA22x2_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_825), .B2(n_826), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_770), .B(n_790), .C(n_791), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_783), .C(n_784), .Y(n_770) );
NOR3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .C(n_781), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_773), .B(n_803), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_799), .C(n_823), .Y(n_793) );
INVxp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_806), .B1(n_816), .B2(n_820), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_801), .A2(n_821), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
A2O1A1Ixp33_ASAP7_75t_L g1045 ( .A1(n_801), .A2(n_1019), .B(n_1046), .C(n_1047), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_802), .A2(n_807), .B1(n_808), .B2(n_811), .Y(n_806) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g881 ( .A(n_809), .Y(n_881) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g1510 ( .A(n_810), .Y(n_1510) );
INVx5_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx6_ASAP7_75t_L g903 ( .A(n_815), .Y(n_903) );
BUFx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
BUFx3_ASAP7_75t_L g1570 ( .A(n_821), .Y(n_1570) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_871), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_862), .C(n_870), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_838), .C(n_845), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .B1(n_834), .B2(n_835), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_832), .A2(n_835), .B1(n_1544), .B2(n_1545), .Y(n_1543) );
AND2x4_ASAP7_75t_L g835 ( .A(n_833), .B(n_836), .Y(n_835) );
AND2x4_ASAP7_75t_L g870 ( .A(n_833), .B(n_861), .Y(n_870) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_840), .B1(n_843), .B2(n_844), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_839), .A2(n_843), .B1(n_886), .B2(n_888), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_840), .B(n_1064), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1581 ( .A1(n_840), .A2(n_844), .B1(n_1561), .B2(n_1564), .Y(n_1581) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g1068 ( .A(n_842), .Y(n_1068) );
AOI33xp33_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_848), .A3(n_850), .B1(n_852), .B2(n_856), .B3(n_859), .Y(n_845) );
INVx1_ASAP7_75t_L g1556 ( .A(n_846), .Y(n_1556) );
BUFx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g1522 ( .A(n_847), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_849), .A2(n_939), .B1(n_940), .B2(n_941), .Y(n_938) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx3_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx3_ASAP7_75t_L g1553 ( .A(n_857), .Y(n_1553) );
BUFx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_861), .A2(n_1107), .B1(n_1149), .B2(n_1161), .Y(n_1183) );
INVx8_ASAP7_75t_L g1540 ( .A(n_863), .Y(n_1540) );
AND2x4_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
INVx1_ASAP7_75t_L g947 ( .A(n_865), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_865), .B(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1069 ( .A(n_867), .Y(n_1069) );
INVx3_ASAP7_75t_L g1538 ( .A(n_868), .Y(n_1538) );
INVx3_ASAP7_75t_L g1546 ( .A(n_870), .Y(n_1546) );
INVx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g1566 ( .A1(n_874), .A2(n_884), .B1(n_1539), .B2(n_1567), .C(n_1568), .Y(n_1566) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_875), .Y(n_1013) );
INVx1_ASAP7_75t_L g1165 ( .A(n_875), .Y(n_1165) );
AOI21xp5_ASAP7_75t_SL g876 ( .A1(n_877), .A2(n_883), .B(n_884), .Y(n_876) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
BUFx6f_ASAP7_75t_L g1565 ( .A(n_890), .Y(n_1565) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx4_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx3_ASAP7_75t_L g1572 ( .A(n_895), .Y(n_1572) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
NOR2x1_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g1047 ( .A(n_899), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_902), .B1(n_903), .B2(n_904), .C(n_905), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_903), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx3_ASAP7_75t_L g1056 ( .A(n_907), .Y(n_1056) );
INVx1_ASAP7_75t_L g1577 ( .A(n_907), .Y(n_1577) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_908), .Y(n_1028) );
XNOR2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_969), .Y(n_908) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_967), .B(n_968), .Y(n_909) );
AND3x1_ASAP7_75t_L g910 ( .A(n_911), .B(n_944), .C(n_951), .Y(n_910) );
AOI31xp33_ASAP7_75t_L g968 ( .A1(n_911), .A2(n_944), .A3(n_951), .B(n_967), .Y(n_968) );
NAND3xp33_ASAP7_75t_SL g912 ( .A(n_913), .B(n_924), .C(n_928), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_919), .B2(n_922), .Y(n_913) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_927), .B(n_1170), .Y(n_1169) );
INVxp67_ASAP7_75t_L g981 ( .A(n_929), .Y(n_981) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_931), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_934), .A2(n_1122), .B1(n_1123), .B2(n_1126), .Y(n_1121) );
INVx3_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
BUFx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g1084 ( .A(n_936), .Y(n_1084) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_937), .Y(n_1116) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_949), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx3_ASAP7_75t_L g1020 ( .A(n_964), .Y(n_1020) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_964), .Y(n_1061) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
NAND3xp33_ASAP7_75t_L g971 ( .A(n_972), .B(n_979), .C(n_1003), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
OAI21xp33_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_993), .B(n_1002), .Y(n_979) );
OAI211xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B(n_984), .C(n_987), .Y(n_980) );
OAI211xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B(n_991), .C(n_992), .Y(n_987) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_988), .A2(n_997), .B1(n_1016), .B2(n_1017), .C(n_1018), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NOR3xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1014), .C(n_1023), .Y(n_1003) );
INVxp67_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
XNOR2xp5_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1143), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
XNOR2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1094), .Y(n_1032) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1062), .Y(n_1036) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1043), .B(n_1044), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1048), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_1049), .A2(n_1051), .B1(n_1052), .B2(n_1053), .Y(n_1048) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1049), .Y(n_1579) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_1053), .A2(n_1066), .B1(n_1067), .B2(n_1069), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1057), .B1(n_1058), .B2(n_1060), .Y(n_1054) );
NAND3xp33_ASAP7_75t_SL g1062 ( .A(n_1063), .B(n_1065), .C(n_1070), .Y(n_1062) );
NOR2xp33_ASAP7_75t_SL g1070 ( .A(n_1071), .B(n_1074), .Y(n_1070) );
OAI33xp33_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1077), .A3(n_1081), .B1(n_1086), .B2(n_1090), .B3(n_1093), .Y(n_1074) );
BUFx4f_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1081) );
INVx8_ASAP7_75t_L g1176 ( .A(n_1083), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_1084), .A2(n_1087), .B1(n_1088), .B2(n_1089), .Y(n_1086) );
NAND4xp75_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1131), .C(n_1139), .D(n_1140), .Y(n_1095) );
OAI21xp5_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1100), .B(n_1105), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_1099), .A2(n_1153), .B1(n_1181), .B2(n_1184), .Y(n_1180) );
A2O1A1Ixp33_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .B(n_1108), .C(n_1109), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1117), .B1(n_1121), .B2(n_1127), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1113), .B1(n_1115), .B2(n_1116), .Y(n_1111) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
BUFx4f_ASAP7_75t_SL g1123 ( .A(n_1124), .Y(n_1123) );
INVx3_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1189), .B1(n_1190), .B2(n_1236), .Y(n_1143) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1144), .Y(n_1236) );
OAI21x1_ASAP7_75t_SL g1144 ( .A1(n_1145), .A2(n_1146), .B(n_1188), .Y(n_1144) );
NAND4xp25_ASAP7_75t_L g1188 ( .A(n_1145), .B(n_1148), .C(n_1150), .D(n_1167), .Y(n_1188) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
NAND3xp33_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1150), .C(n_1167), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1155), .Y(n_1150) );
NAND3xp33_ASAP7_75t_SL g1155 ( .A(n_1156), .B(n_1159), .C(n_1162), .Y(n_1155) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
NAND3xp33_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1173), .C(n_1180), .Y(n_1168) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_1174), .A2(n_1175), .B1(n_1177), .B2(n_1178), .Y(n_1173) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
NOR2x1_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1216), .Y(n_1191) );
A2O1A1Ixp33_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1197), .B(n_1213), .C(n_1214), .Y(n_1192) );
NOR3xp33_ASAP7_75t_SL g1197 ( .A(n_1198), .B(n_1206), .C(n_1207), .Y(n_1197) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1224), .Y(n_1216) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
BUFx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1447), .B1(n_1449), .B2(n_1523), .C(n_1527), .Y(n_1237) );
NOR3xp33_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1385), .C(n_1427), .Y(n_1238) );
A2O1A1Ixp33_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1319), .B(n_1337), .C(n_1341), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_1241), .A2(n_1266), .B1(n_1274), .B2(n_1285), .C(n_1292), .Y(n_1240) );
AOI221xp5_ASAP7_75t_SL g1386 ( .A1(n_1241), .A2(n_1325), .B1(n_1387), .B2(n_1389), .C(n_1391), .Y(n_1386) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1257), .Y(n_1242) );
INVx3_ASAP7_75t_L g1318 ( .A(n_1243), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1243), .B(n_1308), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1243), .B(n_1258), .Y(n_1329) );
INVx3_ASAP7_75t_L g1343 ( .A(n_1243), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1243), .B(n_1351), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1243), .B(n_1299), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1243), .B(n_1258), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1243), .B(n_1306), .Y(n_1446) );
AND2x4_ASAP7_75t_SL g1243 ( .A(n_1244), .B(n_1251), .Y(n_1243) );
AND2x6_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1246), .B(n_1250), .Y(n_1249) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_1246), .B(n_1253), .Y(n_1252) );
AND2x6_ASAP7_75t_L g1255 ( .A(n_1246), .B(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1246), .B(n_1250), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1246), .B(n_1250), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1246), .B(n_1253), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1248), .B(n_1254), .Y(n_1253) );
HB1xp67_ASAP7_75t_L g1584 ( .A(n_1253), .Y(n_1584) );
INVx2_ASAP7_75t_SL g1378 ( .A(n_1257), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1262), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1258), .B(n_1287), .Y(n_1286) );
NAND2xp5_ASAP7_75t_SL g1293 ( .A(n_1258), .B(n_1294), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1258), .B(n_1263), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1258), .B(n_1318), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1258), .B(n_1263), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1258), .B(n_1338), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1261), .Y(n_1258) );
AND2x4_ASAP7_75t_L g1347 ( .A(n_1259), .B(n_1261), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1262), .B(n_1347), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1395 ( .A(n_1262), .B(n_1314), .Y(n_1395) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1262), .B(n_1289), .Y(n_1419) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1263), .Y(n_1299) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1263), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1265), .Y(n_1263) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1266), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1266), .B(n_1336), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1266), .B(n_1302), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1266), .B(n_1354), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1271), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1267), .B(n_1284), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1267), .B(n_1271), .Y(n_1326) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1267), .Y(n_1368) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1268), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1268), .B(n_1271), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1271), .Y(n_1284) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1271), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1430 ( .A(n_1271), .B(n_1297), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1273), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1281), .Y(n_1274) );
OAI22xp33_ASAP7_75t_L g1444 ( .A1(n_1275), .A2(n_1349), .B1(n_1411), .B2(n_1445), .Y(n_1444) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1280), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1276), .B(n_1283), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1276), .B(n_1335), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1279), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1277), .B(n_1279), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1280), .B(n_1305), .Y(n_1304) );
A2O1A1Ixp33_ASAP7_75t_L g1370 ( .A1(n_1281), .A2(n_1371), .B(n_1373), .C(n_1377), .Y(n_1370) );
OAI221xp5_ASAP7_75t_L g1410 ( .A1(n_1281), .A2(n_1411), .B1(n_1412), .B2(n_1413), .C(n_1414), .Y(n_1410) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1282), .B(n_1314), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1283), .B(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1283), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1283), .B(n_1305), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1284), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1287), .B(n_1315), .Y(n_1350) );
AOI32xp33_ASAP7_75t_L g1359 ( .A1(n_1287), .A2(n_1360), .A3(n_1364), .B1(n_1365), .B2(n_1369), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1287), .B(n_1402), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1287), .B(n_1323), .Y(n_1412) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1288), .B(n_1322), .Y(n_1321) );
NAND2xp5_ASAP7_75t_SL g1345 ( .A(n_1288), .B(n_1346), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1288), .B(n_1375), .Y(n_1374) );
NAND2xp5_ASAP7_75t_SL g1436 ( .A(n_1288), .B(n_1325), .Y(n_1436) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1289), .B(n_1299), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1302 ( .A(n_1289), .B(n_1297), .Y(n_1302) );
INVx3_ASAP7_75t_L g1314 ( .A(n_1289), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1289), .B(n_1297), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1289), .B(n_1318), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1291), .Y(n_1289) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1300), .C(n_1307), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1298), .Y(n_1294) );
CKINVDCx14_ASAP7_75t_R g1295 ( .A(n_1296), .Y(n_1295) );
AOI32xp33_ASAP7_75t_L g1377 ( .A1(n_1296), .A2(n_1378), .A3(n_1379), .B1(n_1380), .B2(n_1384), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g1305 ( .A(n_1297), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1297), .B(n_1312), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1297), .B(n_1316), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1297), .B(n_1323), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1297), .B(n_1368), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1297), .B(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1299), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1299), .B(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1299), .Y(n_1382) );
OAI322xp33_ASAP7_75t_L g1391 ( .A1(n_1299), .A2(n_1348), .A3(n_1351), .B1(n_1392), .B2(n_1393), .C1(n_1396), .C2(n_1397), .Y(n_1391) );
O2A1O1Ixp33_ASAP7_75t_L g1420 ( .A1(n_1299), .A2(n_1421), .B(n_1422), .C(n_1425), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_1299), .A2(n_1303), .B1(n_1432), .B2(n_1434), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1299), .B(n_1433), .Y(n_1432) );
OAI21xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1303), .B(n_1306), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1302), .B(n_1325), .Y(n_1384) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1305), .B(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1305), .B(n_1361), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1305), .B(n_1368), .Y(n_1372) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1305), .B(n_1436), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1305), .B(n_1323), .Y(n_1443) );
AOI222xp33_ASAP7_75t_L g1428 ( .A1(n_1306), .A2(n_1322), .B1(n_1346), .B2(n_1354), .C1(n_1378), .C2(n_1429), .Y(n_1428) );
A2O1A1Ixp33_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1310), .B(n_1313), .C(n_1317), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1308), .B(n_1317), .Y(n_1369) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1309), .B(n_1322), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1309), .B(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1312), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1314), .Y(n_1336) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1316), .Y(n_1390) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1317), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1318), .B(n_1375), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1411 ( .A(n_1318), .B(n_1376), .Y(n_1411) );
NOR3xp33_ASAP7_75t_L g1418 ( .A(n_1318), .B(n_1362), .C(n_1419), .Y(n_1418) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1318), .B(n_1440), .Y(n_1439) );
O2A1O1Ixp33_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1324), .B(n_1327), .C(n_1328), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1323), .B(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1323), .Y(n_1363) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1324), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1325), .B(n_1354), .Y(n_1433) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OAI21xp5_ASAP7_75t_L g1328 ( .A1(n_1329), .A2(n_1330), .B(n_1331), .Y(n_1328) );
A2O1A1Ixp33_ASAP7_75t_L g1380 ( .A1(n_1329), .A2(n_1381), .B(n_1382), .C(n_1383), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1333), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1332), .B(n_1336), .Y(n_1417) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1336), .B(n_1367), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1336), .B(n_1430), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1337), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1337), .Y(n_1381) );
AOI221xp5_ASAP7_75t_L g1406 ( .A1(n_1337), .A2(n_1407), .B1(n_1408), .B2(n_1410), .C(n_1420), .Y(n_1406) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
OAI221xp5_ASAP7_75t_L g1385 ( .A1(n_1338), .A2(n_1381), .B1(n_1386), .B2(n_1398), .C(n_1406), .Y(n_1385) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1338), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
AOI211xp5_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1344), .B(n_1355), .C(n_1370), .Y(n_1341) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1343), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1348), .B1(n_1349), .B2(n_1351), .C(n_1352), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1346), .B(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1346), .Y(n_1400) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1347), .Y(n_1351) );
NOR2xp33_ASAP7_75t_L g1408 ( .A(n_1347), .B(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
OAI21xp33_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B(n_1359), .Y(n_1355) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1358), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1363), .Y(n_1361) );
NOR2xp33_ASAP7_75t_L g1394 ( .A(n_1362), .B(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1364), .Y(n_1413) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1379), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1381), .B(n_1396), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1382), .B(n_1404), .Y(n_1403) );
INVxp67_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
AOI31xp33_ASAP7_75t_SL g1414 ( .A1(n_1390), .A2(n_1415), .A3(n_1417), .B(n_1418), .Y(n_1414) );
INVxp67_ASAP7_75t_SL g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1395), .Y(n_1442) );
NOR2xp33_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1403), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1401), .Y(n_1399) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
AOI211xp5_ASAP7_75t_L g1438 ( .A1(n_1405), .A2(n_1426), .B(n_1439), .C(n_1444), .Y(n_1438) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
A2O1A1Ixp33_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1431), .B(n_1437), .C(n_1438), .Y(n_1427) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVxp67_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1443), .Y(n_1441) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
BUFx2_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
HB1xp67_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
NAND4xp75_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1481), .C(n_1506), .D(n_1514), .Y(n_1452) );
AO21x1_ASAP7_75t_L g1453 ( .A1(n_1454), .A2(n_1461), .B(n_1478), .Y(n_1453) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_1455), .A2(n_1456), .B1(n_1458), .B2(n_1459), .Y(n_1454) );
AOI22xp5_ASAP7_75t_L g1482 ( .A1(n_1455), .A2(n_1458), .B1(n_1483), .B2(n_1485), .Y(n_1482) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1475), .Y(n_1461) );
NAND3xp33_ASAP7_75t_L g1462 ( .A(n_1463), .B(n_1469), .C(n_1472), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_1464), .A2(n_1465), .B1(n_1467), .B2(n_1468), .Y(n_1463) );
NAND2xp5_ASAP7_75t_L g1493 ( .A(n_1464), .B(n_1494), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1466), .B(n_1471), .Y(n_1470) );
INVx2_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1474), .Y(n_1472) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
AO21x1_ASAP7_75t_L g1481 ( .A1(n_1482), .A2(n_1487), .B(n_1500), .Y(n_1481) );
INVx2_ASAP7_75t_SL g1483 ( .A(n_1484), .Y(n_1483) );
NOR3xp33_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1496), .C(n_1499), .Y(n_1487) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1492), .Y(n_1490) );
AND2x4_ASAP7_75t_L g1494 ( .A(n_1491), .B(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1504), .Y(n_1501) );
INVx1_ASAP7_75t_SL g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
AOI32xp33_ASAP7_75t_L g1514 ( .A1(n_1515), .A2(n_1516), .A3(n_1518), .B1(n_1520), .B2(n_1521), .Y(n_1514) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
BUFx3_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
BUFx2_ASAP7_75t_SL g1528 ( .A(n_1529), .Y(n_1528) );
BUFx3_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVxp33_ASAP7_75t_SL g1531 ( .A(n_1532), .Y(n_1531) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
NAND2xp67_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1558), .Y(n_1536) );
AOI221xp5_ASAP7_75t_L g1537 ( .A1(n_1538), .A2(n_1539), .B1(n_1540), .B2(n_1541), .C(n_1542), .Y(n_1537) );
NAND3xp33_ASAP7_75t_SL g1542 ( .A(n_1543), .B(n_1546), .C(n_1547), .Y(n_1542) );
AOI222xp33_ASAP7_75t_L g1571 ( .A1(n_1544), .A2(n_1545), .B1(n_1572), .B2(n_1573), .C1(n_1575), .C2(n_1578), .Y(n_1571) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_1548), .A2(n_1551), .B1(n_1555), .B2(n_1557), .Y(n_1547) );
INVx2_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1554), .Y(n_1551) );
BUFx2_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
NAND3xp33_ASAP7_75t_SL g1559 ( .A(n_1560), .B(n_1566), .C(n_1571), .Y(n_1559) );
AOI22xp5_ASAP7_75t_L g1560 ( .A1(n_1561), .A2(n_1562), .B1(n_1564), .B2(n_1565), .Y(n_1560) );
HB1xp67_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
OAI21xp5_ASAP7_75t_L g1582 ( .A1(n_1583), .A2(n_1584), .B(n_1585), .Y(n_1582) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
endmodule