module fake_jpeg_21760_n_143 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_13),
.B1(n_12),
.B2(n_16),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_37),
.B1(n_24),
.B2(n_28),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_16),
.C(n_12),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_27),
.C(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_13),
.B1(n_16),
.B2(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_25),
.B(n_21),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_31),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_19),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_37),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_37),
.B1(n_35),
.B2(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_57),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_64),
.B1(n_35),
.B2(n_39),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_46),
.C(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_36),
.B1(n_23),
.B2(n_27),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_49),
.B1(n_35),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_78),
.B1(n_36),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_26),
.B1(n_36),
.B2(n_24),
.Y(n_78)
);

XOR2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_54),
.Y(n_79)
);

XNOR2x1_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_92),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_57),
.B(n_58),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_85),
.B(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_53),
.B(n_17),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_90),
.B1(n_30),
.B2(n_43),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_27),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_84),
.C(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_102),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_72),
.B(n_11),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_93),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_20),
.B1(n_10),
.B2(n_14),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_91),
.B1(n_89),
.B2(n_84),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_105),
.B(n_90),
.C(n_82),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

AOI211xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_105),
.B(n_23),
.C(n_27),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_98),
.CI(n_104),
.CON(n_119),
.SN(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_100),
.C(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_119),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_109),
.B1(n_107),
.B2(n_30),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_30),
.C(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_109),
.C(n_20),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_128),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_18),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_0),
.C(n_2),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_5),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_119),
.A3(n_122),
.B1(n_120),
.B2(n_121),
.C1(n_5),
.C2(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_7),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_4),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_137),
.C(n_9),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_136),
.B1(n_8),
.B2(n_9),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_127),
.C(n_131),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_138),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_7),
.B(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_7),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_140),
.Y(n_143)
);


endmodule