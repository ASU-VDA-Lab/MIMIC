module fake_jpeg_2789_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_41),
.B(n_58),
.C(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_54),
.B1(n_62),
.B2(n_46),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_46),
.B1(n_57),
.B2(n_54),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_72),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_40),
.B1(n_51),
.B2(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_65),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_73),
.C(n_75),
.Y(n_95)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_88),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_58),
.B1(n_43),
.B2(n_45),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_1),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_55),
.B1(n_53),
.B2(n_52),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_68),
.B1(n_47),
.B2(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_3),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_100),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_8),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_47),
.B(n_6),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_81),
.B(n_86),
.Y(n_115)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_92),
.B1(n_87),
.B2(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_5),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_7),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_92),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_127),
.B(n_14),
.Y(n_136)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_87),
.B1(n_90),
.B2(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_121),
.B1(n_128),
.B2(n_96),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_22),
.B1(n_38),
.B2(n_36),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_97),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_9),
.B(n_10),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_13),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_134),
.B1(n_117),
.B2(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_101),
.B1(n_106),
.B2(n_13),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_29),
.C(n_17),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_143),
.C(n_121),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_30),
.B(n_18),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_39),
.B(n_27),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_20),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_138),
.C(n_143),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_149),
.B(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_139),
.C(n_141),
.Y(n_155)
);

OAI321xp33_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_132),
.A3(n_133),
.B1(n_142),
.B2(n_116),
.C(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_151),
.C(n_112),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_154),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_116),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_116),
.B(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_33),
.C(n_34),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_14),
.Y(n_162)
);


endmodule