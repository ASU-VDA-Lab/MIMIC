module fake_jpeg_5473_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_31),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_31),
.Y(n_57)
);

XNOR2x1_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_27),
.B1(n_18),
.B2(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_34),
.B1(n_31),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_21),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_28),
.B1(n_30),
.B2(n_22),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_34),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_74),
.B(n_26),
.Y(n_105)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_80),
.B1(n_83),
.B2(n_67),
.Y(n_106)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_59),
.B1(n_51),
.B2(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_84),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_51),
.B1(n_50),
.B2(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_17),
.Y(n_93)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx12f_ASAP7_75t_SL g95 ( 
.A(n_68),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_110),
.C(n_29),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_98),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_51),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_119),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_68),
.B1(n_81),
.B2(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_106),
.B1(n_88),
.B2(n_73),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_67),
.B1(n_52),
.B2(n_55),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_114),
.B(n_72),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_25),
.B(n_23),
.C(n_32),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_67),
.B1(n_46),
.B2(n_25),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_25),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_102),
.C(n_105),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_70),
.B(n_90),
.C(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_46),
.B1(n_23),
.B2(n_32),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_65),
.B(n_24),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_121),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_78),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_126),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_123),
.A2(n_143),
.B(n_19),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_33),
.B1(n_75),
.B2(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_77),
.B1(n_69),
.B2(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_141),
.B1(n_142),
.B2(n_149),
.Y(n_164)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_144),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_65),
.B1(n_77),
.B2(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_29),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_82),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_77),
.B1(n_28),
.B2(n_30),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_106),
.B1(n_104),
.B2(n_107),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_166),
.B1(n_176),
.B2(n_131),
.Y(n_181)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_156),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_172),
.Y(n_185)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_168),
.Y(n_188)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_58),
.B1(n_121),
.B2(n_24),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_167),
.B(n_132),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_58),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_177),
.C(n_127),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_118),
.B1(n_99),
.B2(n_21),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_137),
.B(n_139),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_98),
.B(n_33),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_133),
.B(n_134),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_33),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_126),
.B1(n_124),
.B2(n_122),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_33),
.B1(n_75),
.B2(n_8),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_75),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_129),
.B(n_7),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_8),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_184),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

XOR2x1_ASAP7_75t_SL g218 ( 
.A(n_194),
.B(n_161),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_132),
.B1(n_140),
.B2(n_143),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_204),
.B1(n_206),
.B2(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_179),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_132),
.B(n_148),
.C(n_146),
.D(n_147),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_180),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_163),
.C(n_159),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_203),
.B(n_205),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_164),
.B1(n_155),
.B2(n_168),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_151),
.A2(n_132),
.B1(n_125),
.B2(n_2),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_211),
.C(n_228),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_190),
.C(n_185),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_157),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_223),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_227),
.B1(n_216),
.B2(n_221),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_132),
.B1(n_168),
.B2(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_156),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_181),
.A2(n_171),
.B1(n_169),
.B2(n_158),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_7),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_226),
.Y(n_234)
);

XNOR2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_0),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_186),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_230),
.A2(n_214),
.B(n_209),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_191),
.B(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_241),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_183),
.C(n_189),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_182),
.B1(n_184),
.B2(n_2),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_226),
.B1(n_224),
.B2(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_184),
.C(n_1),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_184),
.C(n_1),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_0),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_1),
.C(n_2),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_208),
.C(n_225),
.Y(n_259)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_215),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_255),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_219),
.Y(n_255)
);

OAI211xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_227),
.B(n_244),
.C(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_260),
.B(n_245),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_262),
.B(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_3),
.C(n_4),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_248),
.B1(n_234),
.B2(n_231),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

BUFx4f_ASAP7_75t_SL g265 ( 
.A(n_261),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_282)
);

XNOR2x2_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_241),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_271),
.B(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_239),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_231),
.Y(n_271)
);

XNOR2x2_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_248),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_239),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_278),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_274),
.B1(n_238),
.B2(n_270),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_269),
.B1(n_10),
.B2(n_6),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_246),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_237),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_236),
.C(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_262),
.B1(n_254),
.B2(n_259),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_283),
.B1(n_11),
.B2(n_15),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_9),
.B1(n_12),
.B2(n_6),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_284),
.A3(n_10),
.B1(n_6),
.B2(n_7),
.C1(n_11),
.C2(n_15),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_15),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_289),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_293),
.B(n_285),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_294),
.B(n_298),
.Y(n_301)
);


endmodule