module fake_jpeg_26568_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_0),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_21),
.Y(n_32)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_13),
.C(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_20),
.A2(n_9),
.B1(n_12),
.B2(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_18),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_27),
.B(n_29),
.C(n_33),
.Y(n_53)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_42),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.C(n_39),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_30),
.B(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_45),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_22),
.B(n_27),
.C(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_27),
.B1(n_36),
.B2(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_20),
.C(n_3),
.Y(n_62)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_63),
.B1(n_14),
.B2(n_3),
.C(n_4),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

AOI221xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.C(n_22),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_31),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_18),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_86),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_40),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_81),
.B(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

OAI322xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_72),
.A3(n_18),
.B1(n_23),
.B2(n_6),
.C1(n_7),
.C2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_89),
.B(n_5),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_81),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_90),
.B(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_33),
.B1(n_36),
.B2(n_28),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_94),
.A3(n_33),
.B1(n_6),
.B2(n_1),
.C1(n_5),
.C2(n_24),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_28),
.B(n_31),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_99),
.B(n_1),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.B1(n_104),
.B2(n_28),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_23),
.Y(n_108)
);


endmodule