module fake_aes_2824_n_1364 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1364);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1364;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1275;
wire n_955;
wire n_1093;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx2_ASAP7_75t_L g288 ( .A(n_222), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_163), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_195), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_265), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_131), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_116), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_143), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_84), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_2), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_49), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_186), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_52), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_286), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_248), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_144), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_78), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_170), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_5), .Y(n_306) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_214), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_43), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_225), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_14), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_118), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_21), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_112), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_249), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_63), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_145), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_194), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_169), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_201), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_208), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_279), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_287), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_27), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_34), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_93), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_105), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_11), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_187), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_247), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_9), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_179), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_182), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_207), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_146), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_228), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_53), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_285), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_238), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_141), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_156), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_229), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_74), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_220), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_203), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_50), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_172), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_43), .Y(n_349) );
INVxp33_ASAP7_75t_SL g350 ( .A(n_13), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_269), .Y(n_351) );
INVxp33_ASAP7_75t_SL g352 ( .A(n_40), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_108), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_164), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_2), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_155), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_134), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_234), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_242), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_284), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_151), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_136), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_109), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_273), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_76), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_88), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_99), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_123), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_69), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_137), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_154), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_9), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_274), .B(n_24), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_276), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_254), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_266), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_259), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_264), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_79), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_36), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_49), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_86), .B(n_73), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_261), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_184), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_221), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_165), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_215), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_87), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_90), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_233), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_271), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_260), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_161), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_39), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_96), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_244), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_56), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_245), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_81), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_177), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_29), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_8), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_51), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_54), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_227), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_91), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_189), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_217), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_98), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_16), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_55), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_106), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_198), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_56), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_66), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_27), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_219), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_152), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_183), .Y(n_419) );
BUFx2_ASAP7_75t_SL g420 ( .A(n_175), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_119), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_48), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_199), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_262), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_255), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_14), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_212), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_19), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_13), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_125), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_293), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_312), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_293), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_312), .Y(n_434) );
INVx6_ASAP7_75t_L g435 ( .A(n_300), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_347), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_307), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_380), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_293), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_337), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_324), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_380), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_381), .Y(n_443) );
BUFx8_ASAP7_75t_L g444 ( .A(n_373), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_381), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_293), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_345), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_349), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_345), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_345), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_345), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_347), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_359), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_386), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_359), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_410), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_359), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_359), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_288), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_289), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_295), .B(n_0), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_365), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_297), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_436), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_454), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_461), .B(n_360), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
AO22x2_ASAP7_75t_L g469 ( .A1(n_461), .A2(n_401), .B1(n_429), .B2(n_338), .Y(n_469) );
INVx4_ASAP7_75t_L g470 ( .A(n_435), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_441), .B(n_375), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_439), .Y(n_472) );
AND2x6_ASAP7_75t_L g473 ( .A(n_436), .B(n_373), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_436), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_460), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_460), .Y(n_476) );
NOR2x1p5_ASAP7_75t_L g477 ( .A(n_437), .B(n_306), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
NAND2xp33_ASAP7_75t_L g479 ( .A(n_440), .B(n_292), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
AND2x6_ASAP7_75t_L g481 ( .A(n_462), .B(n_300), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_460), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_460), .B(n_382), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_452), .B(n_306), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_448), .B(n_394), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_454), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_452), .B(n_456), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
AND2x6_ASAP7_75t_L g491 ( .A(n_456), .B(n_305), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_457), .B(n_355), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_431), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_439), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_457), .B(n_355), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_435), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_446), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_432), .B(n_368), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_432), .B(n_411), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_434), .A2(n_352), .B1(n_350), .B2(n_317), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_434), .B(n_296), .Y(n_504) );
AND2x6_ASAP7_75t_L g505 ( .A(n_444), .B(n_305), .Y(n_505) );
AND2x6_ASAP7_75t_L g506 ( .A(n_444), .B(n_314), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_438), .B(n_411), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_438), .B(n_379), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_444), .B(n_292), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_489), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_502), .B(n_309), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_489), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_468), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_502), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_507), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_507), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_473), .A2(n_469), .B1(n_506), .B2(n_505), .Y(n_518) );
XNOR2xp5_ASAP7_75t_L g519 ( .A(n_488), .B(n_464), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_467), .B(n_444), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_473), .B(n_311), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_487), .B(n_316), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_473), .B(n_311), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_465), .A2(n_474), .B(n_468), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_510), .B(n_385), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_487), .A2(n_352), .B1(n_350), .B2(n_309), .Y(n_526) );
INVx5_ASAP7_75t_L g527 ( .A(n_473), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_504), .B(n_299), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_471), .B(n_406), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_483), .B(n_336), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_482), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_471), .A2(n_317), .B1(n_396), .B2(n_384), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_483), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_482), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_484), .B(n_336), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_473), .A2(n_435), .B1(n_325), .B2(n_328), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_483), .B(n_340), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_469), .A2(n_396), .B1(n_425), .B2(n_384), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_473), .B(n_340), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_482), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_475), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_473), .A2(n_425), .B1(n_464), .B2(n_416), .Y(n_543) );
AO22x1_ASAP7_75t_L g544 ( .A1(n_503), .A2(n_351), .B1(n_357), .B2(n_348), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_468), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_475), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_473), .B(n_348), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_492), .B(n_351), .Y(n_548) );
AND3x2_ASAP7_75t_SL g549 ( .A(n_466), .B(n_308), .C(n_297), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_468), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_476), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_491), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_495), .B(n_357), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_497), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_481), .B(n_371), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_481), .B(n_371), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_504), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_469), .A2(n_332), .B1(n_372), .B2(n_310), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_479), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_477), .B(n_442), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_476), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_504), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_469), .A2(n_477), .B1(n_506), .B2(n_505), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_504), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_465), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_474), .Y(n_568) );
NOR2xp33_ASAP7_75t_R g569 ( .A(n_466), .B(n_308), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_469), .Y(n_570) );
INVx5_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
AND2x6_ASAP7_75t_L g572 ( .A(n_505), .B(n_314), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_481), .B(n_376), .Y(n_573) );
BUFx3_ASAP7_75t_L g574 ( .A(n_481), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_500), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_505), .A2(n_402), .B1(n_403), .B2(n_397), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_491), .Y(n_577) );
INVx5_ASAP7_75t_L g578 ( .A(n_505), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_481), .B(n_376), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_509), .B(n_377), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_470), .A2(n_301), .B(n_288), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_481), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_481), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_505), .B(n_442), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_470), .B(n_387), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_491), .A2(n_291), .B(n_290), .Y(n_586) );
BUFx3_ASAP7_75t_L g587 ( .A(n_481), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_470), .B(n_387), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_505), .B(n_391), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_506), .B(n_391), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_491), .Y(n_591) );
NAND3xp33_ASAP7_75t_SL g592 ( .A(n_486), .B(n_399), .C(n_398), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_506), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_506), .B(n_398), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_491), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_493), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_506), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_575), .A2(n_414), .B(n_415), .C(n_404), .Y(n_598) );
AND2x4_ASAP7_75t_SL g599 ( .A(n_512), .B(n_422), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_569), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_563), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_558), .A2(n_428), .B1(n_426), .B2(n_443), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_565), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_520), .B(n_506), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_528), .Y(n_605) );
CKINVDCx16_ASAP7_75t_R g606 ( .A(n_512), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_528), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_520), .B(n_506), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_524), .A2(n_321), .B(n_294), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_566), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_566), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_516), .B(n_491), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_568), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_571), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_533), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_527), .B(n_399), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_570), .A2(n_491), .B1(n_363), .B2(n_435), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_527), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_527), .B(n_443), .Y(n_619) );
BUFx4_ASAP7_75t_SL g620 ( .A(n_515), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_522), .B(n_445), .Y(n_621) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_532), .Y(n_622) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_518), .A2(n_302), .B(n_298), .Y(n_623) );
NAND2x1_ASAP7_75t_L g624 ( .A(n_572), .B(n_491), .Y(n_624) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_557), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_517), .A2(n_445), .B(n_303), .C(n_313), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_545), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_539), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_564), .A2(n_304), .B(n_318), .C(n_315), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_571), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_571), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_527), .B(n_405), .Y(n_632) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_545), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_548), .B(n_405), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_542), .A2(n_551), .B(n_546), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_526), .B(n_412), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_511), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_514), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_539), .A2(n_319), .B(n_322), .C(n_320), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_513), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_548), .A2(n_499), .B(n_486), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_594), .A2(n_501), .B(n_499), .Y(n_644) );
INVx2_ASAP7_75t_SL g645 ( .A(n_561), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_543), .B(n_412), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_544), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_578), .Y(n_648) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_561), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_576), .A2(n_435), .B1(n_327), .B2(n_330), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_529), .A2(n_329), .B(n_333), .C(n_331), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_536), .B(n_417), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_552), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_537), .A2(n_334), .B1(n_341), .B2(n_339), .Y(n_654) );
NOR2xp67_ASAP7_75t_SL g655 ( .A(n_578), .B(n_417), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_578), .B(n_323), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_560), .B(n_326), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_521), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_552), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_553), .B(n_530), .Y(n_660) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_578), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_531), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_592), .A2(n_420), .B1(n_346), .B2(n_354), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_538), .A2(n_342), .B(n_358), .C(n_356), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_519), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_593), .A2(n_362), .B1(n_364), .B2(n_361), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_580), .B(n_389), .Y(n_667) );
AO22x1_ASAP7_75t_L g668 ( .A1(n_549), .A2(n_369), .B1(n_370), .B2(n_366), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_534), .Y(n_669) );
BUFx3_ASAP7_75t_L g670 ( .A(n_535), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_541), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_581), .A2(n_383), .B(n_388), .C(n_378), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_521), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_523), .A2(n_392), .B(n_393), .C(n_390), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_523), .B(n_1), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_584), .B(n_395), .Y(n_676) );
BUFx8_ASAP7_75t_L g677 ( .A(n_549), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_550), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_540), .Y(n_679) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_552), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_554), .Y(n_681) );
BUFx10_ASAP7_75t_L g682 ( .A(n_525), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_586), .A2(n_409), .B1(n_413), .B2(n_407), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_540), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_547), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_547), .A2(n_421), .B1(n_423), .B2(n_419), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_559), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_567), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_585), .B(n_424), .Y(n_689) );
INVx3_ASAP7_75t_L g690 ( .A(n_577), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_577), .A2(n_430), .B1(n_427), .B2(n_343), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_588), .B(n_335), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_555), .B(n_3), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_596), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_583), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_574), .B(n_335), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_582), .B(n_353), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_577), .B(n_301), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_555), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_556), .B(n_353), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_597), .B(n_343), .Y(n_701) );
OR2x6_ASAP7_75t_L g702 ( .A(n_587), .B(n_344), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_556), .B(n_418), .Y(n_703) );
BUFx3_ASAP7_75t_L g704 ( .A(n_573), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_591), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_573), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_594), .A2(n_508), .B(n_400), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_579), .A2(n_400), .B1(n_408), .B2(n_344), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_595), .A2(n_408), .B(n_418), .C(n_451), .Y(n_709) );
AOI221x1_ASAP7_75t_L g710 ( .A1(n_579), .A2(n_365), .B1(n_367), .B2(n_374), .C(n_458), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_590), .Y(n_711) );
OAI21xp33_ASAP7_75t_SL g712 ( .A1(n_589), .A2(n_459), .B(n_458), .Y(n_712) );
NAND2x1p5_ASAP7_75t_L g713 ( .A(n_572), .B(n_365), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_572), .Y(n_714) );
OAI22x1_ASAP7_75t_L g715 ( .A1(n_572), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_561), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_563), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_570), .A2(n_459), .B1(n_458), .B2(n_367), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_524), .A2(n_493), .B(n_480), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_566), .Y(n_720) );
INVx6_ASAP7_75t_L g721 ( .A(n_561), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_512), .B(n_4), .Y(n_722) );
OAI21x1_ASAP7_75t_L g723 ( .A1(n_719), .A2(n_480), .B(n_472), .Y(n_723) );
INVx2_ASAP7_75t_SL g724 ( .A(n_620), .Y(n_724) );
OAI21x1_ASAP7_75t_L g725 ( .A1(n_719), .A2(n_480), .B(n_472), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_707), .A2(n_485), .B(n_472), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_622), .A2(n_365), .B1(n_367), .B2(n_374), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_607), .Y(n_728) );
OAI21x1_ASAP7_75t_L g729 ( .A1(n_713), .A2(n_490), .B(n_485), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_638), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_641), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_605), .Y(n_732) );
NOR2x1_ASAP7_75t_SL g733 ( .A(n_714), .B(n_367), .Y(n_733) );
AO31x2_ASAP7_75t_L g734 ( .A1(n_710), .A2(n_459), .A3(n_494), .B(n_490), .Y(n_734) );
BUFx2_ASAP7_75t_L g735 ( .A(n_615), .Y(n_735) );
OAI21x1_ASAP7_75t_L g736 ( .A1(n_713), .A2(n_490), .B(n_485), .Y(n_736) );
INVx1_ASAP7_75t_SL g737 ( .A(n_721), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_628), .A2(n_374), .B1(n_453), .B2(n_450), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_608), .A2(n_496), .B(n_494), .Y(n_739) );
NAND2x1p5_ASAP7_75t_L g740 ( .A(n_649), .B(n_680), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_649), .Y(n_741) );
INVx5_ASAP7_75t_L g742 ( .A(n_680), .Y(n_742) );
AOI221x1_ASAP7_75t_L g743 ( .A1(n_715), .A2(n_453), .B1(n_446), .B2(n_447), .C(n_449), .Y(n_743) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_677), .A2(n_374), .B1(n_7), .B2(n_8), .Y(n_744) );
OAI21x1_ASAP7_75t_L g745 ( .A1(n_636), .A2(n_496), .B(n_494), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_643), .Y(n_746) );
INVx4_ASAP7_75t_L g747 ( .A(n_619), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_621), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_601), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_603), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_SL g751 ( .A1(n_629), .A2(n_496), .B(n_127), .C(n_85), .Y(n_751) );
O2A1O1Ixp33_ASAP7_75t_L g752 ( .A1(n_598), .A2(n_6), .B(n_7), .C(n_10), .Y(n_752) );
OAI21x1_ASAP7_75t_SL g753 ( .A1(n_636), .A2(n_10), .B(n_11), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g754 ( .A1(n_604), .A2(n_450), .B(n_446), .C(n_463), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_644), .A2(n_447), .B(n_446), .Y(n_755) );
AOI221x1_ASAP7_75t_L g756 ( .A1(n_623), .A2(n_453), .B1(n_447), .B2(n_463), .C(n_455), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_600), .Y(n_757) );
INVx2_ASAP7_75t_SL g758 ( .A(n_721), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_717), .Y(n_759) );
OAI22xp33_ASAP7_75t_SL g760 ( .A1(n_606), .A2(n_12), .B1(n_15), .B2(n_16), .Y(n_760) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_642), .A2(n_449), .B(n_447), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_613), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_722), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_684), .B(n_12), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_699), .B(n_15), .Y(n_765) );
BUFx12f_ASAP7_75t_L g766 ( .A(n_677), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_674), .A2(n_453), .B(n_447), .C(n_463), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_602), .A2(n_453), .B1(n_449), .B2(n_463), .Y(n_768) );
OAI21x1_ASAP7_75t_L g769 ( .A1(n_705), .A2(n_450), .B(n_449), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_637), .B(n_17), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_662), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_624), .A2(n_450), .B(n_449), .Y(n_772) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_668), .A2(n_453), .B1(n_449), .B2(n_463), .C(n_455), .Y(n_773) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_680), .Y(n_774) );
O2A1O1Ixp33_ASAP7_75t_L g775 ( .A1(n_602), .A2(n_17), .B(n_18), .C(n_19), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_716), .Y(n_776) );
OA21x2_ASAP7_75t_L g777 ( .A1(n_709), .A2(n_455), .B(n_450), .Y(n_777) );
NOR2xp67_ASAP7_75t_L g778 ( .A(n_647), .B(n_18), .Y(n_778) );
OAI21x1_ASAP7_75t_L g779 ( .A1(n_619), .A2(n_455), .B(n_450), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_646), .B(n_20), .Y(n_780) );
OAI21x1_ASAP7_75t_L g781 ( .A1(n_656), .A2(n_463), .B(n_455), .Y(n_781) );
OA21x2_ASAP7_75t_L g782 ( .A1(n_700), .A2(n_455), .B(n_433), .Y(n_782) );
BUFx12f_ASAP7_75t_L g783 ( .A(n_645), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_694), .Y(n_784) );
NOR2x1_ASAP7_75t_SL g785 ( .A(n_702), .B(n_433), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_703), .A2(n_71), .B(n_70), .Y(n_786) );
AO21x2_ASAP7_75t_L g787 ( .A1(n_623), .A2(n_433), .B(n_478), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_599), .Y(n_788) );
BUFx12f_ASAP7_75t_L g789 ( .A(n_682), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_669), .Y(n_790) );
AOI21x1_ASAP7_75t_L g791 ( .A1(n_692), .A2(n_433), .B(n_478), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_682), .B(n_20), .Y(n_792) );
AO21x2_ASAP7_75t_L g793 ( .A1(n_718), .A2(n_433), .B(n_478), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_671), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_660), .B(n_21), .Y(n_795) );
OA21x2_ASAP7_75t_L g796 ( .A1(n_718), .A2(n_433), .B(n_478), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_687), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_708), .A2(n_75), .B(n_72), .Y(n_798) );
BUFx3_ASAP7_75t_L g799 ( .A(n_665), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_635), .B(n_22), .Y(n_800) );
OA21x2_ASAP7_75t_L g801 ( .A1(n_689), .A2(n_498), .B(n_478), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_666), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_685), .B(n_22), .Y(n_803) );
BUFx3_ASAP7_75t_L g804 ( .A(n_681), .Y(n_804) );
AOI21xp33_ASAP7_75t_L g805 ( .A1(n_626), .A2(n_23), .B(n_24), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_708), .A2(n_80), .B(n_77), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_688), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_676), .Y(n_808) );
OAI21x1_ASAP7_75t_L g809 ( .A1(n_698), .A2(n_83), .B(n_82), .Y(n_809) );
O2A1O1Ixp33_ASAP7_75t_L g810 ( .A1(n_640), .A2(n_23), .B(n_25), .C(n_26), .Y(n_810) );
BUFx8_ASAP7_75t_L g811 ( .A(n_676), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_701), .A2(n_92), .B(n_89), .Y(n_812) );
AO31x2_ASAP7_75t_L g813 ( .A1(n_686), .A2(n_25), .A3(n_26), .B(n_28), .Y(n_813) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_614), .Y(n_814) );
AO31x2_ASAP7_75t_L g815 ( .A1(n_686), .A2(n_28), .A3(n_29), .B(n_30), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_651), .A2(n_498), .B(n_478), .C(n_32), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_678), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_683), .A2(n_498), .B1(n_31), .B2(n_32), .Y(n_818) );
OAI21x1_ASAP7_75t_L g819 ( .A1(n_618), .A2(n_95), .B(n_94), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_666), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_702), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_658), .B(n_30), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_683), .B(n_31), .Y(n_823) );
OAI21x1_ASAP7_75t_L g824 ( .A1(n_618), .A2(n_100), .B(n_97), .Y(n_824) );
OAI221xp5_ASAP7_75t_L g825 ( .A1(n_663), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_825) );
INVx6_ASAP7_75t_L g826 ( .A(n_614), .Y(n_826) );
AO21x2_ASAP7_75t_L g827 ( .A1(n_672), .A2(n_498), .B(n_158), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_712), .A2(n_498), .B(n_159), .Y(n_828) );
AO31x2_ASAP7_75t_L g829 ( .A1(n_691), .A2(n_33), .A3(n_35), .B(n_37), .Y(n_829) );
O2A1O1Ixp33_ASAP7_75t_L g830 ( .A1(n_654), .A2(n_37), .B(n_38), .C(n_39), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_711), .A2(n_498), .B(n_162), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_712), .A2(n_38), .B(n_40), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_675), .Y(n_833) );
INVx2_ASAP7_75t_SL g834 ( .A(n_702), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_673), .A2(n_41), .B1(n_42), .B2(n_44), .Y(n_835) );
INVx3_ASAP7_75t_L g836 ( .A(n_614), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_695), .A2(n_166), .B(n_282), .Y(n_837) );
OA21x2_ASAP7_75t_L g838 ( .A1(n_693), .A2(n_160), .B(n_281), .Y(n_838) );
BUFx3_ASAP7_75t_L g839 ( .A(n_696), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_706), .A2(n_41), .B1(n_42), .B2(n_44), .Y(n_840) );
INVx1_ASAP7_75t_SL g841 ( .A(n_679), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_654), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_627), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_625), .B(n_45), .Y(n_844) );
OR2x2_ASAP7_75t_L g845 ( .A(n_652), .B(n_45), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g846 ( .A(n_610), .B(n_101), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_691), .A2(n_171), .B(n_280), .Y(n_847) );
BUFx2_ASAP7_75t_SL g848 ( .A(n_696), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g849 ( .A(n_611), .B(n_102), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_720), .A2(n_168), .B(n_278), .Y(n_850) );
INVxp67_ASAP7_75t_L g851 ( .A(n_612), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_639), .Y(n_852) );
NOR2xp67_ASAP7_75t_L g853 ( .A(n_667), .B(n_46), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_650), .B(n_46), .Y(n_854) );
NAND3x1_ASAP7_75t_L g855 ( .A(n_650), .B(n_47), .C(n_48), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_634), .Y(n_856) );
BUFx2_ASAP7_75t_R g857 ( .A(n_704), .Y(n_857) );
CKINVDCx12_ASAP7_75t_R g858 ( .A(n_655), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_748), .A2(n_664), .B1(n_657), .B2(n_609), .C(n_617), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_746), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_820), .A2(n_670), .B1(n_697), .B2(n_617), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_820), .A2(n_697), .B1(n_690), .B2(n_653), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_802), .A2(n_616), .B1(n_632), .B2(n_659), .Y(n_863) );
OR2x6_ASAP7_75t_L g864 ( .A(n_724), .B(n_630), .Y(n_864) );
INVx4_ASAP7_75t_L g865 ( .A(n_747), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_780), .A2(n_690), .B1(n_653), .B2(n_659), .C(n_661), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_841), .B(n_47), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_842), .A2(n_661), .B1(n_648), .B2(n_633), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_841), .B(n_50), .Y(n_869) );
OA21x2_ASAP7_75t_L g870 ( .A1(n_743), .A2(n_661), .B(n_648), .Y(n_870) );
OAI21xp33_ASAP7_75t_L g871 ( .A1(n_780), .A2(n_648), .B(n_633), .Y(n_871) );
OR2x6_ASAP7_75t_L g872 ( .A(n_789), .B(n_630), .Y(n_872) );
BUFx2_ASAP7_75t_SL g873 ( .A(n_788), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_854), .A2(n_633), .B1(n_631), .B2(n_630), .Y(n_874) );
OR2x2_ASAP7_75t_L g875 ( .A(n_728), .B(n_51), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_763), .A2(n_631), .B1(n_53), .B2(n_54), .C(n_55), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_739), .A2(n_631), .B(n_180), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_833), .B(n_52), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_732), .B(n_57), .Y(n_879) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_754), .A2(n_57), .B(n_58), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_770), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_794), .Y(n_882) );
AO221x2_ASAP7_75t_L g883 ( .A1(n_832), .A2(n_59), .B1(n_60), .B2(n_61), .C(n_62), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_811), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_854), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_823), .A2(n_64), .B1(n_65), .B2(n_67), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_739), .A2(n_191), .B(n_277), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_730), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_749), .B(n_67), .Y(n_889) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_825), .A2(n_68), .B1(n_103), .B2(n_104), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_735), .B(n_68), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_792), .B(n_107), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_731), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_762), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_808), .B(n_110), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_771), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_750), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_792), .A2(n_111), .B1(n_113), .B2(n_114), .C(n_115), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_811), .A2(n_117), .B1(n_120), .B2(n_121), .Y(n_899) );
INVx5_ASAP7_75t_L g900 ( .A(n_747), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_726), .A2(n_122), .B(n_124), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_790), .Y(n_902) );
AND2x4_ASAP7_75t_L g903 ( .A(n_741), .B(n_126), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_759), .B(n_128), .Y(n_904) );
NOR2xp67_ASAP7_75t_L g905 ( .A(n_766), .B(n_129), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_795), .A2(n_130), .B1(n_132), .B2(n_133), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_761), .A2(n_135), .B(n_138), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_795), .B(n_139), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_784), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_817), .B(n_140), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_818), .A2(n_142), .B1(n_147), .B2(n_148), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_825), .A2(n_149), .B1(n_150), .B2(n_153), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_852), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_800), .B(n_157), .Y(n_914) );
AO21x2_ASAP7_75t_L g915 ( .A1(n_754), .A2(n_167), .B(n_173), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_726), .A2(n_174), .B(n_176), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_844), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_797), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_805), .A2(n_178), .B1(n_181), .B2(n_185), .C(n_188), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_807), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_856), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_755), .A2(n_190), .B(n_192), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_816), .A2(n_193), .B1(n_196), .B2(n_197), .C(n_200), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_818), .A2(n_202), .B1(n_204), .B2(n_205), .Y(n_924) );
AOI21xp5_ASAP7_75t_L g925 ( .A1(n_751), .A2(n_206), .B(n_209), .Y(n_925) );
OAI21x1_ASAP7_75t_L g926 ( .A1(n_723), .A2(n_210), .B(n_211), .Y(n_926) );
A2O1A1Ixp33_ASAP7_75t_L g927 ( .A1(n_810), .A2(n_213), .B(n_216), .C(n_218), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_844), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_764), .Y(n_929) );
OA21x2_ASAP7_75t_L g930 ( .A1(n_756), .A2(n_223), .B(n_226), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_843), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_764), .B(n_230), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_751), .A2(n_231), .B(n_232), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_765), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_828), .A2(n_235), .B(n_236), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_828), .A2(n_237), .B(n_239), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_804), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_765), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_753), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_821), .A2(n_240), .B1(n_241), .B2(n_243), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_822), .A2(n_246), .B1(n_250), .B2(n_251), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_822), .Y(n_942) );
OAI22xp5_ASAP7_75t_SL g943 ( .A1(n_744), .A2(n_252), .B1(n_253), .B2(n_257), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_848), .B(n_258), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_835), .A2(n_263), .B1(n_267), .B2(n_268), .Y(n_945) );
AO31x2_ASAP7_75t_L g946 ( .A1(n_767), .A2(n_816), .A3(n_733), .B(n_803), .Y(n_946) );
AND2x4_ASAP7_75t_L g947 ( .A(n_834), .B(n_270), .Y(n_947) );
OAI31xp33_ASAP7_75t_L g948 ( .A1(n_760), .A2(n_272), .A3(n_283), .B(n_775), .Y(n_948) );
INVx3_ASAP7_75t_L g949 ( .A(n_740), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_782), .A2(n_801), .B(n_787), .Y(n_950) );
AND2x4_ASAP7_75t_L g951 ( .A(n_785), .B(n_839), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_813), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_853), .A2(n_855), .B1(n_783), .B2(n_803), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_845), .A2(n_805), .B1(n_835), .B2(n_757), .Y(n_954) );
AOI22x1_ASAP7_75t_L g955 ( .A1(n_740), .A2(n_832), .B1(n_774), .B2(n_814), .Y(n_955) );
BUFx2_ASAP7_75t_R g956 ( .A(n_799), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_737), .B(n_776), .Y(n_957) );
OAI21xp33_ASAP7_75t_L g958 ( .A1(n_727), .A2(n_768), .B(n_773), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_744), .A2(n_840), .B1(n_778), .B2(n_758), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_810), .A2(n_775), .B1(n_830), .B2(n_752), .C(n_737), .Y(n_960) );
BUFx3_ASAP7_75t_L g961 ( .A(n_826), .Y(n_961) );
AO22x1_ASAP7_75t_L g962 ( .A1(n_742), .A2(n_857), .B1(n_774), .B2(n_836), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_813), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_742), .B(n_836), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_813), .B(n_815), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_851), .B(n_752), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_813), .Y(n_967) );
OAI22xp33_ASAP7_75t_SL g968 ( .A1(n_826), .A2(n_830), .B1(n_857), .B2(n_849), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_801), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_815), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_773), .A2(n_851), .B1(n_742), .B2(n_838), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_768), .A2(n_767), .B1(n_738), .B2(n_846), .C(n_849), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_738), .A2(n_846), .B1(n_838), .B2(n_777), .C(n_796), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_826), .A2(n_787), .B1(n_847), .B2(n_793), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_847), .A2(n_793), .B1(n_827), .B2(n_814), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_815), .B(n_829), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_814), .B(n_742), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_815), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_827), .A2(n_814), .B1(n_777), .B2(n_796), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_829), .A2(n_858), .B1(n_798), .B2(n_806), .C(n_786), .Y(n_980) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_782), .A2(n_812), .B1(n_809), .B2(n_831), .Y(n_981) );
AOI221xp5_ASAP7_75t_L g982 ( .A1(n_829), .A2(n_734), .B1(n_824), .B2(n_819), .C(n_745), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_829), .B(n_779), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_837), .B(n_850), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_888), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_952), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_893), .B(n_734), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_900), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_896), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_969), .Y(n_990) );
OR2x2_ASAP7_75t_L g991 ( .A(n_942), .B(n_734), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_902), .Y(n_992) );
INVx4_ASAP7_75t_L g993 ( .A(n_900), .Y(n_993) );
INVx2_ASAP7_75t_L g994 ( .A(n_907), .Y(n_994) );
AND2x4_ASAP7_75t_L g995 ( .A(n_900), .B(n_729), .Y(n_995) );
OR2x2_ASAP7_75t_L g996 ( .A(n_963), .B(n_734), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_967), .B(n_725), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_865), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_897), .Y(n_999) );
NAND2xp5_ASAP7_75t_SL g1000 ( .A(n_971), .B(n_791), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_860), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_882), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_883), .B(n_831), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_883), .B(n_736), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_970), .Y(n_1005) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_900), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_894), .B(n_781), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_907), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_909), .B(n_772), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_931), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_913), .B(n_769), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_889), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_889), .Y(n_1013) );
AOI211xp5_ASAP7_75t_SL g1014 ( .A1(n_968), .A2(n_943), .B(n_862), .C(n_885), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_878), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_929), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_878), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_918), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_865), .B(n_964), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_978), .Y(n_1020) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_964), .B(n_977), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_937), .Y(n_1022) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_874), .Y(n_1023) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_872), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_920), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_953), .B(n_917), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_954), .B(n_934), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_921), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_938), .B(n_976), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_965), .B(n_862), .Y(n_1030) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_977), .B(n_951), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_928), .B(n_966), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_947), .B(n_983), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_879), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_947), .B(n_903), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_875), .B(n_873), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_926), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_959), .B(n_957), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_870), .Y(n_1039) );
NOR4xp25_ASAP7_75t_SL g1040 ( .A(n_923), .B(n_980), .C(n_960), .D(n_898), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1041 ( .A(n_966), .B(n_861), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_891), .B(n_867), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_869), .B(n_859), .Y(n_1043) );
INVxp67_ASAP7_75t_L g1044 ( .A(n_872), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_870), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_948), .A2(n_890), .B1(n_892), .B2(n_903), .Y(n_1046) );
AND2x4_ASAP7_75t_L g1047 ( .A(n_951), .B(n_949), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_885), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_948), .A2(n_876), .B1(n_912), .B2(n_958), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_880), .B(n_886), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_949), .B(n_939), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_881), .B(n_884), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_880), .B(n_904), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_872), .B(n_864), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_904), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_930), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_930), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_910), .B(n_944), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_874), .B(n_864), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_984), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_864), .B(n_910), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_914), .B(n_946), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_895), .B(n_961), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_914), .B(n_946), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_955), .Y(n_1065) );
BUFx3_ASAP7_75t_L g1066 ( .A(n_866), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_905), .Y(n_1067) );
NOR2xp33_ASAP7_75t_SL g1068 ( .A(n_956), .B(n_924), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_946), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_932), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_908), .B(n_911), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_915), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_932), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_908), .B(n_911), .Y(n_1074) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_962), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_924), .A2(n_945), .B1(n_941), .B2(n_868), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_915), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_941), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_981), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_871), .B(n_974), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_973), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1082 ( .A(n_950), .B(n_975), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_927), .B(n_945), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_982), .B(n_919), .Y(n_1084) );
NOR2x1p5_ASAP7_75t_L g1085 ( .A(n_899), .B(n_940), .Y(n_1085) );
INVx2_ASAP7_75t_SL g1086 ( .A(n_863), .Y(n_1086) );
NAND3xp33_ASAP7_75t_L g1087 ( .A(n_1014), .B(n_906), .C(n_936), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_990), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_990), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_985), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1022), .B(n_979), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_1050), .A2(n_972), .B1(n_935), .B2(n_901), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1029), .B(n_916), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1029), .B(n_887), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1016), .B(n_877), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1096 ( .A1(n_1052), .A2(n_922), .B1(n_925), .B2(n_933), .C(n_1026), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_989), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1016), .B(n_992), .Y(n_1098) );
NAND3xp33_ASAP7_75t_L g1099 ( .A(n_1068), .B(n_1067), .C(n_998), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1100 ( .A(n_1030), .B(n_1041), .Y(n_1100) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_1060), .B(n_986), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_999), .B(n_1010), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1033), .B(n_1030), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1034), .B(n_1042), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1001), .Y(n_1105) );
NAND2xp33_ASAP7_75t_R g1106 ( .A(n_1075), .B(n_1035), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1031), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1002), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1038), .B(n_1041), .Y(n_1109) );
NOR2x1_ASAP7_75t_L g1110 ( .A(n_993), .B(n_1006), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1018), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1033), .B(n_1060), .Y(n_1112) );
NOR3xp33_ASAP7_75t_L g1113 ( .A(n_1036), .B(n_1044), .C(n_1054), .Y(n_1113) );
NAND3xp33_ASAP7_75t_L g1114 ( .A(n_1046), .B(n_1049), .C(n_1027), .Y(n_1114) );
BUFx3_ASAP7_75t_L g1115 ( .A(n_1019), .Y(n_1115) );
INVx1_ASAP7_75t_SL g1116 ( .A(n_1019), .Y(n_1116) );
OAI31xp33_ASAP7_75t_SL g1117 ( .A1(n_1035), .A2(n_1076), .A3(n_1019), .B(n_1050), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1043), .B(n_1015), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_986), .B(n_1005), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1025), .B(n_1028), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1017), .B(n_1013), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1005), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1020), .Y(n_1123) );
NAND2xp5_ASAP7_75t_SL g1124 ( .A(n_995), .B(n_1003), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1020), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1012), .B(n_1048), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1032), .B(n_1086), .Y(n_1127) );
AOI221xp5_ASAP7_75t_L g1128 ( .A1(n_1086), .A2(n_1078), .B1(n_1032), .B2(n_1070), .C(n_1073), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1039), .Y(n_1129) );
INVx2_ASAP7_75t_SL g1130 ( .A(n_988), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1039), .Y(n_1131) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1045), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_988), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1021), .B(n_1031), .Y(n_1134) );
AOI21xp5_ASAP7_75t_SL g1135 ( .A1(n_1071), .A2(n_1074), .B(n_993), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1053), .B(n_991), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_1084), .A2(n_1053), .B1(n_1055), .B2(n_1003), .C(n_1023), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_988), .Y(n_1138) );
INVx4_ASAP7_75t_L g1139 ( .A(n_993), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1031), .B(n_1021), .Y(n_1140) );
INVx4_ASAP7_75t_L g1141 ( .A(n_1006), .Y(n_1141) );
BUFx2_ASAP7_75t_L g1142 ( .A(n_1021), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_991), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_987), .B(n_1064), .Y(n_1144) );
INVx3_ASAP7_75t_L g1145 ( .A(n_995), .Y(n_1145) );
OAI321xp33_ASAP7_75t_L g1146 ( .A1(n_1059), .A2(n_1004), .A3(n_1075), .B1(n_1083), .B2(n_1023), .C(n_1082), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1024), .Y(n_1147) );
NAND2xp33_ASAP7_75t_R g1148 ( .A(n_1071), .B(n_1074), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1024), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1061), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1061), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1047), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1058), .B(n_1047), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1069), .B(n_1004), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_1047), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1045), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1059), .Y(n_1157) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_995), .Y(n_1158) );
NOR2x1_ASAP7_75t_L g1159 ( .A(n_1066), .B(n_1085), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_1051), .Y(n_1160) );
INVx2_ASAP7_75t_L g1161 ( .A(n_996), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_996), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1058), .B(n_1055), .Y(n_1163) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_1051), .Y(n_1164) );
INVx2_ASAP7_75t_L g1165 ( .A(n_997), .Y(n_1165) );
INVx4_ASAP7_75t_L g1166 ( .A(n_1066), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1090), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1136), .B(n_1069), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_1141), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1145), .B(n_1082), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1136), .B(n_1081), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1100), .B(n_1062), .Y(n_1172) );
AND2x4_ASAP7_75t_L g1173 ( .A(n_1145), .B(n_1081), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1163), .B(n_1084), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1103), .B(n_1062), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_1141), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1118), .B(n_1083), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1097), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1100), .B(n_1064), .Y(n_1179) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_1145), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1129), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_1101), .B(n_1079), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1103), .B(n_1079), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1184 ( .A(n_1101), .B(n_1080), .Y(n_1184) );
NAND2xp33_ASAP7_75t_L g1185 ( .A(n_1110), .B(n_1063), .Y(n_1185) );
INVx1_ASAP7_75t_SL g1186 ( .A(n_1116), .Y(n_1186) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_1114), .A2(n_1080), .B1(n_1000), .B2(n_1007), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1123), .Y(n_1188) );
OR2x6_ASAP7_75t_L g1189 ( .A(n_1135), .B(n_1077), .Y(n_1189) );
AND2x4_ASAP7_75t_L g1190 ( .A(n_1101), .B(n_997), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1102), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1105), .B(n_1007), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1112), .B(n_1077), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1112), .B(n_1072), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_1141), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1108), .B(n_1040), .Y(n_1196) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1131), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_1120), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1111), .B(n_1009), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1098), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1144), .B(n_1072), .Y(n_1201) );
NOR4xp25_ASAP7_75t_SL g1202 ( .A(n_1106), .B(n_1000), .C(n_1065), .D(n_1057), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1131), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1121), .B(n_1009), .Y(n_1204) );
BUFx3_ASAP7_75t_L g1205 ( .A(n_1115), .Y(n_1205) );
INVx6_ASAP7_75t_L g1206 ( .A(n_1139), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1161), .B(n_1065), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1161), .B(n_994), .Y(n_1208) );
NAND4xp25_ASAP7_75t_L g1209 ( .A(n_1117), .B(n_1011), .C(n_1008), .D(n_994), .Y(n_1209) );
INVx4_ASAP7_75t_L g1210 ( .A(n_1139), .Y(n_1210) );
HB1xp67_ASAP7_75t_L g1211 ( .A(n_1139), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1119), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1132), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1162), .B(n_1008), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1162), .B(n_1011), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_1130), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1109), .B(n_1056), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1119), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1122), .Y(n_1219) );
INVx1_ASAP7_75t_SL g1220 ( .A(n_1115), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1123), .Y(n_1221) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_1113), .A2(n_1037), .B1(n_1056), .B2(n_1057), .C(n_1159), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1125), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1127), .B(n_1037), .Y(n_1224) );
NOR3xp33_ASAP7_75t_L g1225 ( .A(n_1099), .B(n_1087), .C(n_1096), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1104), .B(n_1150), .Y(n_1226) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_1130), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1088), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1151), .B(n_1128), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1088), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1175), .B(n_1154), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1198), .B(n_1212), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1188), .Y(n_1233) );
INVx1_ASAP7_75t_SL g1234 ( .A(n_1206), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1172), .B(n_1144), .Y(n_1235) );
INVxp67_ASAP7_75t_SL g1236 ( .A(n_1169), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1175), .B(n_1154), .Y(n_1237) );
INVxp67_ASAP7_75t_L g1238 ( .A(n_1176), .Y(n_1238) );
BUFx2_ASAP7_75t_L g1239 ( .A(n_1195), .Y(n_1239) );
CKINVDCx16_ASAP7_75t_R g1240 ( .A(n_1210), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1218), .B(n_1143), .Y(n_1241) );
OAI21x1_ASAP7_75t_L g1242 ( .A1(n_1196), .A2(n_1095), .B(n_1091), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1191), .B(n_1137), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1244 ( .A(n_1170), .B(n_1158), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1188), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1183), .B(n_1157), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1183), .B(n_1165), .Y(n_1247) );
NAND2xp5_ASAP7_75t_SL g1248 ( .A(n_1210), .B(n_1211), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1226), .B(n_1153), .Y(n_1249) );
NOR2x1_ASAP7_75t_L g1250 ( .A(n_1210), .B(n_1166), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1193), .B(n_1165), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1252 ( .A(n_1174), .B(n_1166), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1181), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1177), .B(n_1126), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1193), .B(n_1135), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1194), .B(n_1124), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1167), .B(n_1166), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1172), .B(n_1156), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1181), .Y(n_1259) );
INVx3_ASAP7_75t_L g1260 ( .A(n_1206), .Y(n_1260) );
INVxp67_ASAP7_75t_L g1261 ( .A(n_1216), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1171), .B(n_1107), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1221), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1186), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1179), .B(n_1156), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1171), .B(n_1149), .Y(n_1266) );
OR2x6_ASAP7_75t_L g1267 ( .A(n_1189), .B(n_1124), .Y(n_1267) );
INVx1_ASAP7_75t_SL g1268 ( .A(n_1206), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1221), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1200), .B(n_1147), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1229), .B(n_1142), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1178), .B(n_1094), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1219), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1179), .B(n_1089), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_1225), .A2(n_1094), .B1(n_1134), .B2(n_1152), .Y(n_1275) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1239), .Y(n_1276) );
OAI22xp33_ASAP7_75t_L g1277 ( .A1(n_1240), .A2(n_1148), .B1(n_1106), .B2(n_1206), .Y(n_1277) );
AOI22xp5_ASAP7_75t_L g1278 ( .A1(n_1252), .A2(n_1148), .B1(n_1185), .B2(n_1184), .Y(n_1278) );
AOI22xp33_ASAP7_75t_SL g1279 ( .A1(n_1255), .A2(n_1185), .B1(n_1205), .B2(n_1227), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1273), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1273), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1235), .B(n_1168), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1235), .Y(n_1283) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1239), .Y(n_1284) );
AOI32xp33_ASAP7_75t_L g1285 ( .A1(n_1250), .A2(n_1146), .A3(n_1220), .B1(n_1168), .B2(n_1205), .Y(n_1285) );
AOI21xp5_ASAP7_75t_L g1286 ( .A1(n_1248), .A2(n_1202), .B(n_1189), .Y(n_1286) );
OAI21xp33_ASAP7_75t_L g1287 ( .A1(n_1255), .A2(n_1187), .B(n_1209), .Y(n_1287) );
AOI322xp5_ASAP7_75t_L g1288 ( .A1(n_1243), .A2(n_1223), .A3(n_1184), .B1(n_1194), .B2(n_1170), .C1(n_1190), .C2(n_1217), .Y(n_1288) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_1271), .A2(n_1199), .B1(n_1184), .B2(n_1222), .C(n_1192), .Y(n_1289) );
INVxp67_ASAP7_75t_L g1290 ( .A(n_1236), .Y(n_1290) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1258), .Y(n_1291) );
NAND4xp25_ASAP7_75t_SL g1292 ( .A(n_1234), .B(n_1140), .C(n_1092), .D(n_1204), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1293 ( .A1(n_1267), .A2(n_1155), .B1(n_1189), .B2(n_1227), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g1294 ( .A(n_1238), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1232), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1270), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1246), .B(n_1207), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1246), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1274), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1274), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1301 ( .A(n_1244), .B(n_1170), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1247), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_1275), .A2(n_1173), .B1(n_1190), .B2(n_1180), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_1267), .A2(n_1173), .B1(n_1190), .B2(n_1180), .Y(n_1304) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_1261), .A2(n_1189), .B1(n_1092), .B2(n_1224), .C(n_1138), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1280), .Y(n_1306) );
AOI31xp33_ASAP7_75t_SL g1307 ( .A1(n_1286), .A2(n_1257), .A3(n_1266), .B(n_1262), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1281), .Y(n_1308) );
NAND3xp33_ASAP7_75t_L g1309 ( .A(n_1285), .B(n_1264), .C(n_1269), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1288), .B(n_1237), .Y(n_1310) );
NOR3xp33_ASAP7_75t_L g1311 ( .A(n_1292), .B(n_1242), .C(n_1254), .Y(n_1311) );
OAI22xp33_ASAP7_75t_SL g1312 ( .A1(n_1290), .A2(n_1267), .B1(n_1268), .B2(n_1260), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1294), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1294), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1283), .Y(n_1315) );
AOI22xp5_ASAP7_75t_L g1316 ( .A1(n_1287), .A2(n_1249), .B1(n_1256), .B2(n_1244), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g1317 ( .A(n_1290), .Y(n_1317) );
XNOR2x1_ASAP7_75t_L g1318 ( .A(n_1295), .B(n_1237), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1296), .B(n_1231), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1289), .B(n_1231), .Y(n_1320) );
OAI21xp33_ASAP7_75t_L g1321 ( .A1(n_1278), .A2(n_1256), .B(n_1242), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1301), .B(n_1244), .Y(n_1322) );
NOR2x1_ASAP7_75t_L g1323 ( .A(n_1286), .B(n_1260), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1297), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1282), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1310), .B(n_1298), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1317), .B(n_1313), .Y(n_1327) );
OAI21xp5_ASAP7_75t_L g1328 ( .A1(n_1323), .A2(n_1279), .B(n_1277), .Y(n_1328) );
O2A1O1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1307), .A2(n_1305), .B(n_1293), .C(n_1276), .Y(n_1329) );
INVx2_ASAP7_75t_SL g1330 ( .A(n_1322), .Y(n_1330) );
AOI21xp5_ASAP7_75t_L g1331 ( .A1(n_1312), .A2(n_1293), .B(n_1279), .Y(n_1331) );
OAI21xp5_ASAP7_75t_L g1332 ( .A1(n_1309), .A2(n_1303), .B(n_1284), .Y(n_1332) );
OAI21xp33_ASAP7_75t_SL g1333 ( .A1(n_1318), .A2(n_1304), .B(n_1267), .Y(n_1333) );
A2O1A1Ixp33_ASAP7_75t_L g1334 ( .A1(n_1311), .A2(n_1301), .B(n_1260), .C(n_1302), .Y(n_1334) );
OAI211xp5_ASAP7_75t_SL g1335 ( .A1(n_1321), .A2(n_1316), .B(n_1311), .C(n_1320), .Y(n_1335) );
AOI211x1_ASAP7_75t_SL g1336 ( .A1(n_1319), .A2(n_1241), .B(n_1272), .C(n_1291), .Y(n_1336) );
NOR3x1_ASAP7_75t_L g1337 ( .A(n_1314), .B(n_1300), .C(n_1299), .Y(n_1337) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_1333), .A2(n_1315), .B(n_1318), .Y(n_1338) );
AOI211xp5_ASAP7_75t_L g1339 ( .A1(n_1335), .A2(n_1324), .B(n_1325), .C(n_1308), .Y(n_1339) );
AOI221xp5_ASAP7_75t_L g1340 ( .A1(n_1329), .A2(n_1306), .B1(n_1269), .B2(n_1233), .C(n_1263), .Y(n_1340) );
AOI21xp5_ASAP7_75t_L g1341 ( .A1(n_1331), .A2(n_1265), .B(n_1258), .Y(n_1341) );
AOI21xp33_ASAP7_75t_L g1342 ( .A1(n_1328), .A2(n_1133), .B(n_1233), .Y(n_1342) );
OAI21xp33_ASAP7_75t_SL g1343 ( .A1(n_1331), .A2(n_1265), .B(n_1247), .Y(n_1343) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_1337), .Y(n_1344) );
NOR2xp67_ASAP7_75t_L g1345 ( .A(n_1332), .B(n_1263), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1344), .B(n_1330), .Y(n_1346) );
NAND4xp75_ASAP7_75t_L g1347 ( .A(n_1343), .B(n_1326), .C(n_1327), .D(n_1334), .Y(n_1347) );
NAND2x1p5_ASAP7_75t_L g1348 ( .A(n_1341), .B(n_1164), .Y(n_1348) );
NOR2x1_ASAP7_75t_L g1349 ( .A(n_1345), .B(n_1336), .Y(n_1349) );
AOI21xp5_ASAP7_75t_L g1350 ( .A1(n_1340), .A2(n_1245), .B(n_1164), .Y(n_1350) );
OAI211xp5_ASAP7_75t_L g1351 ( .A1(n_1346), .A2(n_1339), .B(n_1338), .C(n_1342), .Y(n_1351) );
OAI222xp33_ASAP7_75t_R g1352 ( .A1(n_1347), .A2(n_1160), .B1(n_1253), .B2(n_1259), .C1(n_1228), .C2(n_1230), .Y(n_1352) );
NAND4xp25_ASAP7_75t_SL g1353 ( .A(n_1349), .B(n_1093), .C(n_1251), .D(n_1201), .Y(n_1353) );
NOR3xp33_ASAP7_75t_L g1354 ( .A(n_1349), .B(n_1173), .C(n_1259), .Y(n_1354) );
NOR2x1_ASAP7_75t_L g1355 ( .A(n_1351), .B(n_1350), .Y(n_1355) );
NOR2x1_ASAP7_75t_L g1356 ( .A(n_1353), .B(n_1348), .Y(n_1356) );
OAI21xp5_ASAP7_75t_L g1357 ( .A1(n_1354), .A2(n_1207), .B(n_1201), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_1355), .A2(n_1352), .B1(n_1182), .B2(n_1251), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1356), .Y(n_1359) );
OAI22xp5_ASAP7_75t_SL g1360 ( .A1(n_1359), .A2(n_1357), .B1(n_1182), .B2(n_1228), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1358), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_1361), .A2(n_1197), .B1(n_1213), .B2(n_1203), .Y(n_1362) );
XNOR2xp5_ASAP7_75t_L g1363 ( .A(n_1362), .B(n_1360), .Y(n_1363) );
AOI22xp5_ASAP7_75t_L g1364 ( .A1(n_1363), .A2(n_1215), .B1(n_1214), .B2(n_1208), .Y(n_1364) );
endmodule