module real_jpeg_25510_n_26 (n_17, n_8, n_0, n_21, n_2, n_142, n_143, n_10, n_9, n_12, n_152, n_147, n_24, n_146, n_6, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_145, n_144, n_5, n_4, n_150, n_1, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_26);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_142;
input n_143;
input n_10;
input n_9;
input n_12;
input n_152;
input n_147;
input n_24;
input n_146;
input n_6;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_150;
input n_1;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;

output n_26;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_1),
.B(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_2),
.B(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_4),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_4),
.B(n_106),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_5),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_123),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_6),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_7),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_8),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_9),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_47),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_40),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_13),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_110),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_18),
.B(n_95),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_19),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_20),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_21),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_45),
.C(n_120),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_23),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_24),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_136),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B(n_133),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_30),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_32),
.B(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_34),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_34),
.B(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_36),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_36),
.B(n_139),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_37),
.B(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_37),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_132),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_126),
.B(n_131),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_122),
.B(n_125),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_51),
.B(n_119),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_49),
.B(n_121),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_50),
.B(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_114),
.B(n_118),
.Y(n_51)
);

OAI321xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_105),
.A3(n_109),
.B1(n_112),
.B2(n_113),
.C(n_142),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_99),
.B(n_104),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_94),
.B(n_98),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_88),
.B(n_93),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_87),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_80),
.B(n_86),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_76),
.B(n_79),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B(n_75),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_137),
.B(n_140),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_143),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_144),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_145),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_146),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_147),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_148),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_149),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_150),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_151),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_152),
.Y(n_111)
);


endmodule