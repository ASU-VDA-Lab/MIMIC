module fake_netlist_6_2865_n_1263 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1263);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1263;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_1094;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_177;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_23),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_76),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_8),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_63),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_121),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_144),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_151),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_74),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_73),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_22),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_56),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_98),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_80),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_95),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_49),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_46),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_91),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_55),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_88),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_162),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_19),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_21),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_79),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_35),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_145),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_22),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_142),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_84),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_114),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_112),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_37),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_87),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_25),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_40),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_134),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_125),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_28),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_93),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_70),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_17),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_120),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_175),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_94),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g271 ( 
.A(n_77),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_149),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_136),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_65),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_62),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_50),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_148),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_68),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_127),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_81),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_67),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_143),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_168),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_36),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_46),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_150),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_139),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_157),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_71),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_171),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_39),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_207),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_181),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_177),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_209),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_200),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_218),
.B(n_0),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_217),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_241),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_281),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_223),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_231),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_214),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_268),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_274),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_205),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_179),
.B(n_0),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_203),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_203),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_197),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_265),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_205),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_179),
.B(n_1),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_185),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_186),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_199),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_198),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_202),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_201),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_232),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_189),
.B(n_1),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_189),
.B(n_2),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_205),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_237),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_183),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_210),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_240),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_212),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_238),
.B(n_3),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_238),
.B(n_4),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_245),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_252),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_253),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_213),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_258),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_204),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_264),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_215),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_219),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_257),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_221),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_224),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_206),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_283),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_283),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_225),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_178),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_183),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_230),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_234),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_235),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_243),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_248),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_183),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_255),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_208),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_178),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_270),
.B(n_4),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_380),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_310),
.A2(n_176),
.B1(n_275),
.B2(n_293),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_297),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_SL g399 ( 
.A(n_368),
.B(n_235),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_276),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_374),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_300),
.Y(n_408)
);

BUFx8_ASAP7_75t_L g409 ( 
.A(n_305),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_180),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_307),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_282),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_339),
.B(n_290),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

AND2x2_ASAP7_75t_SL g420 ( 
.A(n_387),
.B(n_235),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_300),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_329),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_298),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_291),
.Y(n_428)
);

AND2x2_ASAP7_75t_SL g429 ( 
.A(n_387),
.B(n_235),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_367),
.A2(n_294),
.B(n_292),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_312),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_330),
.B(n_235),
.Y(n_435)
);

BUFx8_ASAP7_75t_L g436 ( 
.A(n_305),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_331),
.B(n_279),
.Y(n_437)
);

AND3x2_ASAP7_75t_L g438 ( 
.A(n_337),
.B(n_254),
.C(n_211),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_312),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_279),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_334),
.B(n_180),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_354),
.B(n_182),
.Y(n_443)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_309),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_341),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_346),
.B(n_347),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_355),
.B(n_211),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_304),
.B(n_279),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_319),
.B(n_279),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_313),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_313),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_369),
.B(n_182),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_314),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_350),
.B(n_377),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_314),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_308),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_315),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_456),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_446),
.B(n_299),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_303),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_388),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_376),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_386),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_361),
.C(n_358),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_311),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_446),
.B(n_386),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_306),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_419),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_271),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_426),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_298),
.Y(n_476)
);

AO22x2_ASAP7_75t_L g477 ( 
.A1(n_412),
.A2(n_336),
.B1(n_383),
.B2(n_319),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_317),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_420),
.B(n_279),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_432),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_420),
.A2(n_308),
.B1(n_357),
.B2(n_318),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_357),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_414),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

NOR2x1p5_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_317),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_401),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_391),
.B(n_345),
.C(n_320),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_400),
.B(n_315),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_446),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_443),
.A2(n_327),
.B1(n_352),
.B2(n_365),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_443),
.B(n_442),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_426),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_L g512 ( 
.A(n_442),
.B(n_320),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_420),
.B(n_345),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_410),
.B(n_333),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_429),
.B(n_349),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_429),
.B(n_349),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_316),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_406),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_410),
.B(n_340),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_429),
.B(n_352),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_429),
.A2(n_385),
.B1(n_372),
.B2(n_343),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_399),
.B(n_356),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_444),
.B(n_316),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_502),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_462),
.B(n_434),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_481),
.B(n_400),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_412),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_481),
.B(n_400),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_434),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_481),
.B(n_416),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_416),
.Y(n_536)
);

NOR2x1p5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_434),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_499),
.B(n_416),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_487),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_486),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_486),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_428),
.Y(n_543)
);

NOR3xp33_ASAP7_75t_L g544 ( 
.A(n_506),
.B(n_454),
.C(n_426),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_511),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_428),
.B1(n_430),
.B2(n_417),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_428),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_507),
.A2(n_445),
.B1(n_447),
.B2(n_434),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_499),
.B(n_435),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_519),
.A2(n_364),
.B1(n_445),
.B2(n_454),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_499),
.B(n_435),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_499),
.B(n_435),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_507),
.B(n_430),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_507),
.A2(n_441),
.B(n_437),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_514),
.B(n_409),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_513),
.B(n_409),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_463),
.B(n_356),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_488),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_524),
.B(n_476),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_492),
.B(n_504),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_480),
.B(n_359),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_467),
.B(n_430),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_467),
.B(n_435),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_484),
.B(n_409),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_491),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_464),
.B(n_359),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_520),
.A2(n_301),
.B1(n_302),
.B2(n_326),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_525),
.A2(n_324),
.B1(n_444),
.B2(n_417),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_512),
.A2(n_444),
.B1(n_417),
.B2(n_447),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_493),
.A2(n_417),
.B(n_441),
.C(n_437),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_493),
.B(n_430),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_458),
.B(n_409),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_470),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_470),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_503),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_521),
.A2(n_444),
.B1(n_417),
.B2(n_448),
.Y(n_583)
);

INVx8_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_521),
.B(n_409),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_494),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_494),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_496),
.B(n_216),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_495),
.B(n_430),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_469),
.A2(n_444),
.B1(n_448),
.B2(n_396),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_522),
.B(n_435),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_458),
.B(n_396),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_459),
.B(n_425),
.C(n_411),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_360),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_522),
.Y(n_596)
);

BUFx5_ASAP7_75t_L g597 ( 
.A(n_495),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_504),
.B(n_448),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_500),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_500),
.B(n_448),
.Y(n_600)
);

AO221x1_ASAP7_75t_L g601 ( 
.A1(n_477),
.A2(n_438),
.B1(n_436),
.B2(n_408),
.C(n_451),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_528),
.B(n_411),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_528),
.B(n_360),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_505),
.B(n_430),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_477),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_517),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_505),
.B(n_448),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_465),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_528),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_465),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_466),
.B(n_437),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_473),
.B(n_363),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_473),
.B(n_363),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_468),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_515),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_471),
.B(n_425),
.C(n_365),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_471),
.B(n_441),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_L g620 ( 
.A(n_472),
.B(n_348),
.C(n_408),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_473),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_472),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_517),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_473),
.B(n_438),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_477),
.A2(n_496),
.B1(n_457),
.B2(n_421),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_479),
.B(n_423),
.Y(n_626)
);

AND2x2_ASAP7_75t_SL g627 ( 
.A(n_556),
.B(n_461),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_575),
.Y(n_628)
);

BUFx4f_ASAP7_75t_L g629 ( 
.A(n_539),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_554),
.A2(n_482),
.B(n_479),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_554),
.A2(n_485),
.B(n_482),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_531),
.A2(n_485),
.B1(n_489),
.B2(n_490),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_562),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_489),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_578),
.B(n_436),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_436),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_587),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_596),
.B(n_421),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_531),
.A2(n_490),
.B(n_474),
.C(n_478),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_530),
.A2(n_449),
.B(n_439),
.C(n_450),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_536),
.B(n_515),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_555),
.A2(n_516),
.B(n_501),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_565),
.B(n_477),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_549),
.A2(n_516),
.B(n_501),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_533),
.A2(n_518),
.B1(n_509),
.B2(n_508),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_564),
.A2(n_509),
.B(n_508),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_551),
.A2(n_516),
.B(n_501),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_553),
.A2(n_518),
.B(n_515),
.Y(n_650)
);

NAND2x1_ASAP7_75t_L g651 ( 
.A(n_617),
.B(n_599),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_542),
.B(n_439),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_564),
.A2(n_523),
.B(n_474),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_608),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_610),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_547),
.B(n_523),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_598),
.A2(n_592),
.B(n_529),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_543),
.B(n_461),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_533),
.A2(n_478),
.B(n_483),
.C(n_451),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_536),
.A2(n_497),
.B(n_483),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_535),
.A2(n_457),
.B(n_450),
.C(n_422),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_611),
.Y(n_663)
);

AND2x4_ASAP7_75t_SL g664 ( 
.A(n_602),
.B(n_211),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_545),
.B(n_318),
.Y(n_665)
);

NAND2x1_ASAP7_75t_L g666 ( 
.A(n_617),
.B(n_390),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_538),
.A2(n_497),
.B(n_406),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_436),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_538),
.A2(n_497),
.B(n_413),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_577),
.A2(n_395),
.B(n_394),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_563),
.B(n_436),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_593),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_625),
.A2(n_422),
.B(n_431),
.C(n_427),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_605),
.B(n_184),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_577),
.A2(n_405),
.B(n_390),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_625),
.A2(n_422),
.B(n_431),
.C(n_427),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_546),
.A2(n_497),
.B(n_413),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_548),
.B(n_184),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_548),
.B(n_187),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_557),
.B(n_453),
.Y(n_680)
);

OAI321xp33_ASAP7_75t_L g681 ( 
.A1(n_568),
.A2(n_397),
.A3(n_403),
.B1(n_392),
.B2(n_393),
.C(n_402),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_600),
.A2(n_497),
.B(n_413),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_602),
.B(n_550),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_562),
.B(n_392),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_566),
.B(n_567),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_590),
.A2(n_418),
.B(n_415),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_613),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_590),
.A2(n_418),
.B(n_415),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_579),
.B(n_453),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_602),
.B(n_393),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_580),
.B(n_581),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_619),
.B(n_453),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_607),
.A2(n_497),
.B(n_413),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_612),
.A2(n_413),
.B(n_407),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_575),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_604),
.A2(n_418),
.B(n_415),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_619),
.B(n_453),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_620),
.B(n_397),
.Y(n_698)
);

AO21x1_ASAP7_75t_L g699 ( 
.A1(n_558),
.A2(n_398),
.B(n_402),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_576),
.A2(n_413),
.B(n_407),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_604),
.A2(n_418),
.B(n_415),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_603),
.B(n_403),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_616),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_534),
.B(n_413),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_572),
.B(n_398),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_622),
.B(n_453),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_597),
.B(n_413),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_597),
.B(n_455),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_584),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_597),
.B(n_455),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_597),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_544),
.B(n_398),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_624),
.A2(n_595),
.B(n_615),
.C(n_614),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_583),
.A2(n_405),
.B(n_390),
.C(n_433),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_626),
.A2(n_433),
.B(n_395),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_584),
.A2(n_433),
.B(n_395),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_621),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_582),
.A2(n_424),
.B(n_422),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_537),
.A2(n_571),
.B1(n_574),
.B2(n_573),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_584),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_585),
.A2(n_427),
.B(n_424),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_597),
.B(n_455),
.Y(n_722)
);

AOI21x1_ASAP7_75t_L g723 ( 
.A1(n_540),
.A2(n_395),
.B(n_394),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_597),
.B(n_453),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_719),
.B(n_591),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_702),
.B(n_609),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_629),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_668),
.B(n_586),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_641),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_628),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_SL g733 ( 
.A(n_713),
.B(n_594),
.C(n_618),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_641),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_634),
.B(n_609),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_709),
.B(n_541),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_678),
.A2(n_609),
.B(n_589),
.C(n_552),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_713),
.B(n_712),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_711),
.B(n_560),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_711),
.A2(n_623),
.B(n_606),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_637),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_678),
.A2(n_569),
.B(n_570),
.C(n_427),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_644),
.B(n_601),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_672),
.B(n_424),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_659),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_695),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_657),
.A2(n_643),
.B(n_704),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_663),
.B(n_424),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_SL g749 ( 
.A1(n_717),
.A2(n_636),
.B1(n_679),
.B2(n_671),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_704),
.A2(n_394),
.B(n_390),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_646),
.A2(n_394),
.B(n_390),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_687),
.B(n_431),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_679),
.A2(n_431),
.B(n_433),
.C(n_405),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_636),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_652),
.B(n_254),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_645),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_703),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_629),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_659),
.B(n_192),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_712),
.B(n_627),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_665),
.B(n_254),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_683),
.A2(n_705),
.B1(n_698),
.B2(n_633),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_654),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_638),
.B(n_398),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_649),
.A2(n_405),
.B(n_423),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_655),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_695),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_692),
.A2(n_405),
.B(n_423),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_633),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_709),
.B(n_54),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_690),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_698),
.A2(n_260),
.B1(n_220),
.B2(n_222),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_638),
.B(n_398),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_684),
.B(n_453),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_697),
.A2(n_423),
.B(n_401),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_627),
.B(n_423),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_635),
.B(n_193),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_656),
.B(n_658),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_684),
.B(n_194),
.Y(n_779)
);

NAND2x1p5_ASAP7_75t_L g780 ( 
.A(n_651),
.B(n_453),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_681),
.B(n_423),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_674),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_685),
.B(n_455),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_648),
.A2(n_194),
.B(n_195),
.C(n_285),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_674),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_691),
.B(n_195),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_640),
.B(n_455),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_720),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_666),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_673),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_664),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_708),
.A2(n_423),
.B(n_401),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_640),
.B(n_455),
.Y(n_793)
);

INVx5_ASAP7_75t_L g794 ( 
.A(n_699),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_630),
.B(n_455),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_741),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_747),
.A2(n_675),
.B(n_670),
.Y(n_797)
);

AO31x2_ASAP7_75t_L g798 ( 
.A1(n_737),
.A2(n_647),
.A3(n_714),
.B(n_632),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_774),
.Y(n_799)
);

OAI22xp33_ASAP7_75t_L g800 ( 
.A1(n_782),
.A2(n_631),
.B1(n_686),
.B2(n_688),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_765),
.A2(n_700),
.B(n_723),
.Y(n_801)
);

INVx5_ASAP7_75t_L g802 ( 
.A(n_774),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_757),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_782),
.B(n_662),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_SL g805 ( 
.A1(n_738),
.A2(n_714),
.B(n_642),
.C(n_680),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_745),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_751),
.A2(n_694),
.B(n_650),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_725),
.A2(n_677),
.B(n_696),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_725),
.A2(n_701),
.B(n_710),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_778),
.A2(n_724),
.B(n_722),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_777),
.A2(n_653),
.B1(n_689),
.B2(n_642),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_734),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_744),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_SL g814 ( 
.A1(n_738),
.A2(n_707),
.B(n_676),
.C(n_706),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_790),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_771),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_755),
.B(n_285),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_729),
.A2(n_707),
.B(n_661),
.Y(n_818)
);

OAI22xp33_ASAP7_75t_L g819 ( 
.A1(n_788),
.A2(n_286),
.B1(n_293),
.B2(n_295),
.Y(n_819)
);

AO32x2_ASAP7_75t_L g820 ( 
.A1(n_749),
.A2(n_660),
.A3(n_639),
.B1(n_716),
.B2(n_715),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_758),
.B(n_286),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_786),
.B(n_667),
.Y(n_822)
);

AO21x2_ASAP7_75t_L g823 ( 
.A1(n_760),
.A2(n_669),
.B(n_682),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_739),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_729),
.A2(n_693),
.B(n_718),
.Y(n_825)
);

NAND3x1_ASAP7_75t_L g826 ( 
.A(n_762),
.B(n_721),
.C(n_6),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_730),
.Y(n_827)
);

NOR4xp25_ASAP7_75t_L g828 ( 
.A(n_785),
.B(n_5),
.C(n_9),
.D(n_10),
.Y(n_828)
);

AO21x2_ASAP7_75t_L g829 ( 
.A1(n_760),
.A2(n_423),
.B(n_455),
.Y(n_829)
);

INVx5_ASAP7_75t_L g830 ( 
.A(n_774),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_792),
.A2(n_401),
.B(n_97),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_735),
.A2(n_295),
.B1(n_251),
.B2(n_284),
.Y(n_832)
);

HB1xp67_ASAP7_75t_SL g833 ( 
.A(n_727),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_784),
.A2(n_226),
.B(n_280),
.Y(n_834)
);

BUFx12f_ASAP7_75t_L g835 ( 
.A(n_791),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_771),
.B(n_228),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_786),
.A2(n_250),
.B(n_277),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_763),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_737),
.A2(n_401),
.B(n_273),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_784),
.A2(n_229),
.B(n_263),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_795),
.A2(n_401),
.B(n_262),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_726),
.B(n_233),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_775),
.A2(n_401),
.B(n_78),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_743),
.B(n_242),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_733),
.A2(n_261),
.B(n_259),
.C(n_247),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_731),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_776),
.A2(n_244),
.B(n_246),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_766),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_783),
.A2(n_401),
.B(n_64),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_776),
.A2(n_59),
.B(n_169),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_787),
.A2(n_58),
.B(n_167),
.Y(n_851)
);

AOI221x1_ASAP7_75t_L g852 ( 
.A1(n_754),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_793),
.A2(n_768),
.B(n_750),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_837),
.A2(n_761),
.B1(n_759),
.B2(n_756),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_796),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_827),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_799),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_806),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_827),
.Y(n_860)
);

INVx6_ASAP7_75t_L g861 ( 
.A(n_799),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_799),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_799),
.A2(n_731),
.B1(n_759),
.B2(n_772),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_802),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_SL g865 ( 
.A1(n_850),
.A2(n_817),
.B1(n_834),
.B2(n_840),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_802),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_844),
.A2(n_779),
.B1(n_773),
.B2(n_770),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_816),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_813),
.B(n_770),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_844),
.A2(n_736),
.B1(n_764),
.B2(n_769),
.Y(n_870)
);

INVx6_ASAP7_75t_L g871 ( 
.A(n_802),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_802),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_830),
.A2(n_791),
.B1(n_736),
.B2(n_730),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_830),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_803),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_830),
.A2(n_767),
.B1(n_734),
.B2(n_746),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_835),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_815),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_838),
.Y(n_879)
);

INVx2_ASAP7_75t_R g880 ( 
.A(n_830),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_824),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_838),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_804),
.A2(n_767),
.B1(n_746),
.B2(n_769),
.Y(n_883)
);

CKINVDCx11_ASAP7_75t_R g884 ( 
.A(n_835),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_824),
.B(n_769),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_819),
.A2(n_769),
.B1(n_748),
.B2(n_752),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_851),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_848),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_846),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_842),
.A2(n_819),
.B1(n_833),
.B2(n_826),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_812),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_848),
.Y(n_892)
);

CKINVDCx11_ASAP7_75t_R g893 ( 
.A(n_812),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_822),
.A2(n_781),
.B1(n_794),
.B2(n_728),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_801),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_836),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_823),
.Y(n_897)
);

CKINVDCx6p67_ASAP7_75t_R g898 ( 
.A(n_821),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_852),
.A2(n_732),
.B1(n_728),
.B2(n_794),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_828),
.B(n_753),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_L g901 ( 
.A1(n_845),
.A2(n_781),
.B(n_742),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_832),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_847),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_851),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_829),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_829),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_826),
.A2(n_732),
.B1(n_794),
.B2(n_789),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_845),
.B(n_789),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_839),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_811),
.A2(n_794),
.B1(n_780),
.B2(n_740),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_797),
.Y(n_911)
);

CKINVDCx6p67_ASAP7_75t_R g912 ( 
.A(n_814),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_805),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_831),
.Y(n_914)
);

CKINVDCx6p67_ASAP7_75t_R g915 ( 
.A(n_814),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_897),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_889),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_858),
.Y(n_918)
);

BUFx2_ASAP7_75t_SL g919 ( 
.A(n_866),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_865),
.A2(n_800),
.B1(n_808),
.B2(n_811),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_881),
.B(n_800),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_903),
.A2(n_809),
.B1(n_810),
.B2(n_818),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_858),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_878),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_878),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_913),
.B(n_798),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_911),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_905),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_889),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_905),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_906),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_881),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_895),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_895),
.A2(n_853),
.B(n_807),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_897),
.B(n_798),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_884),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_897),
.B(n_798),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_903),
.A2(n_805),
.B1(n_823),
.B2(n_825),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_892),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_910),
.A2(n_853),
.B(n_843),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_904),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_861),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_904),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_902),
.A2(n_849),
.B1(n_780),
.B2(n_841),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_887),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_890),
.B(n_11),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_892),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_861),
.Y(n_949)
);

AO21x2_ASAP7_75t_L g950 ( 
.A1(n_900),
.A2(n_843),
.B(n_820),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_887),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_900),
.A2(n_820),
.B(n_798),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_887),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_912),
.B(n_820),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_887),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_887),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_947),
.A2(n_854),
.B(n_902),
.C(n_909),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_939),
.B(n_863),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_946),
.Y(n_959)
);

AO21x1_ASAP7_75t_L g960 ( 
.A1(n_947),
.A2(n_899),
.B(n_907),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_936),
.B(n_855),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_938),
.B(n_954),
.Y(n_962)
);

AO32x1_ASAP7_75t_L g963 ( 
.A1(n_920),
.A2(n_875),
.A3(n_874),
.B1(n_873),
.B2(n_882),
.Y(n_963)
);

NOR2x1p5_ASAP7_75t_L g964 ( 
.A(n_943),
.B(n_898),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_918),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_938),
.B(n_912),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_920),
.A2(n_867),
.B1(n_898),
.B2(n_896),
.Y(n_967)
);

AOI221xp5_ASAP7_75t_L g968 ( 
.A1(n_922),
.A2(n_909),
.B1(n_869),
.B2(n_868),
.C(n_883),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_918),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_928),
.Y(n_970)
);

AOI211xp5_ASAP7_75t_L g971 ( 
.A1(n_922),
.A2(n_901),
.B(n_876),
.C(n_908),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_938),
.B(n_954),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_955),
.B(n_866),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_928),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_954),
.B(n_915),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_937),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_937),
.A2(n_896),
.B(n_888),
.C(n_879),
.Y(n_977)
);

OAI211xp5_ASAP7_75t_L g978 ( 
.A1(n_939),
.A2(n_893),
.B(n_870),
.C(n_884),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_952),
.B(n_915),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_952),
.B(n_926),
.Y(n_980)
);

NOR2x1_ASAP7_75t_SL g981 ( 
.A(n_919),
.B(n_866),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_917),
.B(n_885),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_SL g983 ( 
.A1(n_943),
.A2(n_877),
.B1(n_860),
.B2(n_856),
.Y(n_983)
);

AOI221xp5_ASAP7_75t_L g984 ( 
.A1(n_945),
.A2(n_885),
.B1(n_908),
.B2(n_894),
.C(n_886),
.Y(n_984)
);

AO21x2_ASAP7_75t_L g985 ( 
.A1(n_941),
.A2(n_908),
.B(n_914),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_936),
.B(n_914),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_917),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_945),
.A2(n_877),
.B1(n_856),
.B2(n_860),
.Y(n_988)
);

AOI221xp5_ASAP7_75t_L g989 ( 
.A1(n_921),
.A2(n_862),
.B1(n_872),
.B2(n_891),
.C(n_857),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_941),
.A2(n_872),
.B(n_862),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_941),
.A2(n_866),
.B(n_862),
.C(n_872),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_952),
.B(n_880),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_929),
.B(n_859),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_952),
.B(n_857),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_943),
.B(n_949),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_929),
.B(n_859),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_959),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_987),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_980),
.B(n_944),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_980),
.B(n_944),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_970),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_958),
.B(n_943),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_970),
.Y(n_1003)
);

AOI222xp33_ASAP7_75t_SL g1004 ( 
.A1(n_967),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_17),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_962),
.B(n_944),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_962),
.B(n_972),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_974),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_974),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_965),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_972),
.B(n_944),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_961),
.B(n_936),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_965),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_994),
.B(n_942),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_959),
.B(n_946),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_969),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_959),
.B(n_946),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_973),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_969),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_961),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_994),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_982),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_992),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_992),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1008),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1008),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_SL g1026 ( 
.A1(n_1002),
.A2(n_957),
.B(n_981),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1022),
.B(n_986),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_SL g1028 ( 
.A(n_1004),
.B(n_960),
.C(n_988),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1006),
.B(n_979),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_1017),
.B(n_981),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1022),
.B(n_986),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_1023),
.B(n_985),
.Y(n_1032)
);

NAND3xp33_ASAP7_75t_L g1033 ( 
.A(n_1004),
.B(n_968),
.C(n_971),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_997),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1002),
.A2(n_960),
.B1(n_984),
.B2(n_1017),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_998),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_998),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1021),
.B(n_996),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1006),
.B(n_979),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_997),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_1023),
.B(n_985),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1006),
.B(n_1020),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_SL g1043 ( 
.A1(n_1017),
.A2(n_978),
.B1(n_983),
.B2(n_976),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1020),
.B(n_985),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1013),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_999),
.B(n_966),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1043),
.B(n_976),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1030),
.B(n_1017),
.Y(n_1048)
);

NOR4xp25_ASAP7_75t_SL g1049 ( 
.A(n_1036),
.B(n_977),
.C(n_991),
.D(n_989),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1042),
.B(n_997),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1024),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1024),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1025),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1038),
.B(n_1021),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1025),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1027),
.B(n_1019),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1027),
.B(n_1019),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1037),
.B(n_999),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_1029),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1048),
.B(n_1030),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1056),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1056),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_1047),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_1054),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1059),
.B(n_1035),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1048),
.B(n_1030),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_1044),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1063),
.B(n_1049),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1064),
.B(n_1029),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1065),
.B(n_1039),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_1060),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1060),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1068),
.A2(n_1028),
.B1(n_1033),
.B2(n_1066),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_1071),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1069),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1072),
.B(n_1062),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1070),
.A2(n_1033),
.B1(n_1026),
.B2(n_1048),
.Y(n_1077)
);

OAI333xp33_ASAP7_75t_L g1078 ( 
.A1(n_1068),
.A2(n_1062),
.A3(n_1061),
.B1(n_1026),
.B2(n_1058),
.B3(n_1066),
.C1(n_1053),
.C2(n_1051),
.C3(n_993),
.Y(n_1078)
);

NOR4xp25_ASAP7_75t_L g1079 ( 
.A(n_1068),
.B(n_1067),
.C(n_1044),
.D(n_16),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1071),
.B(n_1057),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1068),
.A2(n_1030),
.B(n_1067),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1069),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_1068),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1071),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1079),
.B(n_1050),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1074),
.B(n_1050),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_1084),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_1083),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1076),
.Y(n_1089)
);

AOI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1079),
.A2(n_1032),
.B(n_1041),
.C(n_990),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_L g1091 ( 
.A(n_1077),
.B(n_964),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_1080),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1075),
.Y(n_1093)
);

AOI221x1_ASAP7_75t_SL g1094 ( 
.A1(n_1078),
.A2(n_1053),
.B1(n_1051),
.B2(n_1052),
.C(n_1055),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1081),
.B(n_1039),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1082),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1073),
.Y(n_1097)
);

OAI221xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1079),
.A2(n_1032),
.B1(n_1041),
.B2(n_1031),
.C(n_1040),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1076),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1078),
.A2(n_1045),
.B1(n_1034),
.B2(n_1040),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1074),
.Y(n_1101)
);

AOI222xp33_ASAP7_75t_L g1102 ( 
.A1(n_1088),
.A2(n_893),
.B1(n_1042),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1094),
.A2(n_1055),
.B1(n_1052),
.B2(n_1034),
.C(n_1046),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1087),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1085),
.B(n_1046),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1093),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1097),
.B(n_1031),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1093),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1087),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1087),
.B(n_1034),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1097),
.A2(n_1034),
.B(n_891),
.C(n_18),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1096),
.Y(n_1112)
);

AO21x1_ASAP7_75t_L g1113 ( 
.A1(n_1100),
.A2(n_14),
.B(n_15),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1092),
.A2(n_995),
.B1(n_975),
.B2(n_966),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1096),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1101),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1089),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1089),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1099),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1101),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1116),
.B(n_1086),
.Y(n_1121)
);

NAND3x1_ASAP7_75t_L g1122 ( 
.A(n_1106),
.B(n_1091),
.C(n_1086),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1104),
.B(n_1109),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_1120),
.B(n_1095),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1104),
.B(n_1098),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1117),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1107),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_L g1128 ( 
.A(n_1108),
.B(n_1095),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1111),
.A2(n_1102),
.B(n_1113),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1105),
.B(n_1090),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1102),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_SL g1132 ( 
.A(n_1119),
.B(n_874),
.C(n_25),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1105),
.B(n_999),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1118),
.B(n_859),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1114),
.A2(n_1110),
.B1(n_1112),
.B2(n_1115),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1103),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1104),
.B(n_1000),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1131),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1138)
);

NAND2xp33_ASAP7_75t_SL g1139 ( 
.A(n_1121),
.B(n_857),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1125),
.A2(n_955),
.B1(n_1012),
.B2(n_1003),
.C(n_1001),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1129),
.A2(n_1012),
.B1(n_1001),
.B2(n_1003),
.C(n_1009),
.Y(n_1141)
);

AOI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1135),
.A2(n_1003),
.B1(n_1001),
.B2(n_1009),
.C(n_1007),
.Y(n_1142)
);

OAI221xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1136),
.A2(n_949),
.B1(n_1011),
.B2(n_997),
.C(n_975),
.Y(n_1143)
);

OAI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1124),
.A2(n_1127),
.B1(n_1128),
.B2(n_1123),
.C(n_1130),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1122),
.A2(n_997),
.B1(n_1011),
.B2(n_1007),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1126),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1126),
.A2(n_1132),
.B1(n_1134),
.B2(n_1137),
.C(n_1133),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1125),
.A2(n_24),
.B(n_26),
.Y(n_1148)
);

NAND4xp25_ASAP7_75t_SL g1149 ( 
.A(n_1129),
.B(n_1000),
.C(n_1013),
.D(n_1005),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_1135),
.B(n_28),
.C(n_29),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1121),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1125),
.A2(n_1009),
.B1(n_1013),
.B2(n_950),
.C(n_1000),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1125),
.A2(n_1016),
.B1(n_1014),
.B2(n_973),
.Y(n_1153)
);

AOI211xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1129),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1121),
.B(n_1005),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1125),
.A2(n_1016),
.B1(n_1014),
.B2(n_973),
.Y(n_1156)
);

NAND4xp25_ASAP7_75t_L g1157 ( 
.A(n_1129),
.B(n_949),
.C(n_1011),
.D(n_921),
.Y(n_1157)
);

XOR2x2_ASAP7_75t_L g1158 ( 
.A(n_1122),
.B(n_30),
.Y(n_1158)
);

NAND4xp25_ASAP7_75t_L g1159 ( 
.A(n_1129),
.B(n_949),
.C(n_32),
.D(n_33),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1129),
.A2(n_857),
.B(n_864),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1125),
.A2(n_950),
.B1(n_942),
.B2(n_1014),
.C(n_1016),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_866),
.C(n_32),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1150),
.A2(n_950),
.B1(n_951),
.B2(n_956),
.Y(n_1163)
);

AOI222xp33_ASAP7_75t_L g1164 ( 
.A1(n_1158),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.C1(n_35),
.C2(n_36),
.Y(n_1164)
);

AOI211xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1144),
.A2(n_38),
.B(n_41),
.C(n_42),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1148),
.A2(n_38),
.B(n_41),
.C(n_42),
.Y(n_1166)
);

AOI211xp5_ASAP7_75t_L g1167 ( 
.A1(n_1159),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1146),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.C(n_47),
.Y(n_1168)
);

AOI211xp5_ASAP7_75t_L g1169 ( 
.A1(n_1160),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1169)
);

OAI211xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1147),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1138),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1171)
);

AOI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1151),
.A2(n_1145),
.B(n_1142),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_1141),
.B(n_52),
.C(n_1005),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1143),
.A2(n_1016),
.B1(n_1014),
.B2(n_942),
.C(n_1018),
.Y(n_1174)
);

OAI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1153),
.A2(n_857),
.B1(n_864),
.B2(n_861),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1157),
.A2(n_941),
.B(n_1018),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1155),
.Y(n_1177)
);

OAI211xp5_ASAP7_75t_L g1178 ( 
.A1(n_1139),
.A2(n_864),
.B(n_1010),
.C(n_946),
.Y(n_1178)
);

NOR4xp25_ASAP7_75t_L g1179 ( 
.A(n_1149),
.B(n_1008),
.C(n_1015),
.D(n_923),
.Y(n_1179)
);

XNOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1156),
.B(n_57),
.Y(n_1180)
);

AOI211xp5_ASAP7_75t_L g1181 ( 
.A1(n_1140),
.A2(n_864),
.B(n_1010),
.C(n_1014),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1161),
.A2(n_1016),
.B1(n_1014),
.B2(n_950),
.C(n_956),
.Y(n_1182)
);

AOI211xp5_ASAP7_75t_L g1183 ( 
.A1(n_1152),
.A2(n_864),
.B(n_1010),
.C(n_1016),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1154),
.A2(n_953),
.B(n_956),
.Y(n_1184)
);

OAI211xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1144),
.A2(n_951),
.B(n_956),
.C(n_953),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1162),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1177),
.B(n_1015),
.Y(n_1187)
);

NOR4xp75_ASAP7_75t_L g1188 ( 
.A(n_1173),
.B(n_951),
.C(n_916),
.D(n_926),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_L g1189 ( 
.A(n_1170),
.B(n_951),
.C(n_953),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1164),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1180),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1172),
.B(n_1008),
.Y(n_1192)
);

XNOR2xp5_ASAP7_75t_L g1193 ( 
.A(n_1167),
.B(n_66),
.Y(n_1193)
);

XNOR2xp5_ASAP7_75t_L g1194 ( 
.A(n_1169),
.B(n_72),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1184),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1185),
.A2(n_861),
.B1(n_871),
.B2(n_919),
.Y(n_1196)
);

NOR2x1_ASAP7_75t_SL g1197 ( 
.A(n_1178),
.B(n_919),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1176),
.B(n_1015),
.Y(n_1198)
);

NAND4xp75_ASAP7_75t_L g1199 ( 
.A(n_1168),
.B(n_918),
.C(n_923),
.D(n_1015),
.Y(n_1199)
);

XNOR2xp5_ASAP7_75t_L g1200 ( 
.A(n_1163),
.B(n_75),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1183),
.A2(n_871),
.B1(n_953),
.B2(n_951),
.Y(n_1201)
);

XNOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1165),
.B(n_1171),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1175),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1179),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1181),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_L g1206 ( 
.A(n_1166),
.B(n_83),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1174),
.B(n_950),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1186),
.B(n_1182),
.Y(n_1208)
);

NOR4xp25_ASAP7_75t_L g1209 ( 
.A(n_1190),
.B(n_923),
.C(n_948),
.D(n_940),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1202),
.B(n_948),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1206),
.B(n_1195),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_SL g1213 ( 
.A(n_1192),
.B(n_871),
.C(n_86),
.Y(n_1213)
);

NOR4xp75_ASAP7_75t_L g1214 ( 
.A(n_1199),
.B(n_1201),
.C(n_1200),
.D(n_1207),
.Y(n_1214)
);

NOR2x1_ASAP7_75t_L g1215 ( 
.A(n_1193),
.B(n_85),
.Y(n_1215)
);

OAI31xp33_ASAP7_75t_L g1216 ( 
.A1(n_1204),
.A2(n_963),
.A3(n_951),
.B(n_940),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1205),
.A2(n_926),
.B(n_916),
.Y(n_1217)
);

NAND4xp25_ASAP7_75t_L g1218 ( 
.A(n_1189),
.B(n_916),
.C(n_925),
.D(n_924),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1187),
.B(n_933),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1194),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1188),
.B(n_933),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1187),
.A2(n_916),
.B1(n_924),
.B2(n_925),
.C(n_933),
.Y(n_1222)
);

OAI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1211),
.A2(n_1196),
.B1(n_1197),
.B2(n_1198),
.C(n_916),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1212),
.Y(n_1224)
);

XOR2x2_ASAP7_75t_L g1225 ( 
.A(n_1215),
.B(n_1197),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1219),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1220),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1208),
.A2(n_1198),
.B1(n_916),
.B2(n_928),
.Y(n_1228)
);

XNOR2xp5_ASAP7_75t_L g1229 ( 
.A(n_1214),
.B(n_89),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1221),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1210),
.B(n_925),
.C(n_924),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1213),
.A2(n_930),
.B1(n_932),
.B2(n_931),
.Y(n_1232)
);

AOI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1217),
.A2(n_1209),
.B1(n_1218),
.B2(n_1216),
.Y(n_1233)
);

XOR2xp5_ASAP7_75t_L g1234 ( 
.A(n_1222),
.B(n_92),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1211),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1211),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1211),
.B(n_96),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1224),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1235),
.A2(n_930),
.B1(n_932),
.B2(n_931),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1230),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1229),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1225),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1236),
.A2(n_930),
.B1(n_932),
.B2(n_931),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1227),
.A2(n_934),
.B1(n_927),
.B2(n_935),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1237),
.A2(n_963),
.B1(n_102),
.B2(n_103),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1234),
.A2(n_934),
.B1(n_927),
.B2(n_935),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1226),
.A2(n_1228),
.B1(n_1233),
.B2(n_1232),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1240),
.Y(n_1248)
);

XNOR2xp5_ASAP7_75t_L g1249 ( 
.A(n_1242),
.B(n_1233),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1238),
.B(n_1241),
.Y(n_1250)
);

AOI221x1_ASAP7_75t_L g1251 ( 
.A1(n_1247),
.A2(n_1231),
.B1(n_1243),
.B2(n_1223),
.C(n_1245),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1246),
.A2(n_934),
.B1(n_927),
.B2(n_935),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1239),
.A2(n_963),
.B1(n_104),
.B2(n_106),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1248),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1249),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1250),
.A2(n_1244),
.B(n_963),
.Y(n_1256)
);

OAI22x1_ASAP7_75t_L g1257 ( 
.A1(n_1251),
.A2(n_963),
.B1(n_109),
.B2(n_113),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1254),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1258),
.A2(n_1255),
.B(n_1257),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1259),
.A2(n_1256),
.B(n_1252),
.Y(n_1260)
);

XNOR2xp5_ASAP7_75t_L g1261 ( 
.A(n_1260),
.B(n_1253),
.Y(n_1261)
);

OAI221xp5_ASAP7_75t_R g1262 ( 
.A1(n_1261),
.A2(n_101),
.B1(n_116),
.B2(n_117),
.C(n_122),
.Y(n_1262)
);

AOI211xp5_ASAP7_75t_L g1263 ( 
.A1(n_1262),
.A2(n_124),
.B(n_135),
.C(n_138),
.Y(n_1263)
);


endmodule