module fake_jpeg_16067_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_13),
.B(n_6),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_40),
.B(n_13),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_91),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_36),
.B1(n_23),
.B2(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_72),
.A2(n_74),
.B1(n_85),
.B2(n_88),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_20),
.B1(n_18),
.B2(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_76),
.B1(n_86),
.B2(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_23),
.B1(n_18),
.B2(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_18),
.B1(n_35),
.B2(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_37),
.B1(n_13),
.B2(n_10),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_29),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_14),
.C(n_11),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_19),
.B1(n_29),
.B2(n_21),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_101),
.A2(n_105),
.B1(n_113),
.B2(n_118),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_15),
.B1(n_27),
.B2(n_10),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_21),
.B1(n_26),
.B2(n_37),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_14),
.C(n_16),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_14),
.C(n_41),
.Y(n_148)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_27),
.B1(n_15),
.B2(n_28),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_45),
.Y(n_122)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_46),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_54),
.B1(n_51),
.B2(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_104),
.B1(n_102),
.B2(n_75),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_125),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_126),
.B(n_129),
.Y(n_198)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_45),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_148),
.Y(n_206)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_90),
.B(n_54),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_114),
.C(n_84),
.Y(n_195)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_16),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_69),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_141),
.B(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_16),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_144),
.C(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_81),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.Y(n_184)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_95),
.Y(n_149)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_68),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_68),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_71),
.B(n_39),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_88),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_78),
.B(n_27),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_97),
.A2(n_51),
.B1(n_27),
.B2(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_2),
.Y(n_197)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_102),
.A2(n_4),
.B1(n_9),
.B2(n_5),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_93),
.B1(n_12),
.B2(n_9),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_3),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_118),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_111),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_176),
.A2(n_208),
.B1(n_199),
.B2(n_209),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_110),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_204),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_123),
.A2(n_104),
.B1(n_113),
.B2(n_83),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_186),
.B1(n_191),
.B2(n_192),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_184),
.A2(n_203),
.B(n_212),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_108),
.B1(n_82),
.B2(n_116),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_106),
.B1(n_117),
.B2(n_93),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_131),
.A2(n_114),
.B1(n_84),
.B2(n_4),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_194),
.A2(n_200),
.B1(n_201),
.B2(n_205),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_194),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_151),
.B1(n_148),
.B2(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_151),
.A2(n_111),
.B1(n_119),
.B2(n_2),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_132),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_0),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_140),
.A2(n_1),
.B1(n_2),
.B2(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_135),
.B1(n_128),
.B2(n_137),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_147),
.A2(n_1),
.B1(n_2),
.B2(n_163),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_153),
.A2(n_1),
.B1(n_2),
.B2(n_166),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_124),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_125),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_150),
.B1(n_146),
.B2(n_139),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_130),
.C(n_124),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_221),
.B(n_240),
.C(n_258),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_184),
.A2(n_150),
.B1(n_146),
.B2(n_139),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_144),
.B1(n_157),
.B2(n_121),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_157),
.B1(n_133),
.B2(n_120),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_126),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_229),
.A2(n_235),
.B(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_120),
.B1(n_127),
.B2(n_161),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_203),
.B1(n_174),
.B2(n_191),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_182),
.B(n_203),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_233),
.B(n_246),
.Y(n_271)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_203),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_183),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_243),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_203),
.B1(n_193),
.B2(n_185),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_237),
.A2(n_248),
.B1(n_250),
.B2(n_226),
.Y(n_290)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_244),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_193),
.A2(n_210),
.B1(n_218),
.B2(n_219),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_242),
.A2(n_257),
.B1(n_254),
.B2(n_236),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_188),
.B(n_216),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_232),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_173),
.B(n_198),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_181),
.A2(n_197),
.B1(n_186),
.B2(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_185),
.A2(n_179),
.B1(n_187),
.B2(n_181),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_211),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_259),
.B(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_205),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_179),
.B(n_187),
.C(n_172),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_172),
.A2(n_175),
.B(n_189),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_196),
.B(n_189),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_238),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_175),
.B(n_217),
.C(n_214),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_235),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_178),
.B1(n_217),
.B2(n_227),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_272),
.A2(n_283),
.B1(n_287),
.B2(n_288),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_274),
.B(n_281),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_282),
.B(n_286),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_295),
.C(n_274),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_281),
.B(n_264),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_230),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_251),
.A2(n_235),
.B(n_233),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_259),
.B(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_237),
.A2(n_230),
.B(n_250),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_228),
.A2(n_248),
.B1(n_225),
.B2(n_245),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_225),
.A2(n_221),
.B1(n_240),
.B2(n_231),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_222),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_294),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_258),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_224),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_224),
.A2(n_238),
.B1(n_243),
.B2(n_239),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_247),
.B1(n_286),
.B2(n_267),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_298),
.A2(n_301),
.B(n_311),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_286),
.B1(n_270),
.B2(n_287),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_308),
.B1(n_318),
.B2(n_269),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_309),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_275),
.A2(n_291),
.B1(n_290),
.B2(n_265),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_282),
.A2(n_271),
.B(n_264),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_322),
.C(n_295),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_313),
.B(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_323),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_265),
.A2(n_288),
.B1(n_269),
.B2(n_268),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_276),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_272),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_331),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_278),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_280),
.C(n_279),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_289),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_333),
.B(n_336),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_273),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_335),
.A2(n_337),
.B(n_344),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_311),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_317),
.A2(n_271),
.B(n_273),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_297),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_263),
.C(n_318),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_296),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

AOI211xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_263),
.B(n_315),
.C(n_323),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_343),
.A2(n_296),
.B1(n_299),
.B2(n_320),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_339),
.C(n_341),
.Y(n_367)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_348),
.A2(n_349),
.B1(n_356),
.B2(n_357),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_307),
.B1(n_320),
.B2(n_319),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_342),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_351),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_332),
.B(n_306),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_361),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_354),
.A2(n_330),
.B(n_337),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_345),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_334),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_344),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_335),
.A2(n_306),
.B1(n_307),
.B2(n_343),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_367),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_336),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_355),
.C(n_363),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_366),
.A2(n_354),
.B(n_359),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_353),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_370),
.C(n_371),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_348),
.A2(n_331),
.B1(n_329),
.B2(n_332),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_349),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_330),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_327),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_376),
.A2(n_372),
.B(n_363),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_366),
.A2(n_373),
.B1(n_347),
.B2(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_375),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_365),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_385),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_384),
.A2(n_378),
.B1(n_367),
.B2(n_380),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_370),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_389),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_328),
.C(n_351),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_390),
.A2(n_382),
.B(n_362),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_357),
.C(n_381),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_350),
.B(n_338),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_368),
.C(n_371),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_325),
.Y(n_395)
);


endmodule