module fake_jpeg_20_n_212 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_212);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_1),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_4),
.Y(n_94)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_68),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_94),
.B(n_51),
.Y(n_99)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_95),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_74),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_81),
.B1(n_60),
.B2(n_54),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_104),
.B1(n_117),
.B2(n_71),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_60),
.B1(n_66),
.B2(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_66),
.B1(n_69),
.B2(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_69),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_56),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_52),
.B(n_70),
.C(n_62),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_75),
.B1(n_5),
.B2(n_6),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_141),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_55),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_57),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_58),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_59),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_140),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_61),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_65),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_63),
.B1(n_75),
.B2(n_6),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_63),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_145),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_152),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_75),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_153),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_157),
.B1(n_13),
.B2(n_14),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_119),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_25),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_7),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_158),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_120),
.B(n_134),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_10),
.B(n_12),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_29),
.C(n_45),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_9),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_145),
.B1(n_153),
.B2(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_167),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_192),
.C(n_171),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_148),
.A3(n_142),
.B1(n_144),
.B2(n_162),
.C1(n_147),
.C2(n_15),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_17),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_196),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_171),
.Y(n_197)
);

OAI322xp33_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_198),
.A3(n_199),
.B1(n_183),
.B2(n_172),
.C1(n_170),
.C2(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_177),
.C(n_174),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_181),
.CI(n_21),
.CON(n_205),
.SN(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_205),
.A2(n_201),
.B1(n_22),
.B2(n_23),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_204),
.B1(n_205),
.B2(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_200),
.C(n_24),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_18),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_49),
.Y(n_210)
);

AOI321xp33_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_31),
.A3(n_32),
.B1(n_33),
.B2(n_37),
.C(n_38),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_44),
.Y(n_212)
);


endmodule