module fake_jpeg_13139_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g214 ( 
.A(n_58),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_65),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_64),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_19),
.B(n_0),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_68),
.B(n_92),
.Y(n_203)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_81),
.Y(n_138)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_20),
.B(n_0),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_84),
.Y(n_127)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_88),
.Y(n_153)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_1),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_33),
.B(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_95),
.B(n_44),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_101),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_18),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_102),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_36),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_104),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_34),
.B(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_114),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_37),
.B(n_18),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_116),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_40),
.B(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_126),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_56),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_41),
.B(n_52),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_40),
.B(n_4),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_56),
.B1(n_28),
.B2(n_32),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_131),
.A2(n_144),
.B1(n_148),
.B2(n_175),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_82),
.B1(n_71),
.B2(n_73),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_94),
.A2(n_56),
.B1(n_48),
.B2(n_32),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_148),
.A2(n_168),
.B(n_175),
.C(n_179),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_60),
.A2(n_48),
.B1(n_32),
.B2(n_51),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_158),
.A2(n_184),
.B1(n_201),
.B2(n_205),
.Y(n_239)
);

BUFx4f_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_83),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_167),
.B(n_183),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_58),
.A2(n_32),
.B1(n_48),
.B2(n_42),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_47),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_188),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_69),
.A2(n_48),
.B1(n_42),
.B2(n_23),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_54),
.C(n_41),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_182),
.B(n_140),
.C(n_127),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_77),
.B(n_43),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_61),
.A2(n_54),
.B1(n_52),
.B2(n_49),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_100),
.A2(n_42),
.B1(n_45),
.B2(n_49),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_186),
.A2(n_187),
.B(n_9),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_111),
.A2(n_42),
.B1(n_45),
.B2(n_50),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_113),
.B(n_51),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_77),
.B(n_53),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_204),
.Y(n_223)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_64),
.Y(n_192)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_72),
.Y(n_198)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_66),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_80),
.B(n_43),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_75),
.A2(n_53),
.B1(n_50),
.B2(n_44),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_203),
.C(n_172),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_93),
.A2(n_96),
.B1(n_123),
.B2(n_122),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_208),
.A2(n_106),
.B1(n_97),
.B2(n_84),
.Y(n_250)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_90),
.B(n_6),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_212),
.B(n_8),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_222),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_133),
.B(n_118),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_128),
.B(n_6),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_218),
.B(n_220),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_132),
.B(n_7),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_115),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_150),
.B(n_109),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_152),
.B(n_7),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_224),
.B(n_229),
.Y(n_322)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_124),
.B1(n_121),
.B2(n_112),
.Y(n_225)
);

AO22x2_ASAP7_75t_L g323 ( 
.A1(n_225),
.A2(n_164),
.B1(n_196),
.B2(n_206),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_117),
.B1(n_116),
.B2(n_154),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_226),
.A2(n_267),
.B1(n_159),
.B2(n_135),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_R g228 ( 
.A(n_157),
.B(n_83),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_228),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_8),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_145),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_231),
.B(n_237),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_129),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_8),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_236),
.B(n_275),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_162),
.Y(n_237)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_110),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_240),
.B(n_242),
.C(n_259),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_155),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_130),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_243),
.Y(n_336)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_245),
.B(n_253),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_249),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_250),
.A2(n_213),
.B1(n_276),
.B2(n_261),
.Y(n_329)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_260),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_254),
.A2(n_274),
.B(n_250),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_153),
.B(n_10),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_255),
.B(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_10),
.Y(n_257)
);

INVx11_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_143),
.B(n_11),
.Y(n_259)
);

INVx2_ASAP7_75t_R g260 ( 
.A(n_214),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_142),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_262),
.B(n_263),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_134),
.Y(n_264)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_209),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_147),
.B(n_12),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_271),
.B(n_272),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_160),
.B(n_17),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_156),
.B(n_12),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_184),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_274),
.A2(n_276),
.B(n_254),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_177),
.B(n_13),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_194),
.A2(n_13),
.B1(n_15),
.B2(n_200),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_163),
.B(n_181),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_281),
.Y(n_344)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_170),
.Y(n_278)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_187),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_279),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_139),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_280),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_141),
.B(n_15),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_161),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_179),
.B1(n_165),
.B2(n_202),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_174),
.B(n_176),
.Y(n_284)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_135),
.Y(n_285)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_154),
.B(n_127),
.CI(n_166),
.CON(n_286),
.SN(n_286)
);

OAI32xp33_ASAP7_75t_L g342 ( 
.A1(n_286),
.A2(n_258),
.A3(n_219),
.B1(n_260),
.B2(n_235),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_210),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_149),
.B(n_210),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_242),
.B(n_252),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_294),
.B(n_306),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_307),
.A2(n_317),
.B1(n_325),
.B2(n_327),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_261),
.A2(n_200),
.B1(n_194),
.B2(n_136),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_308),
.A2(n_313),
.B(n_240),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_222),
.A2(n_186),
.B(n_170),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_218),
.B(n_169),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_256),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_169),
.B1(n_149),
.B2(n_159),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_323),
.Y(n_375)
);

AO21x2_ASAP7_75t_L g383 ( 
.A1(n_323),
.A2(n_332),
.B(n_302),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_239),
.A2(n_225),
.B1(n_261),
.B2(n_288),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_225),
.A2(n_164),
.B1(n_196),
.B2(n_206),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_329),
.A2(n_338),
.B1(n_251),
.B2(n_268),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_240),
.B(n_259),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_225),
.A2(n_213),
.B1(n_261),
.B2(n_272),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_340),
.B1(n_307),
.B2(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_216),
.A2(n_228),
.B1(n_281),
.B2(n_236),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_272),
.A2(n_259),
.B1(n_220),
.B2(n_224),
.Y(n_340)
);

NOR4xp25_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_286),
.C(n_229),
.D(n_275),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_309),
.Y(n_345)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_266),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_347),
.B(n_354),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_348),
.A2(n_357),
.B(n_358),
.Y(n_394)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_359),
.B1(n_362),
.B2(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_356),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_223),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_249),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_325),
.A2(n_264),
.B1(n_238),
.B2(n_270),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_316),
.B(n_241),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g398 ( 
.A1(n_360),
.A2(n_384),
.B(n_386),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_331),
.A2(n_286),
.B(n_278),
.C(n_231),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_372),
.B(n_379),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_333),
.A2(n_285),
.B1(n_247),
.B2(n_232),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_329),
.A2(n_245),
.B(n_282),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_364),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_234),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_335),
.A2(n_233),
.B1(n_243),
.B2(n_265),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_366),
.B(n_321),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_323),
.B1(n_304),
.B2(n_344),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_317),
.A2(n_248),
.B1(n_230),
.B2(n_244),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_368),
.A2(n_376),
.B1(n_378),
.B2(n_385),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_311),
.A2(n_294),
.B1(n_338),
.B2(n_313),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_369),
.A2(n_370),
.B1(n_383),
.B2(n_343),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_294),
.A2(n_227),
.B1(n_235),
.B2(n_246),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_373),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_306),
.A2(n_227),
.B(n_246),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_374),
.A2(n_375),
.B1(n_377),
.B2(n_380),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_327),
.A2(n_308),
.B1(n_300),
.B2(n_340),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_312),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_344),
.A2(n_322),
.B1(n_337),
.B2(n_305),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_292),
.A2(n_303),
.B(n_290),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_312),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_309),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_381),
.Y(n_399)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_301),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_382),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_295),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_323),
.A2(n_342),
.B1(n_292),
.B2(n_303),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_301),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_406),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_366),
.C(n_289),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_393),
.C(n_410),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_289),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_355),
.A2(n_289),
.B1(n_334),
.B2(n_323),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_401),
.A2(n_402),
.B1(n_421),
.B2(n_422),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_355),
.A2(n_334),
.B1(n_322),
.B2(n_316),
.Y(n_402)
);

XOR2x2_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_305),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_417),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_375),
.A2(n_310),
.B1(n_318),
.B2(n_334),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_411),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_314),
.C(n_339),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_383),
.B1(n_367),
.B2(n_349),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_383),
.A2(n_332),
.B1(n_298),
.B2(n_328),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_413),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_383),
.A2(n_298),
.B1(n_336),
.B2(n_315),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_326),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_418),
.C(n_420),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_383),
.A2(n_315),
.B1(n_330),
.B2(n_336),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_416),
.B(n_362),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_364),
.B(n_319),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_349),
.B(n_319),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_351),
.A2(n_299),
.B1(n_330),
.B2(n_341),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_299),
.B1(n_341),
.B2(n_376),
.Y(n_422)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_390),
.B(n_379),
.CI(n_348),
.CON(n_426),
.SN(n_426)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_426),
.B(n_402),
.CI(n_420),
.CON(n_460),
.SN(n_460)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_428),
.A2(n_396),
.B1(n_422),
.B2(n_421),
.Y(n_464)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_357),
.B(n_361),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_430),
.A2(n_436),
.B(n_445),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_389),
.B(n_384),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_446),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_370),
.B1(n_363),
.B2(n_359),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_432),
.A2(n_434),
.B1(n_365),
.B2(n_386),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_358),
.C(n_352),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_418),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_400),
.A2(n_363),
.B1(n_372),
.B2(n_353),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_391),
.A2(n_394),
.B(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_439),
.Y(n_466)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_397),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_441),
.Y(n_468)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_393),
.B(n_373),
.C(n_374),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_417),
.C(n_408),
.Y(n_454)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_443),
.B(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

AO32x1_ASAP7_75t_L g445 ( 
.A1(n_391),
.A2(n_345),
.A3(n_381),
.B1(n_368),
.B2(n_377),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_397),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_395),
.B(n_380),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_447),
.B(n_412),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_406),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_403),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_452),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_398),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_371),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_453),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_456),
.C(n_457),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_409),
.B1(n_411),
.B2(n_388),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_455),
.A2(n_477),
.B1(n_435),
.B2(n_425),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_417),
.C(n_408),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_394),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_415),
.C(n_418),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_459),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_465),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_400),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_462),
.B(n_474),
.Y(n_493)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_464),
.Y(n_484)
);

XOR2x2_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_420),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_430),
.A2(n_396),
.B(n_419),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_416),
.B1(n_419),
.B2(n_399),
.Y(n_471)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_473),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_399),
.C(n_392),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_448),
.A2(n_413),
.B1(n_392),
.B2(n_407),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_450),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_346),
.C(n_350),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_479),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_426),
.B(n_382),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_431),
.A2(n_435),
.B1(n_446),
.B2(n_440),
.Y(n_480)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_468),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_489),
.B(n_492),
.Y(n_515)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_468),
.Y(n_490)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_490),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_461),
.A2(n_425),
.B1(n_428),
.B2(n_450),
.Y(n_491)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_491),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_466),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_496),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_453),
.Y(n_497)
);

OAI211xp5_ASAP7_75t_L g505 ( 
.A1(n_497),
.A2(n_436),
.B(n_437),
.C(n_445),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_503),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_447),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_500),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_439),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_501),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_470),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_504),
.Y(n_509)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_505),
.B(n_507),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_462),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_474),
.Y(n_531)
);

OAI322xp33_ASAP7_75t_L g507 ( 
.A1(n_482),
.A2(n_426),
.A3(n_457),
.B1(n_460),
.B2(n_456),
.C1(n_454),
.C2(n_479),
.Y(n_507)
);

BUFx12_ASAP7_75t_L g508 ( 
.A(n_501),
.Y(n_508)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_494),
.A2(n_469),
.B(n_476),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_510),
.A2(n_521),
.B(n_488),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_455),
.B1(n_484),
.B2(n_477),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_512),
.A2(n_486),
.B1(n_438),
.B2(n_473),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_458),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_487),
.C(n_483),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_494),
.A2(n_476),
.B(n_445),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_519),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_510),
.A2(n_521),
.B(n_516),
.Y(n_523)
);

AOI211xp5_ASAP7_75t_L g544 ( 
.A1(n_523),
.A2(n_535),
.B(n_514),
.C(n_519),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_515),
.B(n_490),
.Y(n_524)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_526),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_493),
.C(n_487),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_520),
.A2(n_484),
.B1(n_498),
.B2(n_504),
.Y(n_529)
);

OAI321xp33_ASAP7_75t_L g547 ( 
.A1(n_529),
.A2(n_534),
.A3(n_517),
.B1(n_508),
.B2(n_514),
.C(n_459),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_509),
.A2(n_503),
.B(n_500),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_511),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_533),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_483),
.C(n_495),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_478),
.C(n_433),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_520),
.A2(n_486),
.B1(n_460),
.B2(n_438),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_518),
.A2(n_432),
.B1(n_475),
.B2(n_433),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_537),
.B(n_540),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_527),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_511),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_518),
.C(n_512),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_452),
.C(n_465),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_543),
.A2(n_535),
.B(n_449),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_544),
.A2(n_547),
.B1(n_508),
.B2(n_522),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_529),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_546),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_527),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_536),
.A2(n_528),
.B1(n_523),
.B2(n_517),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_548),
.B(n_552),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_530),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_550),
.B(n_551),
.Y(n_560)
);

AOI21x1_ASAP7_75t_SL g563 ( 
.A1(n_553),
.A2(n_441),
.B(n_444),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_541),
.A2(n_534),
.B1(n_532),
.B2(n_525),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_555),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_556),
.A2(n_537),
.B(n_538),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_557),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_554),
.A2(n_538),
.B(n_539),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_558),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_552),
.A2(n_543),
.B(n_467),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_563),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_560),
.B(n_561),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_549),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_568),
.B(n_565),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_567),
.A2(n_562),
.B(n_556),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_569),
.B(n_564),
.C(n_555),
.Y(n_571)
);

AOI21x1_ASAP7_75t_L g572 ( 
.A1(n_570),
.A2(n_571),
.B(n_553),
.Y(n_572)
);

AO21x1_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_551),
.B(n_429),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_443),
.Y(n_574)
);


endmodule