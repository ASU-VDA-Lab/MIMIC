module fake_jpeg_13368_n_195 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_7),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_90),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_1),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_83),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_55),
.B1(n_62),
.B2(n_72),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_103),
.B1(n_105),
.B2(n_71),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_78),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_72),
.B1(n_74),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_58),
.B1(n_63),
.B2(n_73),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_100),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_123),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_127),
.Y(n_136)
);

NAND2x1_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_83),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_67),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_76),
.B1(n_60),
.B2(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_57),
.B1(n_81),
.B2(n_80),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_83),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_28),
.C(n_53),
.Y(n_145)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_92),
.B1(n_68),
.B2(n_65),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_71),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_75),
.B1(n_77),
.B2(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_8),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_75),
.B1(n_77),
.B2(n_6),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_138),
.B1(n_42),
.B2(n_45),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_26),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_112),
.B(n_121),
.C(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_31),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_152),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_27),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_47),
.C(n_48),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_10),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_13),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_129),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_171),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_161),
.B(n_135),
.Y(n_174)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_39),
.B(n_51),
.C(n_18),
.D(n_19),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_166),
.B1(n_138),
.B2(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_14),
.B1(n_22),
.B2(n_23),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_30),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_40),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_133),
.B1(n_158),
.B2(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_144),
.B1(n_143),
.B2(n_151),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_147),
.B(n_137),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_161),
.A3(n_165),
.B1(n_160),
.B2(n_145),
.C(n_159),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_183),
.A2(n_184),
.B1(n_179),
.B2(n_182),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_185),
.B(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_186),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_187),
.C(n_181),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_191),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_178),
.B1(n_172),
.B2(n_176),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_165),
.Y(n_195)
);


endmodule