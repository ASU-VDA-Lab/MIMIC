module fake_netlist_1_10451_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_10), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_4), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_4), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_7), .B(n_1), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_2), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_12), .A2(n_8), .B(n_9), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_12), .B(n_0), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_16), .B1(n_13), .B2(n_14), .Y(n_24) );
NOR3xp33_ASAP7_75t_SL g25 ( .A(n_21), .B(n_11), .C(n_14), .Y(n_25) );
AND2x4_ASAP7_75t_SL g26 ( .A(n_25), .B(n_22), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_22), .Y(n_27) );
OAI22xp33_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_21), .B1(n_20), .B2(n_17), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_19), .B1(n_17), .B2(n_3), .C(n_5), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_26), .B1(n_19), .B2(n_3), .Y(n_30) );
OAI22xp33_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_0), .B1(n_1), .B2(n_5), .Y(n_31) );
BUFx6f_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_31), .Y(n_33) );
NAND3xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_19), .C(n_33), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_32), .B1(n_33), .B2(n_30), .Y(n_35) );
endmodule