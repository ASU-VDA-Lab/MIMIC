module real_jpeg_10358_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_1),
.A2(n_26),
.B1(n_30),
.B2(n_38),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_3),
.B(n_63),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_69),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_36),
.B(n_40),
.C(n_125),
.D(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_36),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_78),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_24),
.B(n_140),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_62),
.B(n_74),
.C(n_92),
.D(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_62),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_4),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_157),
.B(n_181),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_58),
.B1(n_66),
.B2(n_80),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_80),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_11),
.A2(n_26),
.B1(n_30),
.B2(n_80),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_12),
.A2(n_54),
.B1(n_58),
.B2(n_66),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_54),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_26),
.B1(n_30),
.B2(n_46),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_15),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_15),
.A2(n_26),
.B1(n_30),
.B2(n_83),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_83),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_116),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_101),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_21),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.CI(n_84),
.CON(n_21),
.SN(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_24),
.A2(n_25),
.B1(n_100),
.B2(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_24),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_24),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_24),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_25),
.A2(n_147),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_25),
.B(n_65),
.Y(n_161)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_26),
.A2(n_43),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_30),
.B(n_41),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_30),
.B(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_47),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_37),
.B1(n_75),
.B2(n_76),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_36),
.A2(n_173),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_37),
.B(n_76),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_39),
.A2(n_47),
.B1(n_137),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_39),
.A2(n_171),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_53),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_47),
.A2(n_51),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_47),
.B(n_65),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.C(n_71),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_50),
.B1(n_71),
.B2(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_64),
.B(n_67),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_59),
.B(n_65),
.C(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_75),
.B(n_77),
.C(n_78),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_75),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_82),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_77),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_81),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.C(n_106),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_102),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_113),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_108),
.A2(n_109),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_112),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_115),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_196),
.B(n_201),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_184),
.B(n_195),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_165),
.B(n_183),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_143),
.B(n_164),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_136),
.C(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_152),
.B(n_163),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_158),
.B(n_162),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_176),
.B2(n_182),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_175),
.C(n_182),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_186),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_192),
.C(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);


endmodule