module fake_jpeg_23559_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_16),
.A2(n_21),
.B1(n_14),
.B2(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_24),
.Y(n_27)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

OR2x2_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_3),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_14),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_31),
.B(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.C(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_23),
.C(n_20),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_18),
.B1(n_15),
.B2(n_22),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_31),
.C(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_26),
.B(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_18),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_45),
.C(n_46),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_49),
.B(n_24),
.Y(n_52)
);


endmodule