module fake_jpeg_21939_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_9),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_14),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_59),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_21),
.B(n_26),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_60),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_32),
.B(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_17),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_23),
.B(n_14),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_22),
.B(n_16),
.Y(n_84)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_2),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_20),
.B(n_27),
.Y(n_69)
);

OAI21x1_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_79),
.B(n_66),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_30),
.A3(n_13),
.B1(n_23),
.B2(n_17),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_60),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_22),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_19),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_57),
.C(n_47),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_69),
.B(n_15),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_87),
.B1(n_72),
.B2(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_83),
.C(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_78),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_100),
.B1(n_96),
.B2(n_82),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_78),
.B1(n_69),
.B2(n_79),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_73),
.C(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_74),
.C(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_81),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_97),
.C(n_84),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_111),
.B1(n_116),
.B2(n_107),
.C(n_4),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_72),
.C(n_96),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_63),
.B1(n_49),
.B2(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_103),
.C(n_108),
.Y(n_122)
);

OAI221xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_82),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_114),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_115),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_127),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_118),
.B(n_112),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_56),
.C(n_64),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_77),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_61),
.B(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_123),
.B(n_9),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

XNOR2x2_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_64),
.Y(n_136)
);


endmodule