module fake_netlist_1_4572_n_809 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_809);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_809;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_58), .Y(n_107) );
OR2x2_ASAP7_75t_L g108 ( .A(n_54), .B(n_103), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_56), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_13), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_74), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_105), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_34), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_44), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_87), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_91), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_63), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_26), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_50), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_48), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_41), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_7), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_88), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_39), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_84), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_16), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_1), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_100), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_27), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_104), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_75), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_65), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_59), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_85), .Y(n_138) );
BUFx10_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_36), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_10), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_46), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_37), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_5), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_79), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_42), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_106), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g148 ( .A(n_97), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_118), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_120), .Y(n_153) );
AOI22xp5_ASAP7_75t_SL g154 ( .A1(n_110), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_154) );
BUFx12f_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_140), .B(n_0), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
BUFx8_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_118), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_141), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
AOI22x1_ASAP7_75t_SL g168 ( .A1(n_110), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_168) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_136), .A2(n_47), .B(n_99), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_158), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_153), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_155), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_155), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_165), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_157), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_149), .B(n_137), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_167), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_160), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_160), .Y(n_186) );
NOR2xp33_ASAP7_75t_R g187 ( .A(n_160), .B(n_109), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_157), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_168), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_168), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_169), .A2(n_114), .B(n_115), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_154), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_162), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_149), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_150), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_150), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_150), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_150), .B(n_148), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_150), .Y(n_203) );
NAND2xp33_ASAP7_75t_R g204 ( .A(n_150), .B(n_144), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g205 ( .A(n_196), .B(n_135), .C(n_143), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_195), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_178), .B(n_139), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_173), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_177), .Y(n_210) );
NOR3xp33_ASAP7_75t_L g211 ( .A(n_193), .B(n_146), .C(n_127), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_176), .Y(n_212) );
INVxp67_ASAP7_75t_SL g213 ( .A(n_184), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_194), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_195), .B(n_111), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_176), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_192), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_183), .B(n_113), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_176), .Y(n_219) );
NAND3xp33_ASAP7_75t_L g220 ( .A(n_188), .B(n_122), .C(n_121), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_181), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_179), .B(n_123), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_202), .B(n_126), .Y(n_223) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_197), .Y(n_224) );
XOR2xp5_ASAP7_75t_L g225 ( .A(n_172), .B(n_109), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_178), .B(n_128), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_202), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_180), .Y(n_228) );
NAND3xp33_ASAP7_75t_L g229 ( .A(n_192), .B(n_119), .C(n_116), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_192), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_180), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_201), .Y(n_232) );
BUFx5_ASAP7_75t_L g233 ( .A(n_198), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g234 ( .A(n_174), .B(n_3), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_170), .B(n_129), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_174), .B(n_107), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_191), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_198), .B(n_132), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_185), .B(n_133), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_200), .B(n_134), .Y(n_240) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_204), .B(n_147), .C(n_138), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_200), .B(n_142), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_199), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_175), .B(n_117), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_185), .B(n_131), .Y(n_246) );
NAND3xp33_ASAP7_75t_L g247 ( .A(n_186), .B(n_131), .C(n_164), .Y(n_247) );
NAND3xp33_ASAP7_75t_L g248 ( .A(n_175), .B(n_166), .C(n_164), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_187), .B(n_151), .Y(n_249) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_189), .A2(n_166), .B1(n_164), .B2(n_161), .C(n_159), .Y(n_250) );
XNOR2xp5_ASAP7_75t_L g251 ( .A(n_182), .B(n_4), .Y(n_251) );
BUFx6f_ASAP7_75t_SL g252 ( .A(n_190), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_203), .B(n_151), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_205), .A2(n_189), .B1(n_203), .B2(n_164), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_221), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_217), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_217), .B(n_151), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_213), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_213), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_227), .B(n_5), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_208), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_206), .B(n_6), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_233), .B(n_159), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_232), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g267 ( .A1(n_236), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_233), .B(n_159), .Y(n_268) );
AND2x6_ASAP7_75t_SL g269 ( .A(n_252), .B(n_8), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_227), .B(n_9), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_205), .B(n_9), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_211), .A2(n_166), .B1(n_164), .B2(n_161), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_210), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_225), .Y(n_276) );
XOR2x2_ASAP7_75t_L g277 ( .A(n_251), .B(n_10), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
NOR3xp33_ASAP7_75t_L g279 ( .A(n_211), .B(n_199), .C(n_12), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_252), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_228), .B(n_11), .Y(n_281) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_245), .B(n_166), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_233), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_233), .Y(n_284) );
AOI22x1_ASAP7_75t_L g285 ( .A1(n_224), .A2(n_166), .B1(n_161), .B2(n_159), .Y(n_285) );
NOR2x1p5_ASAP7_75t_L g286 ( .A(n_235), .B(n_11), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_233), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_224), .A2(n_161), .B(n_159), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_233), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_219), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_231), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_207), .B(n_12), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_229), .A2(n_161), .B(n_55), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_255), .B(n_220), .Y(n_295) );
NOR3xp33_ASAP7_75t_L g296 ( .A(n_273), .B(n_234), .C(n_215), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_276), .B(n_239), .Y(n_297) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_260), .B(n_207), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_259), .A2(n_230), .B1(n_223), .B2(n_250), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_258), .A2(n_230), .B(n_249), .Y(n_300) );
NOR3xp33_ASAP7_75t_SL g301 ( .A(n_280), .B(n_222), .C(n_246), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_256), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_259), .A2(n_250), .B(n_218), .C(n_241), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_286), .B(n_226), .Y(n_304) );
NOR2xp33_ASAP7_75t_R g305 ( .A(n_280), .B(n_243), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_258), .A2(n_240), .B(n_238), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_262), .B(n_13), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_266), .A2(n_248), .B(n_247), .C(n_244), .Y(n_308) );
NAND3xp33_ASAP7_75t_SL g309 ( .A(n_279), .B(n_242), .C(n_237), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_275), .A2(n_14), .B1(n_15), .B2(n_17), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_265), .A2(n_57), .B(n_98), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_277), .B(n_14), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_290), .B(n_15), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_282), .B(n_18), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
AND2x6_ASAP7_75t_L g319 ( .A(n_284), .B(n_19), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_265), .A2(n_20), .B(n_21), .Y(n_320) );
NOR3xp33_ASAP7_75t_SL g321 ( .A(n_263), .B(n_102), .C(n_23), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_310), .B(n_282), .Y(n_322) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_321), .A2(n_294), .B(n_268), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_306), .A2(n_268), .B(n_288), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_303), .A2(n_271), .B(n_261), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_297), .B(n_254), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_313), .Y(n_327) );
BUFx2_ASAP7_75t_R g328 ( .A(n_315), .Y(n_328) );
BUFx2_ASAP7_75t_SL g329 ( .A(n_319), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_311), .B(n_267), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_302), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_319), .Y(n_332) );
BUFx4f_ASAP7_75t_L g333 ( .A(n_319), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_299), .A2(n_272), .B(n_292), .Y(n_334) );
BUFx2_ASAP7_75t_SL g335 ( .A(n_319), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_318), .B(n_287), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_316), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_300), .A2(n_257), .B(n_285), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_314), .A2(n_257), .B(n_289), .Y(n_341) );
INVx6_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_318), .B(n_289), .Y(n_343) );
AOI21x1_ASAP7_75t_L g344 ( .A1(n_317), .A2(n_287), .B(n_281), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_320), .A2(n_289), .B(n_272), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_298), .B(n_295), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_327), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_333), .Y(n_348) );
BUFx10_ASAP7_75t_L g349 ( .A(n_338), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_339), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_328), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_331), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_332), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_333), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_325), .A2(n_308), .B(n_316), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_333), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_329), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
INVx8_ASAP7_75t_L g361 ( .A(n_338), .Y(n_361) );
BUFx2_ASAP7_75t_R g362 ( .A(n_329), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_322), .B(n_312), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_346), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_345), .A2(n_307), .B(n_299), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_335), .A2(n_312), .B1(n_305), .B2(n_277), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_322), .B(n_291), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_333), .Y(n_369) );
AOI21x1_ASAP7_75t_L g370 ( .A1(n_344), .A2(n_283), .B(n_256), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_336), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
BUFx2_ASAP7_75t_SL g373 ( .A(n_332), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_326), .A2(n_296), .B1(n_309), .B2(n_293), .Y(n_374) );
OA21x2_ASAP7_75t_L g375 ( .A1(n_325), .A2(n_274), .B(n_283), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_337), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_301), .B(n_256), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_330), .B(n_264), .Y(n_381) );
BUFx4_ASAP7_75t_SL g382 ( .A(n_342), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_365), .B(n_342), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_367), .A2(n_334), .B1(n_342), .B2(n_338), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_351), .B(n_334), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_363), .A2(n_342), .B1(n_338), .B2(n_343), .Y(n_387) );
NAND2xp33_ASAP7_75t_R g388 ( .A(n_348), .B(n_269), .Y(n_388) );
NOR3xp33_ASAP7_75t_SL g389 ( .A(n_352), .B(n_324), .C(n_342), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_368), .B(n_343), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_347), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_350), .Y(n_392) );
NAND2xp33_ASAP7_75t_R g393 ( .A(n_348), .B(n_337), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_351), .B(n_323), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_363), .A2(n_323), .B1(n_293), .B2(n_264), .Y(n_395) );
NOR2xp33_ASAP7_75t_R g396 ( .A(n_356), .B(n_344), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_374), .A2(n_323), .B1(n_293), .B2(n_264), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_350), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_382), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
BUFx4f_ASAP7_75t_SL g402 ( .A(n_356), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_362), .Y(n_403) );
NOR2xp33_ASAP7_75t_R g404 ( .A(n_356), .B(n_22), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_368), .B(n_343), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_361), .A2(n_323), .B1(n_293), .B2(n_341), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_349), .B(n_24), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_381), .B(n_361), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_381), .B(n_256), .Y(n_410) );
INVxp33_ASAP7_75t_SL g411 ( .A(n_373), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
OR2x6_ASAP7_75t_L g413 ( .A(n_373), .B(n_341), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_361), .Y(n_414) );
NOR2xp33_ASAP7_75t_R g415 ( .A(n_369), .B(n_25), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_361), .A2(n_340), .B1(n_29), .B2(n_30), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_377), .B(n_340), .Y(n_418) );
AND2x4_ASAP7_75t_SL g419 ( .A(n_349), .B(n_28), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_349), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_360), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
OR2x6_ASAP7_75t_L g423 ( .A(n_369), .B(n_31), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_360), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_358), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_360), .B(n_32), .Y(n_426) );
OR2x2_ASAP7_75t_SL g427 ( .A(n_358), .B(n_33), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_364), .B(n_35), .Y(n_428) );
OR2x6_ASAP7_75t_L g429 ( .A(n_358), .B(n_38), .Y(n_429) );
XNOR2xp5_ASAP7_75t_L g430 ( .A(n_359), .B(n_40), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_355), .B(n_96), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_355), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_364), .B(n_43), .Y(n_433) );
INVx4_ASAP7_75t_SL g434 ( .A(n_358), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_358), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_377), .A2(n_45), .B1(n_49), .B2(n_51), .Y(n_436) );
NOR3xp33_ASAP7_75t_SL g437 ( .A(n_358), .B(n_52), .C(n_53), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_364), .B(n_60), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_371), .B(n_376), .Y(n_439) );
OR2x6_ASAP7_75t_L g440 ( .A(n_380), .B(n_62), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_371), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_371), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_401), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_421), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_392), .B(n_376), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_407), .A2(n_366), .B(n_370), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_416), .B(n_376), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_398), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_383), .B(n_378), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_406), .B(n_378), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_394), .B(n_378), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_391), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_432), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_394), .B(n_372), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_424), .B(n_372), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_441), .B(n_442), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_411), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_386), .B(n_353), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_386), .B(n_439), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_387), .B(n_353), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_384), .B(n_357), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_387), .B(n_357), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_418), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_390), .B(n_357), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_413), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_405), .B(n_357), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_393), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_413), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_395), .B(n_366), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_410), .B(n_380), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_385), .B(n_380), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_385), .B(n_380), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_412), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_440), .B(n_375), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_440), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_440), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_426), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_412), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_409), .B(n_375), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_425), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_435), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_404), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_434), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_434), .Y(n_493) );
INVx4_ASAP7_75t_L g494 ( .A(n_423), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_397), .B(n_375), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_400), .B(n_375), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_427), .B(n_64), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_429), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_389), .B(n_370), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_429), .B(n_66), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_429), .Y(n_503) );
INVxp67_ASAP7_75t_L g504 ( .A(n_388), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_423), .B(n_67), .Y(n_505) );
BUFx3_ASAP7_75t_L g506 ( .A(n_402), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_423), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_415), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_408), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_436), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_419), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_414), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_430), .B(n_68), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_437), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_417), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_403), .B(n_69), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_411), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_392), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_421), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_392), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_385), .A2(n_70), .B1(n_72), .B2(n_73), .C1(n_76), .C2(n_77), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_392), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_421), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_421), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_396), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_392), .B(n_78), .Y(n_526) );
INVx5_ASAP7_75t_L g527 ( .A(n_423), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_421), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_392), .B(n_80), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_392), .B(n_81), .Y(n_530) );
AND2x4_ASAP7_75t_SL g531 ( .A(n_475), .B(n_83), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_494), .B(n_86), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_448), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_444), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_467), .B(n_89), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_453), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_448), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_462), .B(n_90), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_494), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_508), .A2(n_93), .B(n_94), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_467), .B(n_95), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_449), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_518), .Y(n_543) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_494), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_462), .B(n_461), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_469), .B(n_459), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_461), .B(n_454), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_520), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_521), .B(n_507), .C(n_497), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_469), .B(n_459), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_522), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_454), .B(n_455), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_455), .B(n_522), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_446), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_494), .B(n_527), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_446), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_451), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_470), .B(n_509), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_509), .B(n_488), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_509), .B(n_488), .Y(n_561) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_490), .B(n_508), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_451), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_527), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_456), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_456), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_443), .B(n_525), .Y(n_567) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_512), .B(n_511), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_521), .B(n_507), .C(n_501), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_460), .B(n_517), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_452), .B(n_450), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_485), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_445), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_460), .B(n_517), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_460), .B(n_517), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_452), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_450), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_476), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_476), .B(n_487), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_487), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_504), .B(n_498), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_464), .B(n_524), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_519), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_523), .B(n_528), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_481), .B(n_458), .Y(n_587) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_523), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_524), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_489), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_489), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_489), .B(n_481), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_524), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_458), .B(n_443), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_473), .B(n_528), .Y(n_595) );
NOR2xp33_ASAP7_75t_SL g596 ( .A(n_527), .B(n_490), .Y(n_596) );
NAND2xp33_ASAP7_75t_SL g597 ( .A(n_525), .B(n_491), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_463), .B(n_512), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_528), .B(n_479), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_506), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_463), .B(n_512), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_493), .Y(n_602) );
OAI221xp5_ASAP7_75t_SL g603 ( .A1(n_513), .A2(n_506), .B1(n_505), .B2(n_499), .C(n_474), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_479), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_479), .B(n_473), .Y(n_605) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_511), .B(n_491), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_466), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_493), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_465), .B(n_482), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_511), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_465), .B(n_482), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_498), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_486), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_483), .B(n_492), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_457), .B(n_482), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_466), .Y(n_616) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_516), .B(n_486), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_483), .B(n_492), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_501), .B(n_484), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_486), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_567), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_570), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_547), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_546), .B(n_480), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_547), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_612), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_574), .Y(n_627) );
NAND2xp33_ASAP7_75t_R g628 ( .A(n_567), .B(n_480), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_554), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_551), .B(n_457), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_598), .B(n_457), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_574), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_601), .B(n_457), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_537), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_600), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_545), .B(n_468), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_577), .B(n_468), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_618), .B(n_484), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_589), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_554), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_545), .B(n_468), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_619), .B(n_471), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_619), .B(n_471), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_582), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_609), .B(n_471), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_564), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_609), .B(n_478), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_589), .Y(n_649) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_569), .B(n_474), .C(n_477), .D(n_513), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_553), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_544), .B(n_478), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_565), .B(n_477), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_571), .B(n_478), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_611), .B(n_495), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_611), .B(n_495), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_553), .Y(n_657) );
AO22x1_ASAP7_75t_L g658 ( .A1(n_544), .A2(n_527), .B1(n_500), .B2(n_503), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_580), .B(n_472), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_597), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_594), .B(n_500), .Y(n_661) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_540), .B(n_527), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_587), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_587), .Y(n_664) );
INVx8_ASAP7_75t_L g665 ( .A(n_575), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_573), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_537), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_597), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_581), .B(n_472), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_571), .B(n_500), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_605), .B(n_447), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_566), .B(n_503), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_615), .B(n_503), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_559), .B(n_447), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_532), .B(n_499), .Y(n_675) );
NAND2xp67_ASAP7_75t_L g676 ( .A(n_606), .B(n_516), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_578), .B(n_447), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_610), .B(n_447), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_534), .B(n_510), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_595), .B(n_496), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_542), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_595), .B(n_527), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_555), .B(n_510), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_536), .B(n_558), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_583), .B(n_505), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_543), .Y(n_686) );
INVx4_ASAP7_75t_L g687 ( .A(n_531), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_548), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_590), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_536), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_592), .B(n_514), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_655), .B(n_572), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_621), .B(n_576), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_650), .B(n_603), .C(n_549), .D(n_596), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_655), .B(n_563), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_665), .Y(n_696) );
INVxp33_ASAP7_75t_L g697 ( .A(n_687), .Y(n_697) );
AOI32xp33_ASAP7_75t_L g698 ( .A1(n_660), .A2(n_596), .A3(n_617), .B1(n_591), .B2(n_582), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_635), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_637), .B(n_533), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_627), .Y(n_701) );
NAND4xp75_ASAP7_75t_L g702 ( .A(n_662), .B(n_562), .C(n_556), .D(n_532), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_645), .A2(n_562), .B1(n_560), .B2(n_561), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_627), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_656), .B(n_557), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_665), .Y(n_706) );
NOR2x1p5_ASAP7_75t_SL g707 ( .A(n_632), .B(n_620), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_651), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_657), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_632), .Y(n_710) );
AOI32xp33_ASAP7_75t_L g711 ( .A1(n_668), .A2(n_539), .A3(n_568), .B1(n_502), .B2(n_556), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_656), .B(n_614), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_642), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_687), .A2(n_603), .B1(n_539), .B2(n_608), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_665), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_642), .Y(n_716) );
NOR4xp25_ASAP7_75t_L g717 ( .A(n_666), .B(n_602), .C(n_538), .D(n_579), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_629), .Y(n_718) );
AOI21xp33_ASAP7_75t_SL g719 ( .A1(n_665), .A2(n_502), .B(n_514), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_621), .B(n_615), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_687), .B(n_538), .C(n_541), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_636), .B(n_613), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_633), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_621), .B(n_604), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_628), .A2(n_599), .B1(n_515), .B2(n_588), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_641), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_628), .A2(n_535), .B1(n_510), .B2(n_515), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_689), .B(n_616), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g729 ( .A1(n_675), .A2(n_588), .B(n_526), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_689), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_690), .Y(n_731) );
INVx2_ASAP7_75t_SL g732 ( .A(n_622), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_622), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_691), .A2(n_515), .B1(n_552), .B2(n_550), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_670), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_683), .B(n_607), .Y(n_736) );
OAI22xp33_ASAP7_75t_SL g737 ( .A1(n_676), .A2(n_585), .B1(n_593), .B2(n_584), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_643), .A2(n_515), .B1(n_586), .B2(n_529), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_643), .A2(n_515), .B1(n_526), .B2(n_529), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_654), .B(n_515), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_708), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_697), .A2(n_647), .B1(n_633), .B2(n_682), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_733), .Y(n_743) );
CKINVDCx14_ASAP7_75t_R g744 ( .A(n_693), .Y(n_744) );
OAI22xp33_ASAP7_75t_SL g745 ( .A1(n_696), .A2(n_647), .B1(n_633), .B2(n_684), .Y(n_745) );
OAI22x1_ASAP7_75t_L g746 ( .A1(n_730), .A2(n_647), .B1(n_640), .B2(n_652), .Y(n_746) );
AOI22x1_ASAP7_75t_L g747 ( .A1(n_706), .A2(n_630), .B1(n_667), .B2(n_674), .Y(n_747) );
INVx2_ASAP7_75t_SL g748 ( .A(n_715), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_694), .A2(n_714), .B1(n_721), .B2(n_737), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_709), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_703), .A2(n_630), .B1(n_624), .B2(n_639), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_720), .B(n_644), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_718), .Y(n_753) );
AOI211x1_ASAP7_75t_L g754 ( .A1(n_725), .A2(n_658), .B(n_624), .C(n_679), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_717), .A2(n_674), .B(n_671), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_711), .A2(n_653), .B(n_672), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_702), .A2(n_685), .B1(n_623), .B2(n_625), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g758 ( .A1(n_727), .A2(n_663), .B1(n_664), .B2(n_671), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_732), .A2(n_644), .B1(n_683), .B2(n_646), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_719), .A2(n_631), .B1(n_634), .B2(n_649), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_698), .A2(n_626), .B1(n_677), .B2(n_646), .C(n_648), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_728), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_726), .Y(n_763) );
AOI31xp33_ASAP7_75t_L g764 ( .A1(n_729), .A2(n_652), .A3(n_631), .B(n_634), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_731), .A2(n_677), .B1(n_648), .B2(n_669), .C(n_659), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_720), .A2(n_659), .B1(n_669), .B2(n_661), .Y(n_766) );
NAND4xp25_ASAP7_75t_L g767 ( .A(n_739), .B(n_652), .C(n_678), .D(n_673), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_749), .A2(n_734), .B1(n_722), .B2(n_699), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_744), .B(n_692), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_741), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_750), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_753), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_743), .B(n_713), .Y(n_773) );
AOI211x1_ASAP7_75t_L g774 ( .A1(n_755), .A2(n_712), .B(n_705), .C(n_695), .Y(n_774) );
AOI222xp33_ASAP7_75t_L g775 ( .A1(n_761), .A2(n_707), .B1(n_723), .B2(n_735), .C1(n_716), .C2(n_678), .Y(n_775) );
OAI21xp33_ASAP7_75t_SL g776 ( .A1(n_764), .A2(n_723), .B(n_738), .Y(n_776) );
INVxp67_ASAP7_75t_L g777 ( .A(n_748), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_763), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_759), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_752), .B(n_724), .Y(n_780) );
NOR2xp33_ASAP7_75t_SL g781 ( .A(n_747), .B(n_728), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_776), .B(n_757), .C(n_777), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_781), .A2(n_746), .B(n_745), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_781), .A2(n_742), .B(n_764), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_770), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_774), .B(n_754), .C(n_767), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_780), .B(n_762), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g788 ( .A1(n_779), .A2(n_758), .B1(n_767), .B2(n_760), .C(n_756), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g789 ( .A(n_782), .B(n_786), .C(n_788), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_787), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_785), .B(n_778), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_784), .A2(n_768), .B1(n_769), .B2(n_751), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_792), .A2(n_783), .B1(n_771), .B2(n_772), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_789), .B(n_775), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g795 ( .A1(n_790), .A2(n_765), .B(n_773), .C(n_766), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_794), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_793), .Y(n_797) );
OR5x1_ASAP7_75t_L g798 ( .A(n_797), .B(n_795), .C(n_791), .D(n_724), .E(n_740), .Y(n_798) );
INVx4_ASAP7_75t_L g799 ( .A(n_796), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_799), .A2(n_710), .B(n_704), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_798), .Y(n_801) );
OA22x2_ASAP7_75t_L g802 ( .A1(n_801), .A2(n_701), .B1(n_736), .B2(n_673), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_802), .A2(n_800), .B1(n_686), .B2(n_681), .Y(n_803) );
AOI22x1_ASAP7_75t_L g804 ( .A1(n_803), .A2(n_530), .B1(n_700), .B2(n_649), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_804), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_805), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_806), .A2(n_673), .B1(n_680), .B2(n_638), .Y(n_807) );
OR2x6_ASAP7_75t_L g808 ( .A(n_807), .B(n_530), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_808), .A2(n_680), .B1(n_638), .B2(n_688), .Y(n_809) );
endmodule