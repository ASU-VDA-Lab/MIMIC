module fake_ariane_977_n_179 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_179);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_179;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_162;
wire n_112;
wire n_45;
wire n_138;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVxp33_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_R g60 ( 
.A(n_37),
.B(n_15),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_4),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_5),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_34),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_42),
.Y(n_82)
);

AOI22x1_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_50),
.B1(n_49),
.B2(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_55),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_5),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_73),
.Y(n_99)
);

NAND2x1p5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_85),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_58),
.B(n_60),
.C(n_63),
.Y(n_101)
);

AND3x1_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_67),
.C(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_61),
.B1(n_62),
.B2(n_6),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_12),
.B1(n_19),
.B2(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_27),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_30),
.B(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_81),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_88),
.B1(n_96),
.B2(n_85),
.Y(n_115)
);

AO21x2_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_87),
.B(n_80),
.Y(n_116)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_83),
.B(n_87),
.Y(n_117)
);

NAND2x1p5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_92),
.B(n_91),
.Y(n_121)
);

OAI21x1_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_92),
.B(n_91),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_91),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_113),
.B(n_98),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_115),
.B(n_103),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_106),
.B(n_102),
.Y(n_129)
);

OAI21x1_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_103),
.B(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_112),
.B(n_99),
.Y(n_132)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_112),
.B(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_128),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_131),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_130),
.Y(n_136)
);

AND4x1_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_130),
.C(n_129),
.D(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_R g138 ( 
.A(n_129),
.B(n_123),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_121),
.C(n_118),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_121),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_116),
.B(n_132),
.C(n_133),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_145),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

OR2x6_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_153),
.Y(n_162)
);

OR2x6_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_153),
.Y(n_163)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_152),
.B(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_163),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_164),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_163),
.B(n_162),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_162),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_155),
.B1(n_138),
.B2(n_157),
.C(n_143),
.Y(n_171)
);

INVxp33_ASAP7_75t_SL g172 ( 
.A(n_170),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_150),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_172),
.B1(n_150),
.B2(n_137),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_160),
.B1(n_146),
.B2(n_116),
.C(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_154),
.B1(n_141),
.B2(n_127),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_117),
.B(n_132),
.Y(n_179)
);


endmodule