module fake_jpeg_2278_n_517 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_3),
.B(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_52),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_54),
.B(n_44),
.Y(n_159)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_63),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_67),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_85),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_18),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_93),
.Y(n_132)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx2_ASAP7_75t_R g96 ( 
.A(n_41),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_24),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_109),
.B(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_24),
.B1(n_17),
.B2(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_111),
.A2(n_42),
.B1(n_96),
.B2(n_75),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_40),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_119),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_86),
.B(n_46),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_131),
.B(n_159),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_50),
.A2(n_17),
.B1(n_42),
.B2(n_46),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_27),
.B1(n_14),
.B2(n_71),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_67),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_70),
.B1(n_27),
.B2(n_31),
.Y(n_169)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_48),
.B(n_69),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_84),
.B(n_31),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_64),
.B(n_43),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_161),
.B(n_72),
.Y(n_210)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_164),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_84),
.B(n_14),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_178),
.Y(n_215)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_169),
.A2(n_184),
.B1(n_204),
.B2(n_209),
.Y(n_245)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx3_ASAP7_75t_SL g228 ( 
.A(n_170),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_119),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_28),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_174),
.Y(n_231)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_28),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_36),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_177),
.B(n_185),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_103),
.B(n_88),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_179),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_180),
.A2(n_205),
.B1(n_115),
.B2(n_80),
.Y(n_229)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_103),
.A2(n_98),
.B1(n_36),
.B2(n_23),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_23),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_40),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_194),
.Y(n_248)
);

INVx5_ASAP7_75t_SL g189 ( 
.A(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_74),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_104),
.Y(n_214)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_115),
.B1(n_138),
.B2(n_127),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_122),
.B(n_99),
.Y(n_194)
);

CKINVDCx12_ASAP7_75t_R g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_121),
.A2(n_97),
.B(n_92),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_208),
.Y(n_216)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_202),
.Y(n_226)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_207),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_128),
.A2(n_51),
.B1(n_78),
.B2(n_100),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_143),
.A2(n_59),
.B1(n_101),
.B2(n_94),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_105),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g209 ( 
.A(n_124),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_210),
.B(n_212),
.Y(n_222)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_140),
.B1(n_123),
.B2(n_155),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_77),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_139),
.B1(n_127),
.B2(n_113),
.Y(n_213)
);

AO22x1_ASAP7_75t_SL g258 ( 
.A1(n_213),
.A2(n_218),
.B1(n_179),
.B2(n_191),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_214),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_138),
.B1(n_112),
.B2(n_113),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_221),
.A2(n_189),
.B1(n_179),
.B2(n_136),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_172),
.B(n_158),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_232),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_188),
.B(n_135),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_120),
.B1(n_112),
.B2(n_125),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_244),
.B1(n_208),
.B2(n_207),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_125),
.B1(n_155),
.B2(n_137),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_186),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_251),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_165),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_253),
.A2(n_214),
.B1(n_218),
.B2(n_220),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_174),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_185),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_176),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_265),
.C(n_268),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_197),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_264),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_216),
.A2(n_171),
.B1(n_194),
.B2(n_137),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_195),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_266),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_231),
.B(n_200),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_171),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_263),
.B(n_278),
.Y(n_289)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_178),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_237),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_252),
.B1(n_275),
.B2(n_278),
.Y(n_284)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_189),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_274),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_213),
.A2(n_191),
.B1(n_66),
.B2(n_65),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_229),
.B1(n_242),
.B2(n_238),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_182),
.B(n_168),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_221),
.B(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_173),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_238),
.C(n_248),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_298),
.C(n_303),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_274),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_284),
.A2(n_267),
.B1(n_270),
.B2(n_228),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_287),
.A2(n_301),
.B(n_302),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_289),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_297),
.B1(n_308),
.B2(n_252),
.Y(n_314)
);

INVx11_ASAP7_75t_SL g295 ( 
.A(n_279),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_295),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_259),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_252),
.A2(n_232),
.B1(n_239),
.B2(n_226),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_214),
.C(n_227),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_214),
.B(n_225),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_258),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_257),
.A2(n_214),
.B(n_227),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_230),
.C(n_234),
.Y(n_303)
);

XOR2x2_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_151),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_152),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_256),
.B(n_259),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_240),
.C(n_230),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_252),
.A2(n_275),
.B1(n_269),
.B2(n_264),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_320),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_314),
.A2(n_316),
.B1(n_319),
.B2(n_329),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_315),
.A2(n_328),
.B(n_302),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_253),
.B1(n_269),
.B2(n_251),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_289),
.A2(n_276),
.B(n_260),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_318),
.A2(n_336),
.B(n_338),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_281),
.A2(n_272),
.B1(n_258),
.B2(n_277),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_255),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_272),
.B1(n_258),
.B2(n_254),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_321),
.A2(n_297),
.B1(n_303),
.B2(n_294),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_327),
.Y(n_349)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_268),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_304),
.A2(n_225),
.B(n_266),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_258),
.B1(n_267),
.B2(n_273),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_243),
.C(n_240),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_333),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_340),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_273),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_304),
.Y(n_334)
);

BUFx4f_ASAP7_75t_SL g368 ( 
.A(n_334),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_293),
.B(n_270),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_335),
.B(n_285),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_307),
.A2(n_236),
.B(n_181),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_233),
.C(n_234),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_332),
.C(n_333),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_307),
.A2(n_236),
.B(n_235),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_339),
.Y(n_344)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_298),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_348),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_303),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_352),
.B(n_356),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_351),
.A2(n_359),
.B1(n_322),
.B2(n_319),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_313),
.A2(n_300),
.B(n_283),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_357),
.C(n_312),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_313),
.A2(n_291),
.B(n_301),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_291),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_318),
.A2(n_305),
.B(n_287),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_372),
.B(n_315),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_290),
.B1(n_305),
.B2(n_293),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_367),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_312),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_340),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_323),
.B(n_306),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_371),
.B(n_320),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_315),
.A2(n_310),
.B(n_285),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_351),
.A2(n_316),
.B1(n_314),
.B2(n_322),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_356),
.B1(n_347),
.B2(n_358),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_378),
.A2(n_384),
.B1(n_394),
.B2(n_395),
.Y(n_415)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_334),
.Y(n_381)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_327),
.B1(n_331),
.B2(n_329),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_385),
.A2(n_354),
.B(n_309),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_386),
.B(n_397),
.Y(n_423)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_317),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_391),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_219),
.Y(n_417)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_345),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_317),
.B1(n_330),
.B2(n_326),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_362),
.A2(n_338),
.B1(n_341),
.B2(n_288),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_233),
.C(n_235),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_398),
.C(n_353),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_224),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_348),
.B(n_219),
.C(n_309),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_357),
.B(n_224),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_361),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_404),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_345),
.C(n_372),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_414),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_352),
.B(n_347),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_416),
.B(n_418),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_365),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_421),
.Y(n_425)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_410),
.A2(n_422),
.B1(n_391),
.B2(n_394),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_395),
.A2(n_367),
.B1(n_343),
.B2(n_350),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_382),
.B1(n_374),
.B2(n_373),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_366),
.C(n_342),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_419),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_382),
.A2(n_373),
.B(n_374),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_267),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_147),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_375),
.A2(n_206),
.B1(n_228),
.B2(n_108),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_376),
.Y(n_426)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_426),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_427),
.A2(n_429),
.B1(n_432),
.B2(n_424),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_376),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_428),
.B(n_434),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g429 ( 
.A(n_413),
.B(n_392),
.CI(n_381),
.CON(n_429),
.SN(n_429)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_430),
.A2(n_433),
.B1(n_443),
.B2(n_142),
.Y(n_463)
);

AOI321xp33_ASAP7_75t_L g432 ( 
.A1(n_411),
.A2(n_393),
.A3(n_379),
.B1(n_388),
.B2(n_387),
.C(n_383),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_410),
.A2(n_389),
.B1(n_377),
.B2(n_380),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_423),
.Y(n_434)
);

INVx13_ASAP7_75t_L g435 ( 
.A(n_424),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_435),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_249),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_409),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_202),
.C(n_199),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_444),
.C(n_445),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_150),
.B1(n_156),
.B2(n_146),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_441),
.A2(n_136),
.B1(n_144),
.B2(n_146),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_403),
.A2(n_249),
.B1(n_241),
.B2(n_120),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_211),
.C(n_201),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_198),
.C(n_190),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_437),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_452),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_405),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_454),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_449),
.A2(n_456),
.B1(n_90),
.B2(n_73),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_416),
.C(n_418),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_455),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_421),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_422),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_427),
.A2(n_420),
.B1(n_412),
.B2(n_406),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_442),
.A2(n_409),
.B1(n_220),
.B2(n_166),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_458),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_439),
.A2(n_156),
.B1(n_150),
.B2(n_144),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_170),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_460),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_58),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_463),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_175),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_464),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_439),
.C(n_444),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_470),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_435),
.B1(n_441),
.B2(n_429),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_463),
.A2(n_429),
.B1(n_432),
.B2(n_445),
.Y(n_471)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_443),
.C(n_168),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_476),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_449),
.A2(n_192),
.B(n_123),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_475),
.A2(n_461),
.B(n_167),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_448),
.C(n_451),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_79),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_102),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_140),
.C(n_81),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_1),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

AOI31xp67_ASAP7_75t_L g482 ( 
.A1(n_467),
.A2(n_450),
.A3(n_476),
.B(n_472),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_482),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_466),
.A2(n_454),
.B(n_456),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_484),
.B(n_490),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_468),
.A2(n_465),
.B(n_475),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_489),
.Y(n_501)
);

AOI321xp33_ASAP7_75t_L g487 ( 
.A1(n_465),
.A2(n_102),
.A3(n_62),
.B1(n_57),
.B2(n_39),
.C(n_4),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_488),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_0),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_480),
.A2(n_1),
.B(n_2),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_478),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_486),
.A2(n_474),
.B1(n_477),
.B2(n_469),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_495),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_481),
.B(n_477),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_6),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_481),
.B(n_479),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_498),
.A2(n_2),
.B(n_3),
.Y(n_503)
);

AOI322xp5_ASAP7_75t_L g499 ( 
.A1(n_493),
.A2(n_491),
.A3(n_469),
.B1(n_492),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_2),
.B(n_4),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_503),
.B(n_504),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_2),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_508),
.C(n_502),
.Y(n_509)
);

AO21x1_ASAP7_75t_L g507 ( 
.A1(n_497),
.A2(n_4),
.B(n_5),
.Y(n_507)
);

MAJx2_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_500),
.C(n_501),
.Y(n_511)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_509),
.A2(n_511),
.B(n_496),
.Y(n_513)
);

NOR3xp33_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_505),
.C(n_501),
.Y(n_512)
);

AOI322xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_513),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_514)
);

A2O1A1Ixp33_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_515)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_7),
.B(n_8),
.Y(n_516)
);

O2A1O1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_516),
.A2(n_8),
.B(n_10),
.C(n_223),
.Y(n_517)
);


endmodule