module real_aes_1812_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_626;
wire n_400;
wire n_539;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_727;
wire n_397;
wire n_749;
wire n_358;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_0), .A2(n_213), .B1(n_414), .B2(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_1), .A2(n_284), .B1(n_396), .B2(n_646), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_2), .A2(n_58), .B1(n_460), .B2(n_461), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_3), .A2(n_109), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_4), .A2(n_117), .B1(n_565), .B2(n_566), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_5), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_6), .A2(n_233), .B1(n_457), .B2(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_7), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_8), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_9), .A2(n_318), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_10), .A2(n_49), .B1(n_413), .B2(n_829), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_11), .A2(n_188), .B1(n_411), .B2(n_501), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_12), .A2(n_225), .B1(n_646), .B2(n_783), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_13), .A2(n_238), .B1(n_461), .B2(n_583), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_14), .A2(n_294), .B1(n_633), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_15), .A2(n_126), .B1(n_460), .B2(n_461), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_16), .A2(n_169), .B1(n_415), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_17), .A2(n_307), .B1(n_471), .B2(n_520), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_18), .A2(n_174), .B1(n_632), .B2(n_887), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_19), .A2(n_237), .B1(n_471), .B2(n_520), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_20), .B(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_21), .A2(n_271), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_22), .A2(n_203), .B1(n_465), .B2(n_672), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_23), .A2(n_129), .B1(n_465), .B2(n_672), .Y(n_785) );
INVx1_ASAP7_75t_SL g369 ( .A(n_24), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_24), .B(n_38), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_25), .A2(n_110), .B1(n_517), .B2(n_518), .Y(n_606) );
AOI22xp5_ASAP7_75t_SL g767 ( .A1(n_26), .A2(n_239), .B1(n_507), .B2(n_768), .Y(n_767) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_27), .A2(n_288), .B1(n_322), .B2(n_467), .C1(n_469), .C2(n_472), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_28), .B(n_547), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_29), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_30), .A2(n_317), .B1(n_423), .B2(n_748), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_31), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_32), .A2(n_275), .B1(n_463), .B2(n_651), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_33), .A2(n_219), .B1(n_573), .B2(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_34), .A2(n_101), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_35), .A2(n_95), .B1(n_454), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_36), .A2(n_94), .B1(n_573), .B2(n_768), .Y(n_889) );
INVx1_ASAP7_75t_L g932 ( .A(n_37), .Y(n_932) );
AO22x2_ASAP7_75t_L g371 ( .A1(n_38), .A2(n_327), .B1(n_368), .B2(n_372), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_39), .A2(n_197), .B1(n_565), .B2(n_630), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_40), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_41), .A2(n_272), .B1(n_526), .B2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_42), .A2(n_103), .B1(n_573), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_43), .A2(n_87), .B1(n_526), .B2(n_590), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_44), .A2(n_255), .B1(n_420), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_45), .A2(n_262), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_46), .A2(n_258), .B1(n_391), .B2(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g370 ( .A(n_47), .Y(n_370) );
AO222x2_ASAP7_75t_SL g603 ( .A1(n_48), .A2(n_189), .B1(n_266), .B2(n_468), .C1(n_471), .C2(n_520), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_50), .A2(n_319), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g754 ( .A(n_51), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_52), .A2(n_231), .B1(n_532), .B2(n_533), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_53), .A2(n_92), .B1(n_411), .B2(n_414), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_54), .A2(n_299), .B1(n_526), .B2(n_590), .Y(n_903) );
AO222x2_ASAP7_75t_SL g580 ( .A1(n_55), .A2(n_114), .B1(n_148), .B2(n_468), .C1(n_471), .C2(n_520), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_56), .A2(n_273), .B1(n_401), .B2(n_493), .Y(n_744) );
AO22x2_ASAP7_75t_L g378 ( .A1(n_57), .A2(n_180), .B1(n_368), .B2(n_379), .Y(n_378) );
XNOR2x1_ASAP7_75t_L g616 ( .A(n_59), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_60), .A2(n_65), .B1(n_530), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_61), .A2(n_298), .B1(n_428), .B2(n_501), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_62), .B(n_486), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_63), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_64), .A2(n_325), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI221x1_ASAP7_75t_L g631 ( .A1(n_66), .A2(n_74), .B1(n_632), .B2(n_633), .C(n_634), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_67), .A2(n_143), .B1(n_532), .B2(n_533), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_68), .A2(n_228), .B1(n_678), .B2(n_965), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_69), .A2(n_257), .B1(n_461), .B2(n_583), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_70), .A2(n_308), .B1(n_401), .B2(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_71), .A2(n_145), .B1(n_448), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_72), .A2(n_304), .B1(n_528), .B2(n_530), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_73), .A2(n_243), .B1(n_457), .B2(n_502), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_75), .B(n_467), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_76), .A2(n_232), .B1(n_436), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_77), .A2(n_253), .B1(n_439), .B2(n_530), .Y(n_907) );
INVx1_ASAP7_75t_L g637 ( .A(n_78), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_79), .A2(n_348), .B1(n_532), .B2(n_533), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_80), .A2(n_230), .B1(n_650), .B2(n_832), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_81), .A2(n_108), .B1(n_415), .B2(n_454), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_82), .A2(n_241), .B1(n_457), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_83), .A2(n_305), .B1(n_450), .B2(n_887), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_84), .A2(n_935), .B1(n_950), .B2(n_951), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_84), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_85), .A2(n_183), .B1(n_559), .B2(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_86), .B(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_88), .A2(n_127), .B1(n_441), .B2(n_457), .Y(n_812) );
INVx1_ASAP7_75t_L g644 ( .A(n_89), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_90), .A2(n_277), .B1(n_558), .B2(n_655), .Y(n_969) );
INVx1_ASAP7_75t_L g623 ( .A(n_91), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_93), .A2(n_290), .B1(n_517), .B2(n_586), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_96), .A2(n_222), .B1(n_592), .B2(n_595), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_97), .A2(n_309), .B1(n_460), .B2(n_584), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_98), .A2(n_340), .B1(n_694), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_99), .A2(n_276), .B1(n_572), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_100), .A2(n_310), .B1(n_528), .B2(n_530), .Y(n_813) );
AOI222xp33_ASAP7_75t_L g970 ( .A1(n_102), .A2(n_161), .B1(n_313), .B2(n_396), .C1(n_487), .C2(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_104), .A2(n_130), .B1(n_401), .B2(n_556), .Y(n_938) );
OAI22x1_ASAP7_75t_L g356 ( .A1(n_105), .A2(n_357), .B1(n_358), .B2(n_442), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_105), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_106), .A2(n_234), .B1(n_436), .B2(n_507), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_107), .A2(n_247), .B1(n_498), .B2(n_650), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_111), .A2(n_301), .B1(n_504), .B2(n_505), .Y(n_503) );
AO22x2_ASAP7_75t_L g375 ( .A1(n_112), .A2(n_263), .B1(n_368), .B2(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_113), .A2(n_208), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_115), .A2(n_186), .B1(n_428), .B2(n_432), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_116), .A2(n_195), .B1(n_791), .B2(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_118), .A2(n_344), .B1(n_765), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_119), .A2(n_160), .B1(n_471), .B2(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_120), .A2(n_323), .B1(n_528), .B2(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g972 ( .A(n_121), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_122), .A2(n_135), .B1(n_381), .B2(n_386), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_123), .A2(n_246), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_124), .A2(n_141), .B1(n_559), .B2(n_674), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_125), .A2(n_152), .B1(n_517), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_128), .A2(n_194), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_131), .A2(n_292), .B1(n_471), .B2(n_472), .Y(n_897) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_132), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_133), .A2(n_274), .B1(n_533), .B2(n_816), .Y(n_853) );
XOR2x2_ASAP7_75t_L g663 ( .A(n_134), .B(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_136), .A2(n_293), .B1(n_532), .B2(n_533), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_137), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_138), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_139), .A2(n_156), .B1(n_497), .B2(n_498), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_140), .B(n_487), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_142), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_144), .A2(n_209), .B1(n_526), .B2(n_590), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_146), .A2(n_164), .B1(n_592), .B2(n_595), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_147), .A2(n_329), .B1(n_517), .B2(n_586), .Y(n_899) );
INVx1_ASAP7_75t_L g622 ( .A(n_149), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_150), .A2(n_240), .B1(n_621), .B2(n_680), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_151), .A2(n_334), .B1(n_401), .B2(n_405), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_153), .A2(n_187), .B1(n_654), .B2(n_655), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_154), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_155), .A2(n_223), .B1(n_454), .B2(n_455), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_157), .A2(n_264), .B1(n_450), .B2(n_451), .Y(n_449) );
XNOR2x1_ASAP7_75t_L g482 ( .A(n_158), .B(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_159), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_162), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_163), .A2(n_324), .B1(n_528), .B2(n_530), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_165), .A2(n_201), .B1(n_526), .B2(n_590), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_166), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_167), .A2(n_217), .B1(n_498), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_168), .A2(n_227), .B1(n_450), .B2(n_680), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_170), .A2(n_191), .B1(n_401), .B2(n_556), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_171), .A2(n_229), .B1(n_436), .B2(n_439), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_172), .A2(n_216), .B1(n_411), .B2(n_414), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g896 ( .A(n_173), .B(n_487), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_175), .A2(n_303), .B1(n_455), .B2(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_176), .A2(n_268), .B1(n_491), .B2(n_551), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_177), .A2(n_248), .B1(n_502), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_178), .A2(n_341), .B1(n_526), .B2(n_590), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_179), .A2(n_224), .B1(n_621), .B2(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g921 ( .A(n_180), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_181), .A2(n_244), .B1(n_583), .B2(n_584), .Y(n_867) );
INVx1_ASAP7_75t_L g627 ( .A(n_182), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_184), .A2(n_332), .B1(n_533), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_185), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_190), .A2(n_282), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_192), .A2(n_337), .B1(n_505), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_193), .A2(n_226), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_196), .A2(n_345), .B1(n_572), .B2(n_573), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_198), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_199), .A2(n_343), .B1(n_471), .B2(n_520), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_200), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_202), .A2(n_220), .B1(n_396), .B2(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_204), .A2(n_349), .B1(n_448), .B2(n_678), .Y(n_789) );
INVx2_ASAP7_75t_L g931 ( .A(n_205), .Y(n_931) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_206), .B(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_207), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_210), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_211), .A2(n_235), .B1(n_762), .B2(n_829), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_212), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_214), .A2(n_236), .B1(n_528), .B2(n_530), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_215), .A2(n_316), .B1(n_465), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_218), .A2(n_283), .B1(n_532), .B2(n_533), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_221), .A2(n_306), .B1(n_583), .B2(n_584), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_242), .B(n_758), .Y(n_878) );
INVx1_ASAP7_75t_L g626 ( .A(n_245), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_249), .A2(n_297), .B1(n_741), .B2(n_742), .Y(n_740) );
OA22x2_ASAP7_75t_L g443 ( .A1(n_250), .A2(n_444), .B1(n_445), .B2(n_473), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_250), .Y(n_444) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_250), .A2(n_445), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g890 ( .A(n_251), .Y(n_890) );
XNOR2xp5_ASAP7_75t_L g858 ( .A(n_252), .B(n_859), .Y(n_858) );
AOI22x1_ASAP7_75t_L g577 ( .A1(n_254), .A2(n_578), .B1(n_597), .B2(n_598), .Y(n_577) );
INVx1_ASAP7_75t_L g598 ( .A(n_254), .Y(n_598) );
XNOR2x1_ASAP7_75t_L g779 ( .A(n_256), .B(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_259), .A2(n_265), .B1(n_381), .B2(n_493), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_260), .A2(n_315), .B1(n_768), .B2(n_773), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_261), .B(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_263), .B(n_920), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_267), .A2(n_289), .B1(n_457), .B2(n_528), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_269), .B(n_362), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_270), .A2(n_338), .B1(n_517), .B2(n_518), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_278), .A2(n_342), .B1(n_418), .B2(n_423), .Y(n_417) );
OA22x2_ASAP7_75t_L g794 ( .A1(n_279), .A2(n_795), .B1(n_796), .B2(n_818), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_279), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_280), .A2(n_296), .B1(n_505), .B2(n_947), .Y(n_946) );
INVx3_ASAP7_75t_L g368 ( .A(n_281), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_285), .Y(n_719) );
INVx1_ASAP7_75t_L g638 ( .A(n_286), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_287), .A2(n_320), .B1(n_694), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_291), .A2(n_300), .B1(n_391), .B2(n_396), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_295), .A2(n_339), .B1(n_463), .B2(n_465), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_302), .Y(n_724) );
INVx1_ASAP7_75t_L g647 ( .A(n_311), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_312), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_314), .A2(n_321), .B1(n_764), .B2(n_765), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_326), .B(n_547), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_328), .A2(n_335), .B1(n_654), .B2(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_330), .B(n_486), .Y(n_739) );
INVx1_ASAP7_75t_L g916 ( .A(n_331), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g930 ( .A(n_331), .B(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g917 ( .A(n_333), .Y(n_917) );
AND2x2_ASAP7_75t_R g953 ( .A(n_333), .B(n_916), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_336), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g641 ( .A(n_346), .Y(n_641) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_347), .B(n_543), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_912), .B(n_923), .Y(n_350) );
AO21x1_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_728), .B(n_730), .Y(n_351) );
AOI31xp33_ASAP7_75t_L g912 ( .A1(n_352), .A2(n_728), .A3(n_730), .B(n_913), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_538), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_354), .B(n_729), .Y(n_728) );
AO22x2_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_479), .B1(n_536), .B2(n_537), .Y(n_354) );
INVx2_ASAP7_75t_SL g536 ( .A(n_355), .Y(n_536) );
OA22x2_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_443), .B1(n_474), .B2(n_475), .Y(n_355) );
INVx1_ASAP7_75t_SL g474 ( .A(n_356), .Y(n_474) );
INVx2_ASAP7_75t_SL g442 ( .A(n_358), .Y(n_442) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_409), .Y(n_358) );
NAND4xp25_ASAP7_75t_SL g359 ( .A(n_360), .B(n_380), .C(n_390), .D(n_400), .Y(n_359) );
INVx3_ASAP7_75t_L g642 ( .A(n_361), .Y(n_642) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_SL g487 ( .A(n_363), .Y(n_487) );
INVx4_ASAP7_75t_SL g547 ( .A(n_363), .Y(n_547) );
BUFx2_ASAP7_75t_L g667 ( .A(n_363), .Y(n_667) );
INVx3_ASAP7_75t_L g758 ( .A(n_363), .Y(n_758) );
INVx6_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_373), .Y(n_364) );
AND2x4_ASAP7_75t_L g388 ( .A(n_365), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g406 ( .A(n_365), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g461 ( .A(n_365), .B(n_389), .Y(n_461) );
AND2x4_ASAP7_75t_L g468 ( .A(n_365), .B(n_373), .Y(n_468) );
AND2x2_ASAP7_75t_L g518 ( .A(n_365), .B(n_407), .Y(n_518) );
AND2x2_ASAP7_75t_L g584 ( .A(n_365), .B(n_389), .Y(n_584) );
AND2x2_ASAP7_75t_L g586 ( .A(n_365), .B(n_407), .Y(n_586) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_371), .Y(n_365) );
INVx2_ASAP7_75t_L g385 ( .A(n_366), .Y(n_385) );
AND2x2_ASAP7_75t_L g394 ( .A(n_366), .B(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
OAI22x1_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_369), .B2(n_370), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g372 ( .A(n_368), .Y(n_372) );
INVx2_ASAP7_75t_L g376 ( .A(n_368), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_368), .Y(n_379) );
AND2x2_ASAP7_75t_L g384 ( .A(n_371), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
BUFx2_ASAP7_75t_L g426 ( .A(n_371), .Y(n_426) );
AND2x4_ASAP7_75t_L g413 ( .A(n_373), .B(n_394), .Y(n_413) );
AND2x4_ASAP7_75t_L g431 ( .A(n_373), .B(n_416), .Y(n_431) );
AND2x2_ASAP7_75t_L g438 ( .A(n_373), .B(n_384), .Y(n_438) );
AND2x6_ASAP7_75t_L g530 ( .A(n_373), .B(n_384), .Y(n_530) );
AND2x2_ASAP7_75t_L g532 ( .A(n_373), .B(n_394), .Y(n_532) );
AND2x2_ASAP7_75t_L g592 ( .A(n_373), .B(n_416), .Y(n_592) );
AND2x2_ASAP7_75t_L g816 ( .A(n_373), .B(n_394), .Y(n_816) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g383 ( .A(n_375), .B(n_377), .Y(n_383) );
AND2x2_ASAP7_75t_L g398 ( .A(n_375), .B(n_378), .Y(n_398) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
INVxp67_ASAP7_75t_L g389 ( .A(n_377), .Y(n_389) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g403 ( .A(n_378), .B(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g497 ( .A(n_381), .Y(n_497) );
BUFx2_ASAP7_75t_L g654 ( .A(n_381), .Y(n_654) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g558 ( .A(n_382), .Y(n_558) );
BUFx3_ASAP7_75t_L g674 ( .A(n_382), .Y(n_674) );
BUFx2_ASAP7_75t_L g880 ( .A(n_382), .Y(n_880) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g393 ( .A(n_383), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g441 ( .A(n_383), .B(n_416), .Y(n_441) );
AND2x2_ASAP7_75t_L g460 ( .A(n_383), .B(n_384), .Y(n_460) );
AND2x4_ASAP7_75t_L g471 ( .A(n_383), .B(n_394), .Y(n_471) );
AND2x2_ASAP7_75t_L g583 ( .A(n_383), .B(n_384), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_383), .B(n_416), .Y(n_595) );
AND2x2_ASAP7_75t_L g422 ( .A(n_384), .B(n_403), .Y(n_422) );
AND2x2_ASAP7_75t_L g525 ( .A(n_384), .B(n_403), .Y(n_525) );
AND2x2_ASAP7_75t_SL g590 ( .A(n_384), .B(n_403), .Y(n_590) );
AND2x4_ASAP7_75t_L g416 ( .A(n_385), .B(n_395), .Y(n_416) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g498 ( .A(n_387), .Y(n_498) );
INVx2_ASAP7_75t_L g559 ( .A(n_387), .Y(n_559) );
INVx2_ASAP7_75t_L g655 ( .A(n_387), .Y(n_655) );
INVx2_ASAP7_75t_SL g832 ( .A(n_387), .Y(n_832) );
INVx6_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g646 ( .A(n_392), .Y(n_646) );
INVx1_ASAP7_75t_L g971 ( .A(n_392), .Y(n_971) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g491 ( .A(n_393), .Y(n_491) );
BUFx3_ASAP7_75t_L g550 ( .A(n_393), .Y(n_550) );
AND2x2_ASAP7_75t_L g402 ( .A(n_394), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g517 ( .A(n_394), .B(n_403), .Y(n_517) );
INVx2_ASAP7_75t_L g643 ( .A(n_396), .Y(n_643) );
BUFx3_ASAP7_75t_L g771 ( .A(n_396), .Y(n_771) );
BUFx12f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g552 ( .A(n_397), .Y(n_552) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
AND2x4_ASAP7_75t_L g415 ( .A(n_398), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g425 ( .A(n_398), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_398), .B(n_399), .Y(n_472) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_398), .B(n_399), .Y(n_520) );
AND2x4_ASAP7_75t_L g526 ( .A(n_398), .B(n_426), .Y(n_526) );
AND2x4_ASAP7_75t_L g533 ( .A(n_398), .B(n_416), .Y(n_533) );
BUFx6f_ASAP7_75t_SL g650 ( .A(n_401), .Y(n_650) );
INVx1_ASAP7_75t_L g803 ( .A(n_401), .Y(n_803) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g464 ( .A(n_402), .Y(n_464) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_402), .Y(n_672) );
AND2x4_ASAP7_75t_L g434 ( .A(n_403), .B(n_416), .Y(n_434) );
AND2x6_ASAP7_75t_L g528 ( .A(n_403), .B(n_416), .Y(n_528) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_404), .Y(n_408) );
BUFx4f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
INVx2_ASAP7_75t_L g495 ( .A(n_406), .Y(n_495) );
BUFx6f_ASAP7_75t_SL g556 ( .A(n_406), .Y(n_556) );
INVx1_ASAP7_75t_L g652 ( .A(n_406), .Y(n_652) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_417), .C(n_427), .D(n_435), .Y(n_409) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_412), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_412), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
INVx2_ASAP7_75t_L g762 ( .A(n_412), .Y(n_762) );
INVx3_ASAP7_75t_L g791 ( .A(n_412), .Y(n_791) );
INVx6_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g570 ( .A(n_415), .Y(n_570) );
BUFx2_ASAP7_75t_SL g633 ( .A(n_415), .Y(n_633) );
BUFx3_ASAP7_75t_L g793 ( .A(n_415), .Y(n_793) );
BUFx3_ASAP7_75t_L g829 ( .A(n_415), .Y(n_829) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g764 ( .A(n_419), .Y(n_764) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_420), .Y(n_504) );
INVx1_ASAP7_75t_L g636 ( .A(n_420), .Y(n_636) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g563 ( .A(n_421), .Y(n_563) );
INVx1_ASAP7_75t_L g947 ( .A(n_421), .Y(n_947) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_422), .Y(n_678) );
BUFx3_ASAP7_75t_L g885 ( .A(n_422), .Y(n_885) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_424), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_424), .A2(n_700), .B1(n_701), .B2(n_703), .Y(n_699) );
INVx2_ASAP7_75t_L g965 ( .A(n_424), .Y(n_965) );
INVx5_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g505 ( .A(n_425), .Y(n_505) );
BUFx2_ASAP7_75t_L g749 ( .A(n_425), .Y(n_749) );
BUFx3_ASAP7_75t_L g765 ( .A(n_425), .Y(n_765) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g510 ( .A(n_429), .Y(n_510) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g457 ( .A(n_430), .Y(n_457) );
INVx2_ASAP7_75t_SL g572 ( .A(n_430), .Y(n_572) );
INVx3_ASAP7_75t_SL g632 ( .A(n_430), .Y(n_632) );
INVx2_ASAP7_75t_L g768 ( .A(n_430), .Y(n_768) );
INVx2_ASAP7_75t_SL g961 ( .A(n_430), .Y(n_961) );
INVx8_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
INVx2_ASAP7_75t_L g507 ( .A(n_433), .Y(n_507) );
INVx2_ASAP7_75t_L g566 ( .A(n_433), .Y(n_566) );
INVx2_ASAP7_75t_L g680 ( .A(n_433), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_433), .A2(n_705), .B1(n_706), .B2(n_709), .Y(n_704) );
INVx2_ASAP7_75t_SL g887 ( .A(n_433), .Y(n_887) );
INVx2_ASAP7_75t_L g962 ( .A(n_433), .Y(n_962) );
INVx8_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g450 ( .A(n_437), .Y(n_450) );
INVx2_ASAP7_75t_L g565 ( .A(n_437), .Y(n_565) );
INVx2_ASAP7_75t_L g708 ( .A(n_437), .Y(n_708) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g621 ( .A(n_438), .Y(n_621) );
BUFx2_ASAP7_75t_L g683 ( .A(n_438), .Y(n_683) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g455 ( .A(n_440), .Y(n_455) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_441), .Y(n_573) );
BUFx3_ASAP7_75t_L g630 ( .A(n_441), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_443), .A2(n_475), .B1(n_482), .B2(n_511), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_444), .Y(n_478) );
INVx1_ASAP7_75t_L g473 ( .A(n_445), .Y(n_473) );
NOR2x1_ASAP7_75t_SL g477 ( .A(n_445), .B(n_478), .Y(n_477) );
NAND4xp75_ASAP7_75t_L g445 ( .A(n_446), .B(n_452), .C(n_458), .D(n_466), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_455), .Y(n_773) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_462), .Y(n_458) );
INVxp67_ASAP7_75t_L g807 ( .A(n_460), .Y(n_807) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g555 ( .A(n_464), .Y(n_555) );
BUFx6f_ASAP7_75t_SL g760 ( .A(n_465), .Y(n_760) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g862 ( .A(n_468), .Y(n_862) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx4_ASAP7_75t_L g537 ( .A(n_479), .Y(n_537) );
OA22x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_512), .B2(n_535), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_SL g511 ( .A(n_482), .Y(n_511) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_499), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_485), .B(n_488), .C(n_492), .D(n_496), .Y(n_484) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_SL g741 ( .A(n_491), .Y(n_741) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .C(n_506), .D(n_508), .Y(n_499) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g720 ( .A(n_502), .Y(n_720) );
INVx1_ASAP7_75t_L g624 ( .A(n_507), .Y(n_624) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g535 ( .A(n_512), .Y(n_535) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
XNOR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_534), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .C(n_521), .D(n_522), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .C(n_529), .D(n_531), .Y(n_523) );
INVx1_ASAP7_75t_L g945 ( .A(n_530), .Y(n_945) );
INVx1_ASAP7_75t_L g729 ( .A(n_538), .Y(n_729) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_539), .A2(n_660), .B1(n_726), .B2(n_727), .Y(n_538) );
INVx1_ASAP7_75t_L g726 ( .A(n_539), .Y(n_726) );
AO22x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_574), .B1(n_657), .B2(n_658), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g659 ( .A(n_541), .Y(n_659) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_560), .Y(n_543) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_548), .B(n_549), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_550), .Y(n_694) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g743 ( .A(n_552), .Y(n_743) );
INVx2_ASAP7_75t_L g783 ( .A(n_552), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_563), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g718 ( .A(n_572), .Y(n_718) );
INVx2_ASAP7_75t_L g657 ( .A(n_574), .Y(n_657) );
OA22x2_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_616), .B2(n_656), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AO22x2_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_599), .B1(n_600), .B2(n_615), .Y(n_576) );
INVx1_ASAP7_75t_L g615 ( .A(n_577), .Y(n_615) );
INVx1_ASAP7_75t_L g597 ( .A(n_578), .Y(n_597) );
NAND2x1_ASAP7_75t_SL g578 ( .A(n_579), .B(n_587), .Y(n_578) );
NOR2xp67_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
INVxp67_ASAP7_75t_L g809 ( .A(n_584), .Y(n_809) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_593), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
AO22x2_ASAP7_75t_L g662 ( .A1(n_599), .A2(n_600), .B1(n_663), .B2(n_685), .Y(n_662) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
XOR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_614), .Y(n_600) );
NAND2x1_ASAP7_75t_L g601 ( .A(n_602), .B(n_607), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g656 ( .A(n_616), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_631), .C(n_639), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_625), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g714 ( .A(n_633), .Y(n_714) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_648), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_644), .C1(n_645), .C2(n_647), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_642), .A2(n_692), .B1(n_693), .B2(n_695), .C(n_696), .Y(n_691) );
INVx2_ASAP7_75t_L g697 ( .A(n_643), .Y(n_697) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_652), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_801) );
INVx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g727 ( .A(n_660), .Y(n_727) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22x1_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_686), .B1(n_687), .B2(n_725), .Y(n_661) );
INVx2_ASAP7_75t_L g725 ( .A(n_662), .Y(n_725) );
INVx2_ASAP7_75t_L g685 ( .A(n_663), .Y(n_685) );
NAND2x1_ASAP7_75t_SL g664 ( .A(n_665), .B(n_675), .Y(n_664) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_670), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B(n_669), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_681), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_678), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
XNOR2x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_724), .Y(n_688) );
NAND4xp75_ASAP7_75t_L g689 ( .A(n_690), .B(n_698), .C(n_710), .D(n_721), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_704), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_715), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AOI22xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_839), .B1(n_840), .B2(n_911), .Y(n_730) );
INVx1_ASAP7_75t_L g911 ( .A(n_731), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_775), .B2(n_838), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_752), .B1(n_753), .B2(n_774), .Y(n_733) );
INVx3_ASAP7_75t_L g774 ( .A(n_734), .Y(n_774) );
INVx5_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR2x1_ASAP7_75t_L g736 ( .A(n_737), .B(n_745), .Y(n_736) );
NAND4xp25_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .C(n_740), .D(n_744), .Y(n_737) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .C(n_750), .D(n_751), .Y(n_745) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
XNOR2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_766), .Y(n_755) );
NAND4xp25_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .C(n_761), .D(n_763), .Y(n_756) );
NAND4xp25_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .C(n_770), .D(n_772), .Y(n_766) );
INVx1_ASAP7_75t_L g838 ( .A(n_775), .Y(n_838) );
OA22x2_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_820), .B2(n_821), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AO22x2_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_794), .B2(n_819), .Y(n_777) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
OR2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_787), .Y(n_780) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .C(n_785), .D(n_786), .Y(n_781) );
BUFx2_ASAP7_75t_L g834 ( .A(n_783), .Y(n_834) );
NAND4xp25_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .C(n_790), .D(n_792), .Y(n_787) );
INVx2_ASAP7_75t_L g819 ( .A(n_794), .Y(n_819) );
INVx1_ASAP7_75t_L g818 ( .A(n_796), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_810), .Y(n_796) );
NOR3xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .C(n_805), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g798 ( .A(n_799), .B(n_800), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
XNOR2x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_837), .Y(n_821) );
NOR2xp67_ASAP7_75t_L g822 ( .A(n_823), .B(n_830), .Y(n_822) );
NAND4xp25_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .C(n_826), .D(n_827), .Y(n_823) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND4xp25_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .C(n_835), .D(n_836), .Y(n_830) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_855), .B1(n_856), .B2(n_910), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_842), .Y(n_910) );
XNOR2x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
NOR2x1_ASAP7_75t_L g844 ( .A(n_845), .B(n_850), .Y(n_844) );
NAND4xp25_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .C(n_848), .D(n_849), .Y(n_845) );
NAND4xp25_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .C(n_853), .D(n_854), .Y(n_850) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AO22x2_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_891), .B1(n_892), .B2(n_909), .Y(n_856) );
INVx2_ASAP7_75t_L g909 ( .A(n_857), .Y(n_909) );
XOR2x1_ASAP7_75t_SL g857 ( .A(n_858), .B(n_875), .Y(n_857) );
NAND2xp5_ASAP7_75t_SL g859 ( .A(n_860), .B(n_868), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_865), .Y(n_860) );
OAI21xp5_ASAP7_75t_SL g861 ( .A1(n_862), .A2(n_863), .B(n_864), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
XNOR2x1_ASAP7_75t_L g875 ( .A(n_876), .B(n_890), .Y(n_875) );
OR2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_883), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .C(n_881), .D(n_882), .Y(n_877) );
NAND4xp25_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .C(n_888), .D(n_889), .Y(n_883) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
XOR2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_908), .Y(n_892) );
NAND2x1_ASAP7_75t_L g893 ( .A(n_894), .B(n_901), .Y(n_893) );
NOR2x1_ASAP7_75t_L g894 ( .A(n_895), .B(n_898), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
NOR2x1_ASAP7_75t_L g901 ( .A(n_902), .B(n_905), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_914), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_918), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_915), .B(n_919), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g928 ( .A(n_917), .Y(n_928) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_932), .B(n_933), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
BUFx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AND2x2_ASAP7_75t_SL g926 ( .A(n_927), .B(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OR2x2_ASAP7_75t_L g976 ( .A(n_928), .B(n_929), .Y(n_976) );
OA222x2_ASAP7_75t_SL g933 ( .A1(n_934), .A2(n_952), .B1(n_954), .B2(n_972), .C1(n_973), .C2(n_976), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_935), .Y(n_951) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NOR2x1_ASAP7_75t_L g936 ( .A(n_937), .B(n_942), .Y(n_936) );
NAND4xp25_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .C(n_940), .D(n_941), .Y(n_937) );
NAND4xp25_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .C(n_948), .D(n_949), .Y(n_942) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_SL g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx3_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
XOR2x2_ASAP7_75t_L g956 ( .A(n_957), .B(n_972), .Y(n_956) );
NAND4xp75_ASAP7_75t_L g957 ( .A(n_958), .B(n_963), .C(n_967), .D(n_970), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
AND2x2_ASAP7_75t_L g963 ( .A(n_964), .B(n_966), .Y(n_963) );
AND2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
INVx1_ASAP7_75t_SL g973 ( .A(n_974), .Y(n_973) );
CKINVDCx6p67_ASAP7_75t_R g974 ( .A(n_975), .Y(n_974) );
endmodule