module fake_jpeg_26233_n_49 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_49);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_11),
.B1(n_18),
.B2(n_4),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_9),
.B1(n_14),
.B2(n_15),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_2),
.B(n_3),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_12),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.C(n_37),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

OR2x4_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_6),
.Y(n_36)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_40),
.B(n_38),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_46),
.C(n_42),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_34),
.Y(n_49)
);


endmodule