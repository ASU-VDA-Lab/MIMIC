module real_jpeg_12070_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_331, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_331;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_68),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_4),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_120),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_120),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_57),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_253)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_10),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_30),
.C(n_45),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_76),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_10),
.A2(n_111),
.B(n_164),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_10),
.A2(n_59),
.B(n_75),
.C(n_191),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_10),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_10),
.B(n_54),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_11),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_160),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_160),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_160),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_12),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_61),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g249 ( 
.A(n_13),
.B(n_60),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_14),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_14),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_14),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_324)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_16),
.A2(n_54),
.B1(n_55),
.B2(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_16),
.A2(n_40),
.B1(n_42),
.B2(n_78),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_78),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_321),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_308),
.B(n_320),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_136),
.B(n_305),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_123),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_98),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_22),
.B(n_98),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_22),
.Y(n_330)
);

FAx1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_69),
.CI(n_84),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_69),
.C(n_84),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_52),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_24),
.A2(n_25),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_26),
.A2(n_27),
.B1(n_52),
.B2(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_28),
.A2(n_32),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_28),
.B(n_165),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_28),
.A2(n_32),
.B1(n_110),
.B2(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_29),
.B(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_32),
.B(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_34),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_51),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_43),
.B1(n_51),
.B2(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_42),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_40),
.B(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_42),
.A2(n_74),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_51),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_43),
.B(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_43),
.A2(n_51),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_43),
.A2(n_51),
.B1(n_115),
.B2(n_242),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_49),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_47),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_47),
.B(n_148),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_47),
.A2(n_161),
.B(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B(n_62),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_58),
.B1(n_64),
.B2(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_55),
.A2(n_64),
.B(n_148),
.C(n_235),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g248 ( 
.A1(n_55),
.A2(n_59),
.A3(n_61),
.B1(n_236),
.B2(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_67),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_58),
.A2(n_64),
.B1(n_96),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_58),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_58),
.A2(n_62),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_58),
.A2(n_64),
.B1(n_119),
.B2(n_263),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_63),
.A2(n_216),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_63),
.A2(n_216),
.B1(n_315),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_119),
.B(n_121),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_70),
.B(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_81),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_77),
.B1(n_79),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_79),
.B1(n_89),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_71),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_71),
.A2(n_79),
.B1(n_211),
.B2(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_71),
.A2(n_197),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_76),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_72),
.B(n_198),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_72),
.A2(n_76),
.B(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_76),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_79),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_79),
.A2(n_117),
.B(n_212),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_82),
.A2(n_147),
.B(n_149),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_82),
.A2(n_149),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_86),
.B(n_91),
.C(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_91),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_91),
.B(n_128),
.C(n_132),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_95),
.B(n_127),
.C(n_134),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_105),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_104),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_105),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.C(n_118),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_106),
.A2(n_107),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_108),
.A2(n_113),
.B1(n_114),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_108),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_111),
.A2(n_112),
.B1(n_193),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_111),
.A2(n_112),
.B1(n_219),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_112),
.A2(n_170),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_148),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_112),
.A2(n_178),
.B(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_116),
.B(n_118),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_122),
.B(n_234),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_123),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_135),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_124),
.B(n_135),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_129),
.Y(n_314)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_133),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_299),
.B(n_304),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_287),
.B(n_298),
.Y(n_137)
);

OAI321xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_255),
.A3(n_280),
.B1(n_285),
.B2(n_286),
.C(n_331),
.Y(n_138)
);

AOI21x1_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_228),
.B(n_254),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_205),
.B(n_227),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_186),
.B(n_204),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_166),
.B(n_185),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_151),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_146),
.B1(n_151),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_158),
.C(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_163),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_174),
.B(n_184),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_172),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_199),
.C(n_203),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_192),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_207),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_220),
.B2(n_221),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_223),
.C(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_214),
.C(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_244),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_245),
.C(n_246),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_237),
.B2(n_243),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_238),
.C(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.C(n_269),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_258),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_264),
.C(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_266),
.B(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_279),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_274),
.C(n_279),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_297),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_319),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_318),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_313),
.B1(n_316),
.B2(n_317),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_311),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_316),
.C(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_323),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_325),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);


endmodule