module real_jpeg_6895_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_1),
.B(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_1),
.A2(n_203),
.B(n_252),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_1),
.B(n_180),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_1),
.B(n_362),
.C(n_365),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_1),
.A2(n_76),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_1),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_1),
.B(n_136),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_1),
.A2(n_25),
.B1(n_405),
.B2(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_35),
.B1(n_38),
.B2(n_43),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_43),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_2),
.A2(n_43),
.B1(n_76),
.B2(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_2),
.A2(n_43),
.B1(n_139),
.B2(n_222),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_3),
.A2(n_119),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_3),
.A2(n_119),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_119),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_5),
.A2(n_101),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_5),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_5),
.A2(n_185),
.B1(n_247),
.B2(n_284),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_5),
.A2(n_284),
.B1(n_380),
.B2(n_382),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_5),
.A2(n_284),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_6),
.A2(n_75),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_6),
.A2(n_26),
.B1(n_75),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_75),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_7),
.A2(n_47),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_47),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_7),
.A2(n_47),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_8),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_8),
.Y(n_300)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_10),
.Y(n_250)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_12),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_12),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_12),
.A2(n_141),
.B1(n_177),
.B2(n_274),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_12),
.A2(n_27),
.B1(n_177),
.B2(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_12),
.A2(n_52),
.B1(n_177),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_13),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_14),
.A2(n_101),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_14),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_14),
.A2(n_121),
.B1(n_281),
.B2(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_14),
.A2(n_52),
.B1(n_281),
.B2(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_14),
.A2(n_281),
.B1(n_406),
.B2(n_408),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_15),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_488),
.C(n_492),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_486),
.B(n_490),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_476),
.B(n_485),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_209),
.A3(n_232),
.B(n_473),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_188),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_21),
.B(n_188),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_111),
.C(n_151),
.Y(n_21)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_22),
.B(n_111),
.CI(n_151),
.CON(n_350),
.SN(n_350)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_77),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_23),
.A2(n_24),
.B(n_79),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_24),
.A2(n_78),
.B1(n_79),
.B2(n_110),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_24),
.A2(n_44),
.B1(n_78),
.B2(n_342),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_25),
.B(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_25),
.A2(n_255),
.B1(n_261),
.B2(n_265),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_25),
.A2(n_265),
.B(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_25),
.A2(n_160),
.B(n_387),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_25),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_25),
.A2(n_299),
.B1(n_393),
.B2(n_405),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_25),
.A2(n_34),
.B(n_297),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_26),
.Y(n_257)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_29),
.Y(n_270)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_31),
.Y(n_325)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_31),
.Y(n_417)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_34),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_37),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_41),
.Y(n_407)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_42),
.Y(n_260)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_42),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_44),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_55),
.B(n_70),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_46),
.A2(n_56),
.B1(n_71),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_49),
.A2(n_124),
.B1(n_125),
.B2(n_128),
.Y(n_123)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_50),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_50),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_50),
.Y(n_381)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_51),
.Y(n_147)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_55),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_55),
.A2(n_144),
.B(n_145),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_55),
.A2(n_70),
.B(n_145),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_55),
.A2(n_144),
.B1(n_149),
.B2(n_167),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_55),
.A2(n_457),
.B(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_56),
.A2(n_71),
.B1(n_367),
.B2(n_370),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_56),
.A2(n_71),
.B1(n_370),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_56),
.A2(n_71),
.B1(n_379),
.B2(n_444),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_58),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_65),
.Y(n_365)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_98),
.B(n_103),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_80),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_80),
.A2(n_180),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_80),
.A2(n_180),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_80),
.A2(n_98),
.B(n_180),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_81),
.A2(n_174),
.B(n_179),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_81),
.A2(n_109),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_81),
.A2(n_109),
.B1(n_174),
.B2(n_283),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_81),
.A2(n_482),
.B(n_483),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_91)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_93),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_93),
.Y(n_442)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_94),
.Y(n_277)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_94),
.Y(n_333)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_96),
.Y(n_434)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_97),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_98),
.B(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_100),
.Y(n_285)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_103),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_107),
.Y(n_231)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_109),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_109),
.A2(n_199),
.B(n_205),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_142),
.B(n_150),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_142),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_122),
.B1(n_136),
.B2(n_137),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_114),
.A2(n_123),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_122),
.B(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_122),
.A2(n_137),
.B(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_122),
.A2(n_220),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_122),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_122),
.A2(n_136),
.B1(n_330),
.B2(n_441),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_122),
.A2(n_136),
.B(n_480),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_123),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_123),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_123),
.A2(n_292),
.B1(n_293),
.B2(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_124),
.Y(n_369)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_125),
.Y(n_436)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_127),
.Y(n_430)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_184),
.Y(n_195)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g425 ( 
.A1(n_141),
.A2(n_426),
.A3(n_428),
.B1(n_431),
.B2(n_435),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_143),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_144),
.B(n_368),
.Y(n_403)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_146),
.Y(n_437)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_189),
.CI(n_208),
.CON(n_188),
.SN(n_188)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_172),
.C(n_181),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_152),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_164),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_153),
.A2(n_164),
.B1(n_165),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_153),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_155),
.A2(n_256),
.B(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_156),
.Y(n_301)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_162),
.Y(n_413)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_168),
.Y(n_445)
);

INVx5_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_172),
.A2(n_173),
.B1(n_181),
.B2(n_182),
.Y(n_344)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_179),
.B(n_205),
.Y(n_488)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_188),
.B(n_211),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_198),
.B2(n_207),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_197),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_192),
.B(n_217),
.C(n_225),
.Y(n_484)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_197),
.C(n_198),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_195),
.A2(n_221),
.B(n_293),
.Y(n_311)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_207),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_198),
.B(n_212),
.C(n_215),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_210),
.A2(n_474),
.B(n_475),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_225),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_221),
.Y(n_480)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_227),
.Y(n_482)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_351),
.B(n_467),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_336),
.C(n_348),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_315),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_235),
.A2(n_469),
.B(n_470),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_303),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_236),
.B(n_303),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_286),
.C(n_295),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_237),
.B(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_271),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_238),
.B(n_272),
.C(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_254),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_239),
.B(n_254),
.Y(n_318)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_243),
.A3(n_244),
.B1(n_246),
.B2(n_251),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_259),
.Y(n_388)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_268),
.Y(n_394)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_269),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_295),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.C(n_291),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_287),
.B(n_288),
.CI(n_291),
.CON(n_317),
.SN(n_317)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx3_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_300),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_313),
.C(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_334),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_316),
.B(n_334),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.C(n_319),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_317),
.B(n_465),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_317),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_318),
.B(n_319),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_326),
.C(n_328),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_320),
.A2(n_321),
.B1(n_326),
.B2(n_327),
.Y(n_452)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_328),
.B(n_452),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g467 ( 
.A1(n_336),
.A2(n_348),
.B(n_468),
.C(n_471),
.D(n_472),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_347),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_337),
.B(n_347),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_341),
.C(n_346),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_349),
.B(n_350),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_350),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_462),
.B(n_466),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_447),
.B(n_461),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_421),
.B(n_446),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_389),
.B(n_420),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_374),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_374),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_366),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_366),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_368),
.B(n_432),
.Y(n_431)
);

OAI21xp33_ASAP7_75t_SL g441 ( 
.A1(n_368),
.A2(n_431),
.B(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_386),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_385),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_376),
.B(n_385),
.C(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_378),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_401),
.B(n_419),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_400),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_400),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_396),
.B1(n_397),
.B2(n_398),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_394),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_411),
.B(n_418),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_403),
.B(n_404),
.Y(n_418)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_423),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_439),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_440),
.C(n_443),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_438),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_444),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_448),
.B(n_449),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_450),
.A2(n_451),
.B1(n_453),
.B2(n_454),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_456),
.C(n_459),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_459),
.B2(n_460),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_463),
.B(n_464),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_478),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_478),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_478),
.B(n_488),
.Y(n_491)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_481),
.CI(n_484),
.CON(n_478),
.SN(n_478)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_488),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);


endmodule