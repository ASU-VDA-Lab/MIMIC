module fake_jpeg_21528_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_2),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_54),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_44),
.B1(n_43),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_52),
.B1(n_50),
.B2(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_59),
.B1(n_51),
.B2(n_55),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_89),
.B1(n_92),
.B2(n_41),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_43),
.B(n_53),
.C(n_47),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_88),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_62),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_45),
.B1(n_56),
.B2(n_49),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_93),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_10),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_103),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_40),
.B1(n_3),
.B2(n_5),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_35),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_4),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_12),
.C(n_13),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_113),
.C(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_109),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_23),
.B1(n_27),
.B2(n_30),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_32),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_111),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_96),
.C(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_100),
.B(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_122),
.Y(n_123)
);

BUFx4f_ASAP7_75t_SL g124 ( 
.A(n_123),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_114),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_111),
.C(n_120),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_128),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_118),
.Y(n_130)
);


endmodule