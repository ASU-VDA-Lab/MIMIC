module fake_netlist_1_5748_n_624 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_624);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_624;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_178;
wire n_616;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_521;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g177 ( .A(n_7), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_31), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_88), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_174), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
NOR2xp67_ASAP7_75t_L g182 ( .A(n_108), .B(n_138), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_34), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_50), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_141), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_130), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_41), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_126), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_37), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_46), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_8), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_86), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_43), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_142), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_102), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_40), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_66), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_161), .Y(n_200) );
INVx1_ASAP7_75t_SL g201 ( .A(n_98), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_143), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_27), .B(n_33), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_124), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_65), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_120), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_131), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_25), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_95), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_9), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_91), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_73), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_1), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_57), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_3), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_42), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_160), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_122), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_112), .Y(n_221) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_39), .B(n_12), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_48), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_149), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_117), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_96), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_94), .B(n_109), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_111), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_90), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_60), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_5), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_146), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g234 ( .A(n_152), .B(n_147), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_5), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_76), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_157), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_103), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_148), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_129), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_164), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_118), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_97), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_140), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_84), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_0), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_99), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_150), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_116), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_137), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_9), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_170), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_135), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_11), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_89), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_101), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_113), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_169), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_156), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_159), .Y(n_261) );
INVxp33_ASAP7_75t_SL g262 ( .A(n_22), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_132), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_110), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_145), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_72), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_153), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_173), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_154), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_59), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_81), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_83), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_68), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_53), .Y(n_275) );
INVxp33_ASAP7_75t_L g276 ( .A(n_100), .Y(n_276) );
NOR2xp67_ASAP7_75t_L g277 ( .A(n_166), .B(n_1), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_38), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_144), .Y(n_279) );
INVxp33_ASAP7_75t_SL g280 ( .A(n_236), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_188), .A2(n_92), .B(n_172), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_199), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_199), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_236), .B(n_0), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_270), .B(n_2), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_270), .Y(n_288) );
OAI22xp5_ASAP7_75t_SL g289 ( .A1(n_232), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_289) );
OAI22x1_ASAP7_75t_SL g290 ( .A1(n_192), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_178), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_207), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_207), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_247), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_223), .B(n_6), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_189), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_177), .B(n_8), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
INVx5_ASAP7_75t_L g299 ( .A(n_223), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_288), .B(n_187), .Y(n_300) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_288), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_292), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_283), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_280), .B(n_218), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_296), .B(n_198), .Y(n_306) );
BUFx4f_ASAP7_75t_L g307 ( .A(n_292), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_293), .B(n_276), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_291), .B(n_211), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_293), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_286), .B(n_214), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_310), .B(n_284), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_301), .B(n_297), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_302), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_302), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_311), .B(n_294), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_301), .B(n_297), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_312), .B(n_298), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_309), .B(n_196), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_306), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_309), .A2(n_281), .B(n_235), .C(n_252), .Y(n_323) );
BUFx2_ASAP7_75t_SL g324 ( .A(n_321), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_314), .A2(n_300), .B(n_305), .C(n_306), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_314), .B(n_319), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_320), .A2(n_308), .B(n_216), .Y(n_327) );
NAND3x1_ASAP7_75t_L g328 ( .A(n_321), .B(n_289), .C(n_290), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_315), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_323), .A2(n_307), .B(n_308), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_313), .A2(n_295), .B(n_262), .C(n_180), .Y(n_331) );
OAI22xp5_ASAP7_75t_SL g332 ( .A1(n_317), .A2(n_289), .B1(n_237), .B2(n_239), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_322), .A2(n_307), .B(n_181), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_316), .B(n_202), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_316), .A2(n_210), .B1(n_224), .B2(n_228), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_326), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_329), .Y(n_337) );
AO31x2_ASAP7_75t_L g338 ( .A1(n_330), .A2(n_240), .A3(n_183), .B(n_184), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_333), .A2(n_318), .B(n_186), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_335), .B(n_242), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_325), .A2(n_194), .B(n_179), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_324), .B(n_257), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_331), .A2(n_204), .B(n_197), .Y(n_343) );
OAI22x1_ASAP7_75t_L g344 ( .A1(n_332), .A2(n_244), .B1(n_241), .B2(n_201), .Y(n_344) );
AO32x2_ASAP7_75t_L g345 ( .A1(n_335), .A2(n_327), .A3(n_277), .B1(n_283), .B2(n_287), .Y(n_345) );
OAI22x1_ASAP7_75t_L g346 ( .A1(n_334), .A2(n_244), .B1(n_201), .B2(n_241), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_SL g347 ( .A1(n_328), .A2(n_243), .B(n_279), .C(n_278), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_329), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_208), .B(n_205), .Y(n_349) );
BUFx8_ASAP7_75t_SL g350 ( .A(n_326), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_326), .B(n_259), .Y(n_351) );
BUFx4_ASAP7_75t_SL g352 ( .A(n_324), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_326), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_353), .B(n_10), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_350), .A2(n_261), .B1(n_230), .B2(n_231), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_352), .B(n_245), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_336), .A2(n_182), .B(n_234), .C(n_222), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_336), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_349), .A2(n_209), .B(n_206), .Y(n_359) );
INVx4_ASAP7_75t_SL g360 ( .A(n_340), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
AO31x2_ASAP7_75t_L g362 ( .A1(n_346), .A2(n_256), .A3(n_213), .B(n_215), .Y(n_362) );
BUFx10_ASAP7_75t_L g363 ( .A(n_342), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_348), .B(n_217), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_341), .A2(n_220), .B(n_219), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_339), .A2(n_225), .B(n_221), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_351), .B(n_10), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_343), .A2(n_273), .B(n_233), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_344), .B(n_226), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_338), .B(n_238), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_347), .B(n_246), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_255), .B(n_250), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_345), .A2(n_266), .B1(n_268), .B2(n_258), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g376 ( .A1(n_345), .A2(n_260), .B(n_267), .C(n_265), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_338), .B(n_272), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_338), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_353), .Y(n_379) );
AOI21x1_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_275), .B(n_303), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_336), .A2(n_249), .B1(n_263), .B2(n_269), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_353), .B(n_185), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_336), .A2(n_227), .B(n_203), .Y(n_384) );
AOI21x1_ASAP7_75t_L g385 ( .A1(n_349), .A2(n_303), .B(n_287), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_253), .B1(n_193), .B2(n_195), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_353), .B(n_191), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_336), .A2(n_299), .B(n_282), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_376), .A2(n_287), .B(n_285), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
AO21x2_ASAP7_75t_L g393 ( .A1(n_375), .A2(n_285), .B(n_283), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_360), .B(n_13), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_388), .Y(n_396) );
BUFx12f_ASAP7_75t_L g397 ( .A(n_388), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_360), .B(n_200), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_374), .A2(n_285), .B(n_299), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
INVx4_ASAP7_75t_L g402 ( .A(n_356), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_364), .B(n_212), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_382), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_369), .B(n_229), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_377), .A2(n_299), .B(n_282), .Y(n_410) );
AOI21xp5_ASAP7_75t_SL g411 ( .A1(n_372), .A2(n_271), .B(n_264), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_368), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_383), .B(n_248), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
OR2x6_ASAP7_75t_L g417 ( .A(n_387), .B(n_14), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_355), .B(n_251), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_363), .B(n_254), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_367), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_367), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_389), .B(n_274), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_381), .B(n_15), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_370), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_359), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_373), .Y(n_426) );
NAND2xp33_ASAP7_75t_L g427 ( .A(n_386), .B(n_16), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_365), .A2(n_17), .B(n_18), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_380), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_384), .B(n_19), .Y(n_430) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_385), .A2(n_20), .B(n_21), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_390), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_385), .A2(n_23), .B(n_24), .Y(n_434) );
OA21x2_ASAP7_75t_L g435 ( .A1(n_357), .A2(n_26), .B(n_28), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_368), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_364), .B(n_175), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_358), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_358), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_358), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_360), .A2(n_29), .B1(n_30), .B2(n_32), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_358), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_358), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_379), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_358), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_364), .B(n_171), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_358), .B(n_35), .Y(n_447) );
OAI21x1_ASAP7_75t_L g448 ( .A1(n_385), .A2(n_36), .B(n_44), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_394), .Y(n_449) );
NAND4xp25_ASAP7_75t_SL g450 ( .A(n_411), .B(n_45), .C(n_47), .D(n_49), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_438), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_402), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_439), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_444), .B(n_51), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_392), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_392), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_168), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_440), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_442), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_401), .B(n_52), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_416), .B(n_54), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_443), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_445), .B(n_55), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_412), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_412), .B(n_56), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_407), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_437), .A2(n_58), .B1(n_61), .B2(n_62), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_436), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_436), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_414), .B(n_63), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_394), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_414), .B(n_64), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_447), .B(n_67), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_405), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_409), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_446), .B(n_69), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_406), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_403), .B(n_167), .C(n_71), .D(n_74), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_421), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_426), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_399), .B(n_70), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_404), .B(n_75), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_396), .B(n_77), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_397), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_418), .B(n_78), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_432), .B(n_79), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_421), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_429), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_430), .B(n_80), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_410), .B(n_82), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_433), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_430), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_410), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_489), .B(n_393), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_451), .B(n_423), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_462), .B(n_393), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_453), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_466), .B(n_461), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_471), .B(n_391), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_457), .B(n_424), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_472), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_496), .B(n_424), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_477), .B(n_391), .Y(n_517) );
AND2x4_ASAP7_75t_SL g518 ( .A(n_469), .B(n_441), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_474), .B(n_400), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_497), .B(n_503), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_459), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_475), .B(n_400), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_454), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_480), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_469), .B(n_435), .C(n_427), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_481), .B(n_425), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_460), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_482), .Y(n_530) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_487), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_468), .B(n_435), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_488), .B(n_425), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_468), .B(n_434), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_488), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_468), .B(n_434), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_449), .B(n_431), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_449), .B(n_431), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_465), .B(n_419), .Y(n_540) );
NOR2xp67_ASAP7_75t_SL g541 ( .A(n_486), .B(n_428), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_499), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_483), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_519), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_529), .B(n_483), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_508), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_544), .B(n_502), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_509), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_510), .B(n_502), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_538), .B(n_504), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_543), .B(n_495), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_516), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_522), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_525), .Y(n_557) );
NAND2x1_ASAP7_75t_L g558 ( .A(n_543), .B(n_495), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_527), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_515), .B(n_476), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_505), .B(n_452), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_531), .B(n_485), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_531), .B(n_493), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_513), .B(n_455), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_535), .B(n_458), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_530), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_540), .Y(n_567) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_524), .B(n_492), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_535), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_521), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_548), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_551), .B(n_521), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_555), .A2(n_526), .B(n_486), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_554), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_559), .B(n_517), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_557), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_566), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g578 ( .A1(n_563), .A2(n_473), .B(n_494), .C(n_491), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_547), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_561), .A2(n_518), .B1(n_541), .B2(n_567), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_559), .B(n_533), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_553), .B(n_520), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_558), .A2(n_450), .B(n_533), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_570), .B(n_511), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_546), .B(n_523), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_553), .A2(n_518), .B1(n_479), .B2(n_494), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_584), .B(n_572), .Y(n_587) );
AO22x2_ASAP7_75t_L g588 ( .A1(n_574), .A2(n_562), .B1(n_550), .B2(n_545), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_586), .A2(n_568), .B1(n_565), .B2(n_569), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_573), .A2(n_549), .B(n_560), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_582), .A2(n_564), .B1(n_560), .B2(n_479), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_580), .A2(n_506), .B1(n_549), .B2(n_484), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_581), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g594 ( .A1(n_578), .A2(n_450), .B(n_473), .C(n_552), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_575), .B(n_537), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_571), .Y(n_596) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_592), .A2(n_583), .B(n_582), .C(n_585), .Y(n_597) );
NOR3x1_ASAP7_75t_L g598 ( .A(n_589), .B(n_579), .C(n_577), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_590), .B(n_576), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_593), .B(n_476), .Y(n_600) );
OAI322xp33_ASAP7_75t_L g601 ( .A1(n_587), .A2(n_552), .A3(n_512), .B1(n_514), .B2(n_556), .C1(n_500), .C2(n_478), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g602 ( .A1(n_591), .A2(n_539), .A3(n_507), .B1(n_490), .B2(n_514), .C1(n_500), .C2(n_542), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_594), .A2(n_470), .B(n_463), .C(n_464), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_596), .A2(n_413), .B(n_408), .C(n_501), .Y(n_604) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_588), .B(n_532), .C(n_536), .D(n_534), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_588), .A2(n_542), .B1(n_528), .B2(n_522), .C(n_467), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_599), .B(n_606), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_598), .Y(n_608) );
NAND3xp33_ASAP7_75t_SL g609 ( .A(n_597), .B(n_603), .C(n_604), .Y(n_609) );
AND4x1_ASAP7_75t_L g610 ( .A(n_608), .B(n_605), .C(n_595), .D(n_602), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_609), .B(n_601), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_611), .Y(n_612) );
XNOR2xp5_ASAP7_75t_L g613 ( .A(n_610), .B(n_607), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_612), .B(n_528), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_613), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_615), .A2(n_422), .B(n_448), .C(n_600), .Y(n_616) );
AOI22x1_ASAP7_75t_L g617 ( .A1(n_614), .A2(n_85), .B1(n_87), .B2(n_93), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_616), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_617), .A2(n_104), .B(n_105), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_618), .A2(n_106), .B(n_107), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_619), .A2(n_114), .B(n_115), .Y(n_621) );
OAI222xp33_ASAP7_75t_SL g622 ( .A1(n_620), .A2(n_119), .B1(n_121), .B2(n_123), .C1(n_125), .C2(n_127), .Y(n_622) );
AO21x2_ASAP7_75t_L g623 ( .A1(n_622), .A2(n_621), .B(n_133), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_623), .A2(n_128), .B1(n_134), .B2(n_136), .Y(n_624) );
endmodule