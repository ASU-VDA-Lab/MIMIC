module fake_aes_2289_n_708 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_708);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_708;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_49), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_16), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_62), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_59), .Y(n_84) );
CKINVDCx14_ASAP7_75t_R g85 ( .A(n_72), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_68), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_45), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_41), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_9), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_56), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_12), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_39), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_16), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_42), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_23), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_54), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_46), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_1), .B(n_69), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_64), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_30), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_34), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_44), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_57), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_27), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_51), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_66), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_15), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_101), .B(n_0), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_101), .B(n_0), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_98), .B(n_3), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_98), .B(n_4), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
AND3x2_ASAP7_75t_L g138 ( .A(n_87), .B(n_5), .C(n_6), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_105), .B(n_5), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_106), .Y(n_140) );
INVxp67_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_93), .B(n_7), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_84), .A2(n_36), .B(n_76), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_91), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_97), .B(n_10), .Y(n_147) );
OR2x2_ASAP7_75t_L g148 ( .A(n_97), .B(n_11), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_126), .Y(n_149) );
INVx2_ASAP7_75t_SL g150 ( .A(n_99), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_108), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_120), .B(n_11), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_115), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_119), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_82), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_85), .B(n_12), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_89), .Y(n_164) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_89), .A2(n_40), .B(n_75), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_90), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_90), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_113), .B(n_13), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_122), .B(n_13), .Y(n_169) );
XOR2xp5_ASAP7_75t_L g170 ( .A(n_160), .B(n_100), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_130), .B(n_131), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_157), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_141), .B(n_127), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_141), .B(n_79), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_168), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_127), .B(n_124), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_132), .B(n_123), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_130), .B(n_80), .Y(n_181) );
NAND3xp33_ASAP7_75t_L g182 ( .A(n_128), .B(n_125), .C(n_82), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
OR2x2_ASAP7_75t_SL g187 ( .A(n_148), .B(n_122), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_132), .B(n_124), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_133), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_146), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_131), .B(n_113), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_135), .B(n_114), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
INVxp33_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_148), .B(n_104), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_146), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_153), .B(n_117), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_135), .B(n_111), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_166), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_137), .B(n_114), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_137), .B(n_123), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_146), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_159), .B(n_121), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_149), .Y(n_220) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_142), .B(n_121), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_159), .B(n_111), .Y(n_222) );
INVx5_ASAP7_75t_L g223 ( .A(n_146), .Y(n_223) );
INVxp33_ASAP7_75t_L g224 ( .A(n_142), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_147), .A2(n_95), .B(n_96), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g227 ( .A(n_161), .B(n_95), .C(n_96), .Y(n_227) );
INVx5_ASAP7_75t_L g228 ( .A(n_149), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_161), .B(n_92), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_163), .B(n_92), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_149), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_163), .B(n_94), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_134), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_171), .A2(n_143), .B(n_165), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_174), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_170), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_174), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_224), .B(n_175), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_198), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_203), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_224), .B(n_164), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_187), .A2(n_145), .B1(n_91), .B2(n_147), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_214), .B(n_164), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_199), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_222), .B(n_169), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_198), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_221), .B(n_169), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_208), .B(n_145), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_178), .B(n_150), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_221), .B(n_156), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_175), .B(n_156), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_179), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_177), .Y(n_257) );
OAI22xp5_ASAP7_75t_SL g258 ( .A1(n_187), .A2(n_165), .B1(n_143), .B2(n_94), .Y(n_258) );
INVx6_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_199), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_219), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_200), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_179), .B(n_219), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_180), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_177), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_173), .B(n_167), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_179), .B(n_138), .Y(n_267) );
INVx5_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_205), .Y(n_269) );
CKINVDCx11_ASAP7_75t_R g270 ( .A(n_188), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_180), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_180), .A2(n_150), .B1(n_138), .B2(n_86), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_196), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_213), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_L g275 ( .A1(n_217), .A2(n_152), .B(n_154), .C(n_158), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_183), .B(n_150), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_188), .B(n_151), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_218), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_215), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_200), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_219), .B(n_151), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_216), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_230), .B(n_151), .Y(n_284) );
INVx4_ASAP7_75t_L g285 ( .A(n_173), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
AOI211xp5_ASAP7_75t_L g287 ( .A1(n_202), .A2(n_107), .B(n_155), .C(n_151), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_211), .B(n_155), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_230), .B(n_155), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_188), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_230), .B(n_155), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_218), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_189), .B(n_167), .Y(n_295) );
INVx4_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_210), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_232), .B(n_152), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_202), .B(n_152), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_210), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_232), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_261), .B(n_211), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_273), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_242), .A2(n_182), .B(n_186), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_288), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_261), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_263), .A2(n_192), .B1(n_194), .B2(n_191), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_259), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_270), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_296), .A2(n_189), .B1(n_176), .B2(n_227), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_245), .A2(n_226), .B1(n_189), .B2(n_181), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_243), .B(n_226), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_235), .A2(n_226), .B1(n_217), .B2(n_229), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_239), .B(n_171), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_241), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_241), .Y(n_319) );
AND3x1_ASAP7_75t_SL g320 ( .A(n_244), .B(n_116), .C(n_118), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_238), .A2(n_229), .B1(n_167), .B2(n_231), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_288), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_250), .A2(n_197), .B1(n_154), .B2(n_158), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_248), .B(n_256), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_241), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_259), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_268), .B(n_197), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_255), .B(n_158), .Y(n_329) );
CKINVDCx8_ASAP7_75t_R g330 ( .A(n_237), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_257), .A2(n_165), .B1(n_143), .B2(n_102), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_299), .B(n_154), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_240), .B(n_109), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_249), .B(n_110), .Y(n_336) );
CKINVDCx11_ASAP7_75t_R g337 ( .A(n_270), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_288), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_268), .B(n_223), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_241), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_280), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_280), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_264), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_264), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_264), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_267), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_271), .Y(n_350) );
AND3x1_ASAP7_75t_SL g351 ( .A(n_237), .B(n_112), .C(n_103), .Y(n_351) );
O2A1O1Ixp5_ASAP7_75t_L g352 ( .A1(n_234), .A2(n_231), .B(n_209), .C(n_212), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_271), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_268), .B(n_207), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_306), .A2(n_301), .B1(n_290), .B2(n_253), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_315), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
BUFx12f_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_326), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_306), .A2(n_298), .B1(n_271), .B2(n_278), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_302), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_315), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_309), .A2(n_257), .B1(n_265), .B2(n_267), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_324), .B(n_246), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
NOR2xp33_ASAP7_75t_SL g367 ( .A(n_330), .B(n_271), .Y(n_367) );
OAI222xp33_ASAP7_75t_L g368 ( .A1(n_309), .A2(n_265), .B1(n_251), .B2(n_272), .C1(n_262), .C2(n_247), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_349), .B(n_283), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_311), .A2(n_278), .B1(n_282), .B2(n_284), .Y(n_371) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_338), .A2(n_277), .B1(n_286), .B2(n_268), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_338), .A2(n_277), .B1(n_252), .B2(n_258), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_317), .B(n_254), .Y(n_374) );
NOR2x1p5_ASAP7_75t_L g375 ( .A(n_331), .B(n_333), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_305), .B(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_303), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_317), .B(n_291), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_311), .A2(n_276), .B1(n_281), .B2(n_260), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_336), .A2(n_259), .B1(n_252), .B2(n_293), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_322), .B(n_266), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_335), .A2(n_266), .B1(n_236), .B2(n_292), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_326), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_304), .A2(n_269), .B1(n_292), .B2(n_279), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_313), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_325), .Y(n_387) );
NOR3xp33_ASAP7_75t_L g388 ( .A(n_368), .B(n_287), .C(n_329), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_330), .B1(n_314), .B2(n_307), .C(n_312), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_375), .B(n_346), .Y(n_390) );
OAI33xp33_ASAP7_75t_L g391 ( .A1(n_379), .A2(n_323), .A3(n_334), .B1(n_310), .B2(n_346), .B3(n_351), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_332), .B(n_321), .C(n_320), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_362), .A2(n_341), .B1(n_325), .B2(n_343), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_376), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_365), .A2(n_331), .B1(n_333), .B2(n_327), .Y(n_396) );
OAI33xp33_ASAP7_75t_L g397 ( .A1(n_371), .A2(n_295), .A3(n_129), .B1(n_140), .B2(n_144), .B3(n_136), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_365), .A2(n_331), .B1(n_333), .B2(n_327), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_376), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_358), .A2(n_352), .B(n_275), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_367), .A2(n_341), .B1(n_343), .B2(n_326), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_356), .B(n_348), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_356), .B(n_348), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_374), .B(n_308), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_359), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g408 ( .A1(n_363), .A2(n_326), .B1(n_345), .B2(n_342), .C1(n_308), .C2(n_316), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_374), .A2(n_316), .B1(n_328), .B2(n_342), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_374), .A2(n_275), .B1(n_167), .B2(n_295), .C(n_328), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_378), .A2(n_316), .B1(n_328), .B2(n_345), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_378), .A2(n_328), .B1(n_236), .B2(n_269), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_389), .A2(n_381), .B(n_361), .C(n_355), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_388), .A2(n_380), .B1(n_372), .B2(n_375), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_409), .B1(n_399), .B2(n_395), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_404), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_393), .A2(n_359), .B1(n_383), .B2(n_387), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_406), .A2(n_167), .B1(n_387), .B2(n_382), .C(n_386), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_404), .Y(n_422) );
NOR2x1_ASAP7_75t_SL g423 ( .A(n_394), .B(n_357), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_394), .Y(n_424) );
OAI222xp33_ASAP7_75t_L g425 ( .A1(n_403), .A2(n_360), .B1(n_386), .B2(n_358), .C1(n_370), .C2(n_384), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_403), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_392), .A2(n_385), .B1(n_149), .B2(n_360), .C(n_231), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_384), .B1(n_370), .B2(n_347), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_402), .B(n_143), .Y(n_429) );
OAI321xp33_ASAP7_75t_L g430 ( .A1(n_396), .A2(n_129), .A3(n_144), .B1(n_140), .B2(n_136), .C(n_134), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_390), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_390), .A2(n_398), .B1(n_397), .B2(n_405), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_402), .B(n_143), .Y(n_433) );
OAI33xp33_ASAP7_75t_L g434 ( .A1(n_412), .A2(n_129), .A3(n_136), .B1(n_140), .B2(n_144), .B3(n_220), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_407), .A2(n_165), .B1(n_357), .B2(n_366), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_415), .A2(n_209), .B(n_212), .C(n_220), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_414), .B(n_14), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_410), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_411), .B(n_15), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_400), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_407), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_410), .B(n_165), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_413), .A2(n_319), .B1(n_279), .B2(n_340), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_410), .B(n_366), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_401), .Y(n_449) );
AOI21xp5_ASAP7_75t_SL g450 ( .A1(n_393), .A2(n_366), .B(n_357), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_394), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_426), .B(n_134), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_448), .A2(n_353), .B1(n_347), .B2(n_366), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_426), .B(n_366), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_451), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_419), .B(n_357), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_451), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_424), .B(n_17), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_424), .B(n_19), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_422), .B(n_184), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_419), .B(n_21), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_440), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_440), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_417), .A2(n_353), .B1(n_344), .B2(n_340), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_423), .B(n_25), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_441), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_441), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_442), .B(n_184), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_420), .A2(n_344), .B1(n_340), .B2(n_318), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_442), .B(n_172), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_446), .B(n_172), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_418), .B(n_344), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_431), .B(n_206), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_429), .B(n_433), .Y(n_478) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_444), .A2(n_206), .B(n_190), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_449), .B(n_326), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_438), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_431), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_447), .B(n_26), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_438), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_447), .B(n_28), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_425), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_429), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_437), .A2(n_350), .B1(n_318), .B2(n_228), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_433), .Y(n_489) );
OAI31xp33_ASAP7_75t_L g490 ( .A1(n_439), .A2(n_354), .A3(n_339), .B(n_185), .Y(n_490) );
OAI21x1_ASAP7_75t_L g491 ( .A1(n_450), .A2(n_185), .B(n_190), .Y(n_491) );
NAND2x1p5_ASAP7_75t_SL g492 ( .A(n_444), .B(n_204), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_450), .B(n_350), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_416), .B(n_228), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_29), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_428), .B(n_204), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_421), .A2(n_350), .B1(n_318), .B2(n_354), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_209), .Y(n_499) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_430), .A2(n_300), .B(n_297), .Y(n_500) );
OAI33xp33_ASAP7_75t_L g501 ( .A1(n_436), .A2(n_300), .A3(n_32), .B1(n_33), .B2(n_38), .B3(n_43), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_427), .B(n_228), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_455), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_462), .B(n_445), .Y(n_504) );
NOR2xp33_ASAP7_75t_SL g505 ( .A(n_486), .B(n_434), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_455), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_478), .B(n_228), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_486), .B(n_350), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_462), .B(n_31), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_478), .B(n_228), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_494), .A2(n_223), .B1(n_207), .B2(n_201), .C(n_195), .Y(n_511) );
AOI322xp5_ASAP7_75t_L g512 ( .A1(n_457), .A2(n_339), .A3(n_354), .B1(n_53), .B2(n_55), .C1(n_60), .C2(n_61), .Y(n_512) );
NAND2xp33_ASAP7_75t_L g513 ( .A(n_496), .B(n_350), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_464), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_478), .B(n_47), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_489), .B(n_50), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_489), .B(n_63), .Y(n_518) );
NOR2x1p5_ASAP7_75t_L g519 ( .A(n_486), .B(n_354), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_486), .A2(n_339), .B1(n_223), .B2(n_207), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_452), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_487), .B(n_65), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_482), .B(n_67), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_487), .B(n_71), .Y(n_524) );
OA211x2_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_73), .B(n_77), .C(n_223), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_494), .B(n_193), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_452), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_495), .A2(n_339), .B(n_207), .Y(n_528) );
INVxp67_ASAP7_75t_SL g529 ( .A(n_477), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_482), .B(n_233), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_477), .B(n_233), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_495), .A2(n_207), .B(n_223), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_452), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_477), .B(n_233), .Y(n_534) );
OAI33xp33_ASAP7_75t_L g535 ( .A1(n_499), .A2(n_193), .A3(n_195), .B1(n_201), .B2(n_233), .B3(n_475), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_463), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_454), .B(n_233), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_454), .B(n_201), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_475), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g540 ( .A1(n_496), .A2(n_193), .B(n_195), .C(n_201), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_454), .B(n_193), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_463), .B(n_195), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_464), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_456), .B(n_483), .Y(n_544) );
OR2x6_ASAP7_75t_L g545 ( .A(n_493), .B(n_491), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_456), .B(n_483), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_456), .B(n_485), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_484), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_499), .B(n_490), .C(n_465), .Y(n_550) );
OAI31xp33_ASAP7_75t_L g551 ( .A1(n_498), .A2(n_466), .A3(n_485), .B(n_480), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_469), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_492), .B(n_484), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_464), .B(n_467), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_492), .B(n_481), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_467), .B(n_481), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_468), .B(n_467), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_468), .B(n_479), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_468), .B(n_479), .Y(n_559) );
BUFx3_ASAP7_75t_L g560 ( .A(n_468), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_458), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_554), .B(n_479), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_520), .B(n_466), .C(n_474), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_503), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_506), .Y(n_565) );
AND2x2_ASAP7_75t_SL g566 ( .A(n_513), .B(n_458), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_539), .B(n_550), .Y(n_567) );
OA211x2_ASAP7_75t_L g568 ( .A1(n_551), .A2(n_471), .B(n_453), .C(n_474), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_529), .B(n_492), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_515), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_520), .A2(n_488), .B1(n_460), .B2(n_476), .C(n_498), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_517), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_536), .B(n_461), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_546), .B(n_461), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_514), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_549), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_515), .B(n_460), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_508), .A2(n_476), .B1(n_493), .B2(n_497), .C(n_459), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_552), .B(n_479), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_554), .B(n_479), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_491), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_556), .B(n_491), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_549), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_514), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_557), .B(n_459), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_557), .B(n_470), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_553), .B(n_470), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_557), .B(n_470), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_543), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_558), .B(n_472), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_558), .B(n_472), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_543), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_559), .B(n_472), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_540), .B(n_497), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_560), .B(n_497), .Y(n_597) );
BUFx3_ASAP7_75t_L g598 ( .A(n_560), .Y(n_598) );
NOR2xp33_ASAP7_75t_SL g599 ( .A(n_507), .B(n_501), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_521), .B(n_473), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_544), .B(n_501), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_527), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_519), .A2(n_502), .B1(n_473), .B2(n_500), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_533), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_559), .B(n_473), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_561), .B(n_502), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_530), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_531), .Y(n_609) );
INVx5_ASAP7_75t_L g610 ( .A(n_545), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_545), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_547), .B(n_502), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_526), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_548), .B(n_500), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_598), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_564), .Y(n_616) );
AOI321xp33_ASAP7_75t_L g617 ( .A1(n_602), .A2(n_508), .A3(n_510), .B1(n_507), .B2(n_504), .C(n_522), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_567), .B(n_505), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_599), .B(n_512), .C(n_510), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_564), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_588), .B(n_600), .Y(n_621) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_576), .B(n_513), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_598), .Y(n_623) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_611), .A2(n_523), .B(n_518), .Y(n_624) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_611), .A2(n_516), .B(n_528), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_572), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_572), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_565), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_587), .Y(n_629) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_576), .B(n_545), .Y(n_630) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_566), .B(n_525), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_591), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_583), .Y(n_633) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_566), .B(n_524), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_588), .B(n_538), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_603), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_610), .B(n_541), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_603), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_595), .B(n_570), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_605), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_591), .B(n_542), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_593), .Y(n_642) );
OA22x2_ASAP7_75t_L g643 ( .A1(n_583), .A2(n_541), .B1(n_532), .B2(n_531), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_592), .B(n_537), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_596), .A2(n_534), .B(n_511), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_592), .B(n_534), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_593), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_594), .B(n_500), .Y(n_648) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_569), .A2(n_500), .B(n_535), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_606), .Y(n_650) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_563), .B(n_569), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_613), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g653 ( .A(n_568), .B(n_612), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_608), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_594), .B(n_562), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_SL g656 ( .A1(n_604), .A2(n_578), .B(n_608), .C(n_577), .Y(n_656) );
INVx2_ASAP7_75t_SL g657 ( .A(n_587), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g658 ( .A(n_612), .B(n_589), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_571), .A2(n_584), .B(n_579), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_601), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_606), .B(n_562), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_606), .A2(n_610), .B1(n_597), .B2(n_573), .Y(n_662) );
NAND2xp33_ASAP7_75t_SL g663 ( .A(n_580), .B(n_589), .Y(n_663) );
OAI32xp33_ASAP7_75t_L g664 ( .A1(n_574), .A2(n_580), .A3(n_614), .B1(n_581), .B2(n_582), .Y(n_664) );
XNOR2xp5_ASAP7_75t_L g665 ( .A(n_586), .B(n_597), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_614), .A2(n_597), .B1(n_607), .B2(n_586), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_609), .B(n_581), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_609), .B(n_610), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_575), .B(n_585), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_610), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_585), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_590), .B(n_582), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_633), .Y(n_673) );
OAI31xp33_ASAP7_75t_L g674 ( .A1(n_663), .A2(n_653), .A3(n_656), .B(n_619), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_651), .A2(n_618), .B(n_624), .C(n_630), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_615), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_659), .A2(n_619), .B(n_631), .Y(n_677) );
NOR2xp33_ASAP7_75t_SL g678 ( .A(n_623), .B(n_670), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_643), .A2(n_639), .B1(n_625), .B2(n_659), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_621), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_625), .A2(n_622), .B(n_672), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_664), .A2(n_624), .B(n_662), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_617), .A2(n_666), .B1(n_662), .B2(n_650), .C(n_654), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_617), .A2(n_632), .B(n_645), .C(n_661), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_657), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_652), .B(n_660), .Y(n_686) );
NAND5xp2_ASAP7_75t_L g687 ( .A(n_674), .B(n_645), .C(n_649), .D(n_668), .E(n_648), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_677), .A2(n_637), .B(n_628), .C(n_640), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_683), .A2(n_634), .B1(n_610), .B2(n_635), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_682), .A2(n_667), .B(n_658), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g691 ( .A1(n_675), .A2(n_646), .B(n_655), .C(n_626), .Y(n_691) );
OAI22xp5_ASAP7_75t_SL g692 ( .A1(n_679), .A2(n_665), .B1(n_629), .B2(n_644), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_681), .A2(n_636), .B1(n_638), .B2(n_627), .C(n_616), .Y(n_693) );
NAND3xp33_ASAP7_75t_SL g694 ( .A(n_678), .B(n_641), .C(n_620), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_692), .Y(n_695) );
NOR3xp33_ASAP7_75t_SL g696 ( .A(n_687), .B(n_684), .C(n_686), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_694), .A2(n_676), .B1(n_680), .B2(n_685), .Y(n_697) );
NAND3xp33_ASAP7_75t_SL g698 ( .A(n_691), .B(n_673), .C(n_669), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_690), .B(n_673), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_695), .B(n_688), .C(n_693), .Y(n_700) );
XOR2xp5_ASAP7_75t_L g701 ( .A(n_697), .B(n_689), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_699), .Y(n_702) );
AO22x2_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_698), .B1(n_696), .B2(n_647), .Y(n_703) );
XNOR2xp5_ASAP7_75t_L g704 ( .A(n_701), .B(n_642), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_703), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_705), .Y(n_706) );
XNOR2xp5_ASAP7_75t_L g707 ( .A(n_706), .B(n_704), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_700), .B(n_671), .Y(n_708) );
endmodule