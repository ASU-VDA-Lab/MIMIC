module fake_jpeg_26611_n_260 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_34),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_13),
.B1(n_24),
.B2(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_25),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_25),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_57),
.B1(n_60),
.B2(n_62),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_55),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_43),
.B(n_46),
.C(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_52),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_58),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_30),
.B1(n_31),
.B2(n_26),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_31),
.B1(n_36),
.B2(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_64),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_31),
.B1(n_19),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_36),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_45),
.C(n_39),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_72),
.C(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_60),
.B1(n_40),
.B2(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_78),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_29),
.A3(n_20),
.B1(n_45),
.B2(n_15),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_35),
.C(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_22),
.B(n_18),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_45),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_48),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_52),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_102),
.B(n_106),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_52),
.C(n_58),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_110),
.C(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_99),
.Y(n_117)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_49),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_61),
.Y(n_103)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_45),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_78),
.B1(n_79),
.B2(n_85),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_60),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_54),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_122),
.B1(n_123),
.B2(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_87),
.B1(n_81),
.B2(n_79),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_120),
.B1(n_16),
.B2(n_32),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_71),
.B1(n_70),
.B2(n_74),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_71),
.B1(n_62),
.B2(n_66),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_71),
.B1(n_62),
.B2(n_67),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_128),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_11),
.B(n_10),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_1),
.C(n_2),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_11),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_91),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_56),
.B1(n_20),
.B2(n_22),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_137),
.B1(n_141),
.B2(n_32),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_142),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_16),
.B1(n_22),
.B2(n_18),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_102),
.B1(n_100),
.B2(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_15),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_18),
.B(n_16),
.C(n_21),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_96),
.B(n_18),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_93),
.C(n_90),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_147),
.C(n_170),
.Y(n_179)
);

XOR2x2_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_91),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_169),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_90),
.C(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_155),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_153),
.B(n_162),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_95),
.B(n_98),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_168),
.B(n_171),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_1),
.B(n_2),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_14),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_15),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_163),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_21),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_15),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_12),
.B1(n_32),
.B2(n_14),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_125),
.C(n_120),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_32),
.B1(n_21),
.B2(n_5),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_3),
.B(n_4),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_137),
.B(n_4),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_145),
.C(n_147),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_190),
.C(n_163),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_131),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_193),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_144),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_191),
.B1(n_151),
.B2(n_118),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_172),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_122),
.C(n_123),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_159),
.B(n_140),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_139),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_167),
.B1(n_185),
.B2(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_158),
.C(n_148),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_197),
.C(n_174),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_149),
.C(n_161),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_165),
.B1(n_157),
.B2(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_149),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_153),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_196),
.C(n_199),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_174),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_215),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_192),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_190),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_183),
.B1(n_182),
.B2(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_188),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_226),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_207),
.C(n_189),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_192),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_219),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_215),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_212),
.C(n_211),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_231),
.B1(n_216),
.B2(n_230),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_239),
.C(n_134),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_238),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_213),
.B(n_175),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_173),
.B(n_186),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_214),
.C(n_118),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_134),
.B(n_5),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_3),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_5),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_6),
.C(n_7),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_238),
.B1(n_239),
.B2(n_8),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_249),
.B(n_250),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_243),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_252),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_6),
.B(n_7),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_256),
.C(n_9),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_9),
.Y(n_260)
);


endmodule