module fake_ariane_2839_n_1920 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1920);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1920;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_62),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_77),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_97),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_71),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_90),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_78),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_22),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_15),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_53),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_122),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_11),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_119),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_74),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_44),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_79),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_37),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_88),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_80),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_91),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_41),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_3),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_47),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_63),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_166),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_106),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_2),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_134),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_148),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_50),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_59),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_101),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_130),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_41),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_155),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_151),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_139),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_85),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_59),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_157),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_51),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_24),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_118),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_100),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_96),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_133),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_98),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_123),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_165),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_23),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_86),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_141),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_51),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_128),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_63),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_187),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_162),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_93),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_64),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_92),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_23),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_6),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_0),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_138),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_62),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_107),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_161),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_176),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_35),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_34),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_66),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_186),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_185),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_73),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_110),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_82),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_104),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_124),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_102),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_168),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_19),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_181),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_20),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_129),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_53),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_83),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_21),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_28),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_4),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_6),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_64),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_15),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_188),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_54),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_31),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_127),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_52),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_156),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_54),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_16),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_0),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_81),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_95),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_89),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_47),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_66),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_65),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_180),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_120),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_125),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_9),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_179),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_29),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_29),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_158),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_103),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_24),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_70),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_46),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_184),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_31),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_75),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_45),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_50),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_55),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_149),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_69),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_20),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_28),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_65),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_174),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_109),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_8),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_17),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_115),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_114),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_126),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_154),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_121),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_45),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_164),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_150),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_68),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_105),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_172),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_61),
.Y(n_369)
);

BUFx10_ASAP7_75t_L g370 ( 
.A(n_160),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_33),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_19),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_57),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_38),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_26),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_170),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_61),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_72),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_140),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_48),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_14),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_67),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_236),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_236),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_278),
.B(n_1),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_212),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_220),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_269),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_257),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_220),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_232),
.Y(n_392)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_225),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_257),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_229),
.B(n_2),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_225),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_242),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_370),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_246),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_272),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_247),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_208),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_273),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_285),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_208),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_209),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_308),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_209),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_272),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_325),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_365),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_370),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_370),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_190),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_7),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_248),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_202),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_248),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_282),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_308),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_282),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_353),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_308),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_203),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_377),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_206),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_287),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_206),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_229),
.B(n_7),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_195),
.B(n_10),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_204),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_207),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_287),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_291),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_291),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_305),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_293),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_305),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_307),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_214),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_216),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_293),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_298),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_218),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_298),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_307),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_195),
.B(n_12),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_224),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_322),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_322),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_334),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_328),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_357),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_227),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_334),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_329),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_328),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_329),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_234),
.B(n_12),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_333),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_333),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_234),
.B(n_13),
.Y(n_467)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_196),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_351),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_228),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_196),
.B(n_14),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_230),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_329),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_351),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_329),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_352),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_252),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_238),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_211),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_434),
.A2(n_200),
.B(n_199),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_419),
.A2(n_200),
.B(n_199),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_222),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_406),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_409),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_468),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_427),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_383),
.B(n_211),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_357),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_468),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_420),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_357),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_431),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_441),
.B(n_357),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_388),
.B(n_217),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_412),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_444),
.Y(n_518)
);

BUFx8_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_395),
.B(n_217),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_454),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_455),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_457),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_462),
.B(n_280),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_474),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_476),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_396),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_452),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_471),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_388),
.B(n_250),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_398),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_397),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_466),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_393),
.B(n_312),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_402),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_432),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_391),
.B(n_280),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_416),
.B(n_223),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_391),
.B(n_250),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_433),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_467),
.B(n_318),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_394),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_394),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_438),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_399),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_389),
.B(n_222),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_417),
.B(n_219),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_417),
.B(n_252),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_413),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_418),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_536),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_556),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_555),
.B(n_404),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_501),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_480),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_557),
.B(n_421),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_548),
.A2(n_318),
.B1(n_314),
.B2(n_276),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_482),
.Y(n_570)
);

BUFx6f_ASAP7_75t_SL g571 ( 
.A(n_552),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_487),
.A2(n_447),
.B1(n_448),
.B2(n_442),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_557),
.B(n_421),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_539),
.B(n_428),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_494),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_539),
.B(n_540),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_480),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_531),
.B(n_428),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_531),
.B(n_435),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_494),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_536),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_539),
.B(n_223),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_494),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_494),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_553),
.B(n_435),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_480),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_481),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_539),
.B(n_436),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_556),
.Y(n_596)
);

NOR2x1p5_ASAP7_75t_L g597 ( 
.A(n_501),
.B(n_436),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_494),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_481),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_445),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_495),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_516),
.B(n_405),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_501),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_481),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_495),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_533),
.B(n_219),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_487),
.A2(n_456),
.B1(n_460),
.B2(n_450),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_555),
.A2(n_326),
.B1(n_243),
.B2(n_254),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_487),
.A2(n_312),
.B1(n_344),
.B2(n_352),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_495),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_553),
.B(n_445),
.Y(n_613)
);

OAI21xp33_ASAP7_75t_SL g614 ( 
.A1(n_532),
.A2(n_374),
.B(n_356),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_532),
.A2(n_374),
.B1(n_356),
.B2(n_245),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_498),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_488),
.A2(n_331),
.B(n_378),
.C(n_376),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_495),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_540),
.B(n_446),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_495),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_507),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_543),
.B(n_446),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_499),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_489),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_490),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_536),
.B(n_344),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_507),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_507),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_516),
.B(n_449),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_499),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_484),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_507),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_484),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_498),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_507),
.Y(n_638)
);

NOR2x1p5_ASAP7_75t_L g639 ( 
.A(n_501),
.B(n_449),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_484),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_487),
.A2(n_461),
.B1(n_463),
.B2(n_475),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_491),
.B(n_453),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_499),
.Y(n_644)
);

CKINVDCx6p67_ASAP7_75t_R g645 ( 
.A(n_541),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_484),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_536),
.B(n_453),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_541),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_540),
.B(n_459),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_507),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_540),
.B(n_459),
.Y(n_651)
);

AND3x2_ASAP7_75t_L g652 ( 
.A(n_515),
.B(n_549),
.C(n_548),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_543),
.B(n_470),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_515),
.B(n_472),
.C(n_470),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_540),
.B(n_472),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_549),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_541),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_487),
.A2(n_473),
.B1(n_478),
.B2(n_252),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_520),
.B(n_277),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_485),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_507),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_551),
.B(n_478),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_500),
.B(n_194),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_507),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_485),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_551),
.B(n_415),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_554),
.Y(n_667)
);

INVxp33_ASAP7_75t_L g668 ( 
.A(n_538),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_485),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_512),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_538),
.B(n_239),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_498),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_538),
.B(n_255),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_512),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_512),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_554),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_483),
.B(n_256),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_535),
.B(n_266),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_485),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_486),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_486),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_512),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_486),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_500),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_504),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_545),
.B(n_270),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_483),
.B(n_279),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_493),
.B(n_237),
.Y(n_689)
);

INVxp33_ASAP7_75t_L g690 ( 
.A(n_537),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_487),
.A2(n_362),
.B1(n_277),
.B2(n_477),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_504),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_542),
.B(n_288),
.C(n_283),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_486),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_490),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_504),
.Y(n_696)
);

NOR2x1p5_ASAP7_75t_L g697 ( 
.A(n_541),
.B(n_550),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_546),
.B(n_289),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_486),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_512),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_542),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_546),
.B(n_292),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_504),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_512),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_552),
.A2(n_533),
.B1(n_544),
.B2(n_490),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_512),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_512),
.Y(n_707)
);

BUFx4f_ASAP7_75t_L g708 ( 
.A(n_490),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_486),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_486),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_624),
.B(n_544),
.C(n_493),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_688),
.B(n_647),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_483),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_653),
.B(n_526),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_603),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_561),
.B(n_526),
.Y(n_716)
);

AND2x6_ASAP7_75t_SL g717 ( 
.A(n_560),
.B(n_558),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_691),
.A2(n_552),
.B1(n_547),
.B2(n_490),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_561),
.B(n_526),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_568),
.B(n_387),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_565),
.B(n_493),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_587),
.B(n_526),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_574),
.B(n_392),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_587),
.B(n_526),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_565),
.B(n_591),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_562),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_647),
.B(n_493),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_577),
.B(n_493),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_564),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_607),
.A2(n_552),
.B1(n_547),
.B2(n_490),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_577),
.B(n_493),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_565),
.B(n_493),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_626),
.B(n_493),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_686),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_570),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_562),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_626),
.B(n_493),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_592),
.B(n_401),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_567),
.Y(n_739)
);

AND2x6_ASAP7_75t_SL g740 ( 
.A(n_613),
.B(n_558),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_596),
.B(n_537),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_642),
.B(n_547),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_550),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_591),
.B(n_498),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_583),
.B(n_585),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_690),
.B(n_403),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_567),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_570),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_642),
.B(n_547),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_575),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_596),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_603),
.Y(n_752)
);

CKINVDCx11_ASAP7_75t_R g753 ( 
.A(n_645),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_668),
.B(n_537),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_588),
.B(n_705),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_L g756 ( 
.A1(n_609),
.A2(n_534),
.B1(n_522),
.B2(n_527),
.C(n_529),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_631),
.B(n_407),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_685),
.B(n_547),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_575),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_686),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_566),
.B(n_550),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_671),
.B(n_550),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_591),
.B(n_498),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_591),
.B(n_506),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_685),
.B(n_547),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_566),
.B(n_537),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_692),
.B(n_504),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_604),
.B(n_408),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_563),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_625),
.B(n_506),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_696),
.B(n_504),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_L g772 ( 
.A(n_588),
.B(n_490),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_695),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_703),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_703),
.B(n_552),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_663),
.B(n_552),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_628),
.B(n_552),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_654),
.B(n_523),
.C(n_522),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_662),
.B(n_414),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_604),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_701),
.B(n_426),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_625),
.B(n_506),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_657),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_666),
.B(n_527),
.C(n_523),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_588),
.B(n_490),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_628),
.B(n_643),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_582),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_625),
.B(n_506),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_614),
.A2(n_488),
.B(n_513),
.C(n_510),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_593),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_593),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_594),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_628),
.B(n_552),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_671),
.B(n_525),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_708),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_607),
.A2(n_490),
.B1(n_552),
.B2(n_529),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_594),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_628),
.B(n_552),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_607),
.B(n_508),
.Y(n_799)
);

OR2x2_ASAP7_75t_SL g800 ( 
.A(n_678),
.B(n_429),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_625),
.B(n_506),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_600),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_605),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_605),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_615),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_701),
.B(n_534),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_659),
.B(n_508),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_659),
.B(n_508),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_708),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_673),
.B(n_525),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_708),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_659),
.A2(n_490),
.B1(n_518),
.B2(n_510),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_615),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_688),
.B(n_525),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_659),
.B(n_510),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_659),
.A2(n_490),
.B1(n_518),
.B2(n_511),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_578),
.B(n_511),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_633),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_620),
.B(n_511),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_632),
.B(n_492),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_633),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_636),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_632),
.B(n_492),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_695),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_609),
.B(n_518),
.C(n_513),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_632),
.B(n_492),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_632),
.B(n_492),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_695),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_636),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_601),
.B(n_513),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_640),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_649),
.B(n_530),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_651),
.B(n_530),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_640),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_656),
.B(n_667),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_588),
.A2(n_525),
.B1(n_524),
.B2(n_521),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_656),
.B(n_530),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_588),
.B(n_519),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_695),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_588),
.B(n_519),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_588),
.B(n_519),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_617),
.A2(n_488),
.B(n_496),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_646),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_637),
.B(n_519),
.Y(n_845)
);

O2A1O1Ixp5_ASAP7_75t_L g846 ( 
.A1(n_581),
.A2(n_497),
.B(n_496),
.C(n_505),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_672),
.B(n_519),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_667),
.B(n_677),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_648),
.B(n_517),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_576),
.B(n_496),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_652),
.B(n_519),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_646),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_660),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_658),
.B(n_525),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_678),
.B(n_525),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_644),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_660),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_610),
.B(n_528),
.Y(n_858)
);

NAND2x1_ASAP7_75t_L g859 ( 
.A(n_559),
.B(n_486),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_569),
.A2(n_616),
.B1(n_673),
.B2(n_573),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_579),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_571),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_595),
.B(n_528),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_579),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_616),
.B(n_528),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_580),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_693),
.A2(n_524),
.B1(n_521),
.B2(n_517),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_580),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_648),
.A2(n_517),
.B1(n_524),
.B2(n_521),
.Y(n_869)
);

INVxp33_ASAP7_75t_L g870 ( 
.A(n_608),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_584),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_614),
.B(n_528),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_669),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_679),
.B(n_530),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_669),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_726),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_729),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_846),
.A2(n_618),
.B(n_589),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_745),
.A2(n_644),
.B1(n_572),
.B2(n_635),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_821),
.A2(n_644),
.B(n_589),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_735),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_713),
.A2(n_698),
.B(n_702),
.C(n_687),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_712),
.B(n_641),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_836),
.B(n_697),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_843),
.A2(n_590),
.B(n_584),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_712),
.B(n_569),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_753),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_821),
.A2(n_644),
.B(n_598),
.Y(n_888)
);

AO21x1_ASAP7_75t_L g889 ( 
.A1(n_755),
.A2(n_598),
.B(n_590),
.Y(n_889)
);

NOR2x1_ASAP7_75t_L g890 ( 
.A(n_814),
.B(n_697),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_838),
.B(n_806),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_755),
.A2(n_606),
.B(n_611),
.C(n_602),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_824),
.A2(n_606),
.B(n_602),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_824),
.A2(n_612),
.B(n_611),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_827),
.A2(n_619),
.B(n_612),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_827),
.A2(n_621),
.B(n_619),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_828),
.A2(n_622),
.B(n_621),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_715),
.B(n_627),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_828),
.A2(n_623),
.B(n_622),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_734),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_714),
.A2(n_629),
.B(n_623),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_715),
.B(n_627),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_836),
.B(n_741),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_744),
.A2(n_680),
.B(n_675),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_848),
.A2(n_521),
.B(n_524),
.C(n_517),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_720),
.A2(n_303),
.B(n_301),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_815),
.B(n_569),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_763),
.A2(n_694),
.B(n_684),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_856),
.A2(n_572),
.B1(n_635),
.B2(n_559),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_SL g910 ( 
.A1(n_725),
.A2(n_629),
.B(n_634),
.C(n_630),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_815),
.B(n_569),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_764),
.A2(n_634),
.B(n_630),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_752),
.B(n_597),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_752),
.A2(n_683),
.B(n_661),
.C(n_707),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_739),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_809),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_723),
.B(n_639),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_855),
.A2(n_683),
.B(n_661),
.C(n_707),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_780),
.B(n_639),
.Y(n_919)
);

OAI22xp33_ASAP7_75t_L g920 ( 
.A1(n_780),
.A2(n_372),
.B1(n_309),
.B2(n_310),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_748),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_783),
.B(n_528),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_786),
.B(n_528),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_825),
.B(n_627),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_753),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_742),
.B(n_528),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_764),
.A2(n_709),
.B(n_699),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_749),
.B(n_689),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_825),
.B(n_627),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_814),
.B(n_502),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_734),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_747),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_809),
.B(n_627),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_747),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_757),
.A2(n_664),
.B1(n_706),
.B2(n_704),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_770),
.A2(n_650),
.B(n_638),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_782),
.A2(n_710),
.B(n_670),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_795),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_738),
.A2(n_664),
.B1(n_706),
.B2(n_704),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_795),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_782),
.A2(n_674),
.B(n_670),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_825),
.B(n_627),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_794),
.A2(n_700),
.B(n_674),
.C(n_676),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_788),
.A2(n_700),
.B(n_676),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_820),
.A2(n_710),
.B(n_682),
.C(n_681),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_758),
.B(n_765),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_754),
.B(n_572),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_746),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_767),
.B(n_635),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_788),
.A2(n_801),
.B(n_799),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_801),
.A2(n_681),
.B(n_665),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_825),
.B(n_576),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_829),
.B(n_576),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_750),
.A2(n_681),
.B1(n_665),
.B2(n_682),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_800),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_850),
.A2(n_682),
.B(n_665),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_850),
.A2(n_497),
.B(n_496),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_766),
.B(n_502),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_727),
.A2(n_503),
.B(n_497),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_716),
.A2(n_503),
.B(n_497),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_771),
.B(n_810),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_736),
.B(n_576),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_719),
.A2(n_505),
.B(n_503),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_849),
.A2(n_779),
.B1(n_756),
.B2(n_860),
.Y(n_964)
);

NAND2x1_ASAP7_75t_L g965 ( 
.A(n_829),
.B(n_576),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_751),
.B(n_586),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_725),
.A2(n_505),
.B(n_503),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_722),
.A2(n_724),
.B(n_721),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_760),
.B(n_509),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_807),
.A2(n_262),
.B(n_245),
.C(n_251),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_808),
.A2(n_262),
.B(n_251),
.C(n_253),
.Y(n_971)
);

INVx11_ASAP7_75t_L g972 ( 
.A(n_862),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_721),
.A2(n_505),
.B(n_586),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_732),
.A2(n_599),
.B(n_586),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_816),
.A2(n_263),
.B(n_253),
.C(n_284),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_732),
.A2(n_831),
.B(n_818),
.Y(n_976)
);

BUFx4f_ASAP7_75t_L g977 ( 
.A(n_743),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_711),
.A2(n_520),
.B(n_514),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_795),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_743),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_759),
.A2(n_509),
.B(n_514),
.C(n_263),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_778),
.A2(n_315),
.B(n_311),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_863),
.A2(n_599),
.B(n_586),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_743),
.B(n_502),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_872),
.A2(n_789),
.B(n_861),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_781),
.B(n_509),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_859),
.A2(n_599),
.B(n_514),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_787),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_795),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_853),
.A2(n_599),
.B(n_514),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_826),
.A2(n_320),
.B(n_316),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_853),
.A2(n_599),
.B(n_514),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_762),
.B(n_509),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_789),
.A2(n_514),
.B(n_509),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_857),
.A2(n_509),
.B(n_290),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_768),
.B(n_321),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_857),
.A2(n_290),
.B(n_284),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_774),
.B(n_327),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_761),
.B(n_335),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_792),
.Y(n_1000)
);

AOI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_870),
.A2(n_337),
.B(n_336),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_833),
.A2(n_295),
.B(n_350),
.C(n_354),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_743),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_870),
.B(n_340),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_873),
.A2(n_192),
.B(n_191),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_769),
.B(n_342),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_811),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_784),
.B(n_346),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_811),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_834),
.B(n_348),
.C(n_347),
.Y(n_1010)
);

BUFx12f_ASAP7_75t_L g1011 ( 
.A(n_717),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_869),
.A2(n_295),
.B(n_324),
.C(n_331),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_854),
.B(n_363),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_837),
.B(n_366),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_SL g1015 ( 
.A(n_862),
.B(n_571),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_867),
.A2(n_369),
.B(n_371),
.Y(n_1016)
);

OAI22x1_ASAP7_75t_L g1017 ( 
.A1(n_812),
.A2(n_817),
.B1(n_796),
.B2(n_740),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_865),
.B(n_874),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_730),
.B(n_373),
.Y(n_1019)
);

AOI33xp33_ASAP7_75t_L g1020 ( 
.A1(n_864),
.A2(n_324),
.A3(n_332),
.B1(n_339),
.B2(n_350),
.B3(n_354),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_866),
.A2(n_378),
.B(n_376),
.C(n_368),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_858),
.A2(n_479),
.B(n_332),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_790),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_773),
.A2(n_339),
.B(n_368),
.C(n_382),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_791),
.B(n_380),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_718),
.B(n_479),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_862),
.B(n_851),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_811),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_775),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_797),
.B(n_479),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_873),
.A2(n_205),
.B(n_379),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_868),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_773),
.A2(n_571),
.B1(n_210),
.B2(n_213),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_803),
.B(n_813),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_811),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_829),
.B(n_193),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_728),
.B(n_197),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_875),
.A2(n_201),
.B(n_361),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_871),
.A2(n_198),
.B(n_360),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_875),
.A2(n_367),
.B(n_359),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_773),
.A2(n_358),
.B1(n_355),
.B2(n_349),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_731),
.B(n_215),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_802),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_840),
.A2(n_345),
.B(n_343),
.C(n_341),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_813),
.B(n_221),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_840),
.A2(n_338),
.B(n_330),
.C(n_319),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_819),
.B(n_226),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_804),
.B(n_18),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_772),
.B(n_313),
.C(n_244),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_772),
.A2(n_785),
.B(n_737),
.C(n_733),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_840),
.A2(n_306),
.B(n_249),
.C(n_241),
.Y(n_1051)
);

OAI21xp33_ASAP7_75t_SL g1052 ( 
.A1(n_985),
.A2(n_847),
.B(n_845),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_948),
.B(n_805),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_876),
.B(n_822),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_892),
.A2(n_785),
.B(n_832),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_964),
.B(n_839),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_930),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_906),
.A2(n_776),
.B(n_835),
.C(n_842),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_1012),
.A2(n_841),
.B(n_793),
.C(n_777),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1001),
.A2(n_798),
.B(n_844),
.C(n_830),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_959),
.A2(n_852),
.B(n_844),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_961),
.A2(n_830),
.B1(n_823),
.B2(n_819),
.Y(n_1062)
);

INVx8_ASAP7_75t_L g1063 ( 
.A(n_1028),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_881),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_920),
.A2(n_852),
.B(n_823),
.C(n_25),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_917),
.B(n_231),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_SL g1067 ( 
.A(n_999),
.B(n_233),
.C(n_235),
.Y(n_1067)
);

OA22x2_ASAP7_75t_L g1068 ( 
.A1(n_903),
.A2(n_240),
.B1(n_259),
.B2(n_260),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_877),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_930),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_921),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_887),
.B(n_261),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_900),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_996),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_1003),
.B(n_222),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_984),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1008),
.A2(n_21),
.B(n_22),
.C(n_25),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_986),
.B(n_27),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_958),
.B(n_264),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_958),
.B(n_281),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_884),
.B(n_30),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_882),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_886),
.B(n_32),
.Y(n_1083)
);

INVx6_ASAP7_75t_L g1084 ( 
.A(n_925),
.Y(n_1084)
);

AOI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_1017),
.A2(n_222),
.B(n_258),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_900),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_883),
.B(n_35),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_993),
.A2(n_286),
.B1(n_304),
.B2(n_265),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_890),
.B(n_36),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_959),
.A2(n_294),
.B(n_317),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1004),
.B(n_37),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_962),
.B(n_38),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1023),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1006),
.B(n_267),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_913),
.B(n_268),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_955),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1043),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_900),
.Y(n_1098)
);

OAI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_982),
.A2(n_296),
.B1(n_300),
.B2(n_271),
.C(n_274),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_979),
.B(n_275),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_919),
.A2(n_302),
.B1(n_299),
.B2(n_297),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_939),
.A2(n_258),
.B1(n_40),
.B2(n_42),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_972),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1025),
.B(n_39),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_901),
.A2(n_258),
.B(n_116),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_977),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_1032),
.B(n_40),
.C(n_42),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_SL g1108 ( 
.A(n_977),
.B(n_258),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_976),
.A2(n_117),
.B(n_183),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_946),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_1110)
);

AO21x1_ASAP7_75t_L g1111 ( 
.A1(n_1018),
.A2(n_323),
.B(n_250),
.Y(n_1111)
);

BUFx8_ASAP7_75t_L g1112 ( 
.A(n_1011),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_966),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_935),
.A2(n_994),
.B1(n_1048),
.B2(n_1024),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_928),
.B(n_323),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_976),
.A2(n_135),
.B(n_175),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_907),
.B(n_43),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_915),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_931),
.B(n_49),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_979),
.B(n_323),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_885),
.A2(n_113),
.B(n_173),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1014),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_932),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_980),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_922),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1029),
.B(n_323),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_980),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_931),
.B(n_56),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_879),
.A2(n_136),
.B(n_167),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_934),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_979),
.B(n_323),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1010),
.B(n_56),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_916),
.B(n_989),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_1015),
.B(n_142),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_L g1135 ( 
.A(n_991),
.B(n_57),
.C(n_58),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_911),
.A2(n_1016),
.B1(n_1041),
.B2(n_1039),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_943),
.A2(n_323),
.B(n_250),
.C(n_67),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_998),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_SL g1139 ( 
.A(n_1044),
.B(n_58),
.C(n_60),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_989),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_988),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1020),
.B(n_60),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_989),
.Y(n_1143)
);

AO32x1_ASAP7_75t_L g1144 ( 
.A1(n_954),
.A2(n_68),
.A3(n_323),
.B1(n_250),
.B2(n_144),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1027),
.A2(n_250),
.B1(n_99),
.B2(n_145),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_914),
.A2(n_250),
.B(n_159),
.C(n_163),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1013),
.B(n_94),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_1007),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_968),
.A2(n_250),
.B(n_960),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_968),
.A2(n_950),
.B(n_878),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_L g1151 ( 
.A(n_1007),
.B(n_1049),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1002),
.A2(n_978),
.B(n_918),
.C(n_1050),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1007),
.B(n_938),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_960),
.A2(n_963),
.B(n_956),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_940),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_905),
.A2(n_970),
.B(n_971),
.C(n_975),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_933),
.B(n_940),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_947),
.B(n_1000),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_963),
.A2(n_956),
.B(n_967),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1009),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_898),
.A2(n_902),
.B1(n_1037),
.B2(n_1042),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_949),
.A2(n_1019),
.B1(n_969),
.B2(n_923),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1009),
.B(n_1035),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_SL g1164 ( 
.A(n_1046),
.B(n_1051),
.C(n_1040),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1033),
.B(n_909),
.Y(n_1166)
);

O2A1O1Ixp5_ASAP7_75t_L g1167 ( 
.A1(n_1036),
.A2(n_889),
.B(n_953),
.C(n_952),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_981),
.B(n_933),
.Y(n_1168)
);

NOR2x1_ASAP7_75t_L g1169 ( 
.A(n_1031),
.B(n_1040),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1034),
.B(n_926),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1031),
.B(n_1038),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_965),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1022),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_990),
.B(n_992),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_924),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_SL g1176 ( 
.A(n_974),
.B(n_987),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_997),
.B(n_990),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_992),
.B(n_1030),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1038),
.B(n_941),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1026),
.A2(n_945),
.B1(n_987),
.B2(n_880),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_912),
.B(n_936),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_895),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_904),
.A2(n_927),
.B(n_908),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1021),
.A2(n_910),
.B(n_1005),
.C(n_951),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_951),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_929),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_995),
.B(n_944),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_944),
.A2(n_973),
.B(n_974),
.C(n_893),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_973),
.A2(n_899),
.B(n_897),
.C(n_893),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_894),
.B(n_896),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_995),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_983),
.A2(n_897),
.B(n_899),
.Y(n_1192)
);

CKINVDCx6p67_ASAP7_75t_R g1193 ( 
.A(n_942),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_894),
.B(n_896),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1106),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1103),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1150),
.A2(n_983),
.B(n_957),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1190),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1070),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1190),
.Y(n_1200)
);

BUFx10_ASAP7_75t_L g1201 ( 
.A(n_1084),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1057),
.B(n_1054),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_1063),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1154),
.A2(n_937),
.B(n_888),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1159),
.A2(n_1149),
.B(n_1183),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1114),
.A2(n_1102),
.B(n_1056),
.Y(n_1206)
);

AO32x2_ASAP7_75t_L g1207 ( 
.A1(n_1102),
.A2(n_1180),
.A3(n_1162),
.B1(n_1110),
.B2(n_1114),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1150),
.A2(n_1052),
.B(n_1178),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1063),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1053),
.B(n_1113),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1066),
.B(n_1138),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1063),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1188),
.A2(n_1189),
.B(n_1061),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1132),
.A2(n_1122),
.B1(n_1104),
.B2(n_1135),
.C(n_1107),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1174),
.A2(n_1166),
.B(n_1162),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1170),
.A2(n_1194),
.B(n_1177),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_SL g1217 ( 
.A1(n_1082),
.A2(n_1122),
.B1(n_1110),
.B2(n_1137),
.C(n_1077),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1170),
.A2(n_1187),
.B(n_1181),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1084),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1173),
.A2(n_1105),
.B(n_1109),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1152),
.A2(n_1136),
.B(n_1167),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1176),
.A2(n_1111),
.B(n_1179),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1182),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1091),
.A2(n_1065),
.B(n_1171),
.C(n_1161),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1121),
.A2(n_1055),
.B(n_1129),
.Y(n_1225)
);

INVx3_ASAP7_75t_SL g1226 ( 
.A(n_1128),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1076),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1124),
.B(n_1127),
.Y(n_1228)
);

AO22x2_ASAP7_75t_L g1229 ( 
.A1(n_1074),
.A2(n_1165),
.B1(n_1083),
.B2(n_1125),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1095),
.A2(n_1089),
.B1(n_1119),
.B2(n_1081),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1106),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1062),
.A2(n_1115),
.A3(n_1146),
.B(n_1156),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1071),
.B(n_1093),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1092),
.A2(n_1055),
.B(n_1067),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1062),
.A2(n_1186),
.A3(n_1160),
.B1(n_1140),
.B2(n_1192),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_L g1236 ( 
.A(n_1155),
.B(n_1072),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1097),
.B(n_1106),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1059),
.A2(n_1078),
.B(n_1090),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1184),
.A2(n_1185),
.B(n_1116),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1125),
.B(n_1128),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1089),
.Y(n_1241)
);

AO32x2_ASAP7_75t_L g1242 ( 
.A1(n_1192),
.A2(n_1144),
.A3(n_1085),
.B1(n_1117),
.B2(n_1139),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1069),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1115),
.A2(n_1126),
.A3(n_1158),
.B(n_1087),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1164),
.C(n_1058),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1175),
.B(n_1096),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1148),
.B(n_1098),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1073),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1108),
.A2(n_1168),
.B(n_1157),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1118),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1112),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1123),
.B(n_1130),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1169),
.A2(n_1060),
.B(n_1126),
.Y(n_1253)
);

O2A1O1Ixp5_ASAP7_75t_SL g1254 ( 
.A1(n_1133),
.A2(n_1153),
.B(n_1131),
.C(n_1120),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1141),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1191),
.A2(n_1142),
.B(n_1145),
.C(n_1151),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1148),
.B(n_1098),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1068),
.B(n_1086),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1079),
.A2(n_1080),
.B1(n_1088),
.B2(n_1193),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1163),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1108),
.A2(n_1101),
.B(n_1100),
.C(n_1157),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1068),
.A2(n_1075),
.B(n_1144),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1144),
.A2(n_1075),
.A3(n_1172),
.B(n_1099),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_SL g1264 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1086),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1098),
.A2(n_1148),
.B(n_1143),
.C(n_1134),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1075),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1143),
.A2(n_1112),
.B(n_891),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1269)
);

BUFx8_ASAP7_75t_L g1270 ( 
.A(n_1057),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1094),
.A2(n_891),
.B(n_745),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1094),
.A2(n_891),
.B1(n_720),
.B2(n_723),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1176),
.A2(n_1154),
.B(n_1159),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1094),
.A2(n_723),
.B(n_720),
.C(n_653),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1190),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1063),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1149),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1094),
.A2(n_745),
.B(n_653),
.C(n_624),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1111),
.A2(n_1171),
.A3(n_889),
.B(n_1162),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1063),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1094),
.B(n_720),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1149),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1053),
.B(n_903),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1094),
.B(n_720),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1111),
.A2(n_1085),
.B(n_1154),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1149),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1190),
.Y(n_1291)
);

OAI22x1_ASAP7_75t_L g1292 ( 
.A1(n_1094),
.A2(n_609),
.B1(n_723),
.B2(n_720),
.Y(n_1292)
);

BUFx5_ASAP7_75t_L g1293 ( 
.A(n_1191),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1190),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1063),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1094),
.A2(n_745),
.B(n_653),
.C(n_624),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1094),
.B(n_720),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1111),
.A2(n_1171),
.A3(n_889),
.B(n_1162),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1053),
.B(n_903),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_SL g1301 ( 
.A1(n_1137),
.A2(n_891),
.B(n_1152),
.C(n_1181),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1094),
.A2(n_891),
.B(n_745),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1094),
.A2(n_745),
.B(n_653),
.C(n_624),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1094),
.A2(n_891),
.B1(n_720),
.B2(n_723),
.Y(n_1305)
);

O2A1O1Ixp5_ASAP7_75t_L g1306 ( 
.A1(n_1176),
.A2(n_1166),
.B(n_720),
.C(n_723),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1114),
.A2(n_891),
.B(n_1178),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1149),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1057),
.B(n_715),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1111),
.A2(n_1171),
.A3(n_889),
.B(n_1162),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1190),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1150),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1111),
.A2(n_1171),
.A3(n_889),
.B(n_1162),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1124),
.B(n_1127),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1053),
.B(n_903),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1094),
.A2(n_723),
.B(n_720),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1063),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1149),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1069),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1111),
.A2(n_1171),
.A3(n_889),
.B(n_1162),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1063),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1094),
.A2(n_738),
.B1(n_720),
.B2(n_723),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1190),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_SL g1329 ( 
.A1(n_1137),
.A2(n_891),
.B(n_1152),
.C(n_1181),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1064),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1063),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1332)
);

AO22x2_ASAP7_75t_L g1333 ( 
.A1(n_1114),
.A2(n_1102),
.B1(n_886),
.B2(n_911),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1054),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1053),
.B(n_903),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1150),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1150),
.A2(n_891),
.B(n_1052),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1106),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1106),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1069),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1053),
.B(n_903),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1094),
.A2(n_891),
.B1(n_720),
.B2(n_723),
.Y(n_1342)
);

OAI22x1_ASAP7_75t_L g1343 ( 
.A1(n_1094),
.A2(n_609),
.B1(n_723),
.B2(n_720),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1094),
.A2(n_891),
.B(n_745),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1203),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1284),
.A2(n_1288),
.B1(n_1298),
.B2(n_1342),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1273),
.A2(n_1305),
.B1(n_1327),
.B2(n_1292),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1233),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1230),
.A2(n_1344),
.B1(n_1272),
.B2(n_1303),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1201),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1320),
.A2(n_1343),
.B1(n_1214),
.B2(n_1206),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1201),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1330),
.Y(n_1353)
);

BUFx4_ASAP7_75t_SL g1354 ( 
.A(n_1251),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1196),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1287),
.A2(n_1341),
.B1(n_1300),
.B2(n_1335),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1219),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1226),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1221),
.B2(n_1211),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1270),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1319),
.A2(n_1210),
.B1(n_1334),
.B2(n_1215),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1270),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1250),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1278),
.Y(n_1364)
);

INVx8_ASAP7_75t_L g1365 ( 
.A(n_1247),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1333),
.A2(n_1229),
.B1(n_1234),
.B2(n_1240),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1259),
.A2(n_1286),
.B1(n_1309),
.B2(n_1271),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1250),
.Y(n_1368)
);

BUFx4f_ASAP7_75t_L g1369 ( 
.A(n_1195),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1255),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_1212),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1195),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1209),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1255),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1283),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1280),
.A2(n_1304),
.B1(n_1297),
.B2(n_1275),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1252),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1202),
.B(n_1199),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_SL g1379 ( 
.A(n_1228),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1241),
.A2(n_1258),
.B1(n_1337),
.B2(n_1269),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1296),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1321),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1340),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1326),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1246),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1307),
.A2(n_1224),
.B1(n_1323),
.B2(n_1295),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1223),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1241),
.A2(n_1332),
.B1(n_1277),
.B2(n_1282),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1227),
.B(n_1310),
.Y(n_1390)
);

CKINVDCx11_ASAP7_75t_R g1391 ( 
.A(n_1331),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1302),
.A2(n_1313),
.B1(n_1315),
.B2(n_1318),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1267),
.B(n_1264),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1238),
.A2(n_1328),
.B1(n_1312),
.B2(n_1198),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1267),
.A2(n_1207),
.B1(n_1217),
.B2(n_1249),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1195),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_1317),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1256),
.A2(n_1268),
.B1(n_1225),
.B2(n_1245),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1267),
.A2(n_1262),
.B1(n_1207),
.B2(n_1208),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1317),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1247),
.B(n_1257),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1231),
.B(n_1339),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1231),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1339),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1266),
.A2(n_1261),
.B(n_1216),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1207),
.A2(n_1237),
.B1(n_1239),
.B2(n_1306),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1339),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1248),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1260),
.Y(n_1409)
);

INVx6_ASAP7_75t_L g1410 ( 
.A(n_1293),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1198),
.A2(n_1291),
.B1(n_1200),
.B2(n_1276),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1200),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1338),
.A2(n_1329),
.B1(n_1301),
.B2(n_1236),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1276),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1291),
.Y(n_1415)
);

BUFx2_ASAP7_75t_SL g1416 ( 
.A(n_1338),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1294),
.A2(n_1328),
.B1(n_1312),
.B2(n_1293),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1294),
.A2(n_1293),
.B1(n_1218),
.B2(n_1289),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1197),
.A2(n_1265),
.B1(n_1336),
.B2(n_1314),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1235),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1235),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1293),
.A2(n_1242),
.B1(n_1314),
.B2(n_1253),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1213),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1254),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1222),
.A2(n_1274),
.B1(n_1242),
.B2(n_1232),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1204),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1232),
.A2(n_1263),
.B1(n_1325),
.B2(n_1316),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1235),
.Y(n_1428)
);

OAI22x1_ASAP7_75t_L g1429 ( 
.A1(n_1263),
.A2(n_1232),
.B1(n_1244),
.B2(n_1316),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1244),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1220),
.A2(n_1205),
.B1(n_1279),
.B2(n_1322),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1281),
.A2(n_1299),
.B1(n_1311),
.B2(n_1316),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1325),
.Y(n_1433)
);

BUFx2_ASAP7_75t_R g1434 ( 
.A(n_1281),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1299),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1299),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1325),
.Y(n_1437)
);

AOI22x1_ASAP7_75t_SL g1438 ( 
.A1(n_1311),
.A2(n_1285),
.B1(n_1290),
.B2(n_1308),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1311),
.A2(n_569),
.B1(n_1288),
.B2(n_1284),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1440)
);

BUFx10_ASAP7_75t_L g1441 ( 
.A(n_1251),
.Y(n_1441)
);

INVx4_ASAP7_75t_SL g1442 ( 
.A(n_1226),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1251),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1230),
.A2(n_1342),
.B1(n_1273),
.B2(n_1305),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1201),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1201),
.Y(n_1446)
);

CKINVDCx6p67_ASAP7_75t_R g1447 ( 
.A(n_1226),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1284),
.A2(n_1288),
.B1(n_1298),
.B2(n_1327),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1450)
);

BUFx8_ASAP7_75t_SL g1451 ( 
.A(n_1251),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1284),
.A2(n_1288),
.B1(n_1298),
.B2(n_1327),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1230),
.A2(n_1342),
.B1(n_1273),
.B2(n_1305),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1284),
.A2(n_1288),
.B1(n_1298),
.B2(n_1327),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1201),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1201),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1202),
.Y(n_1457)
);

INVx4_ASAP7_75t_SL g1458 ( 
.A(n_1226),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1243),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1201),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1201),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1463)
);

BUFx10_ASAP7_75t_L g1464 ( 
.A(n_1251),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1284),
.A2(n_1288),
.B1(n_1298),
.B2(n_1327),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1219),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1240),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1243),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1219),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1284),
.A2(n_569),
.B1(n_1298),
.B2(n_1288),
.Y(n_1470)
);

BUFx5_ASAP7_75t_L g1471 ( 
.A(n_1198),
.Y(n_1471)
);

BUFx8_ASAP7_75t_L g1472 ( 
.A(n_1212),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1230),
.A2(n_1342),
.B1(n_1273),
.B2(n_1305),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1284),
.A2(n_1298),
.B1(n_1288),
.B2(n_860),
.Y(n_1475)
);

CKINVDCx16_ASAP7_75t_R g1476 ( 
.A(n_1360),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1346),
.A2(n_1454),
.B1(n_1452),
.B2(n_1449),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1412),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1423),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1387),
.A2(n_1392),
.B(n_1367),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1431),
.A2(n_1419),
.B(n_1425),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1388),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1418),
.A2(n_1422),
.B(n_1389),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1414),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1398),
.A2(n_1376),
.B(n_1429),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1418),
.A2(n_1422),
.B(n_1389),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1415),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1363),
.Y(n_1488)
);

AOI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1436),
.A2(n_1435),
.B(n_1433),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1457),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1368),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1370),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1346),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1436),
.B(n_1421),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1374),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1353),
.B(n_1471),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1471),
.B(n_1394),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1430),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1410),
.Y(n_1499)
);

OR2x2_ASAP7_75t_SL g1500 ( 
.A(n_1420),
.B(n_1378),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1471),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1471),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1380),
.A2(n_1405),
.B(n_1394),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1471),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1390),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1471),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1417),
.A2(n_1413),
.B(n_1393),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1420),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1393),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1411),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1411),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1428),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1437),
.A2(n_1426),
.B(n_1366),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1432),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1432),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1366),
.A2(n_1351),
.B(n_1347),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1440),
.A2(n_1475),
.B1(n_1463),
.B2(n_1448),
.C(n_1462),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1424),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1427),
.A2(n_1367),
.B(n_1399),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1427),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1381),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1434),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1438),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1403),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1442),
.B(n_1458),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1395),
.B(n_1406),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1364),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1401),
.A2(n_1348),
.B(n_1377),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1399),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1395),
.B(n_1406),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1451),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1365),
.B(n_1467),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1345),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1467),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1383),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1401),
.A2(n_1402),
.B(n_1407),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1384),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1372),
.Y(n_1538)
);

AO21x1_ASAP7_75t_L g1539 ( 
.A1(n_1444),
.A2(n_1474),
.B(n_1453),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1409),
.A2(n_1459),
.B(n_1468),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1361),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1361),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1359),
.B(n_1450),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1472),
.Y(n_1544)
);

OR2x6_ASAP7_75t_L g1545 ( 
.A(n_1365),
.B(n_1416),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1442),
.B(n_1458),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1440),
.A2(n_1475),
.B(n_1450),
.C(n_1473),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1356),
.B(n_1349),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1349),
.B(n_1474),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1396),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1359),
.B(n_1463),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1444),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1439),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1439),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1442),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1445),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1448),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1462),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1473),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1458),
.B(n_1404),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1385),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1470),
.B(n_1386),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1470),
.B(n_1469),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1408),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1379),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1369),
.A2(n_1379),
.B(n_1391),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1357),
.B(n_1466),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1445),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1445),
.Y(n_1569)
);

INVx5_ASAP7_75t_L g1570 ( 
.A(n_1397),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1382),
.A2(n_1461),
.B(n_1400),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1456),
.B(n_1460),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1456),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1447),
.A2(n_1382),
.B1(n_1375),
.B2(n_1373),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1350),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1352),
.Y(n_1576)
);

AO32x1_ASAP7_75t_L g1577 ( 
.A1(n_1477),
.A2(n_1371),
.A3(n_1354),
.B1(n_1358),
.B2(n_1362),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1481),
.A2(n_1455),
.B(n_1446),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1493),
.A2(n_1354),
.B(n_1441),
.C(n_1464),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1505),
.B(n_1441),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1534),
.B(n_1490),
.Y(n_1581)
);

AO32x2_ASAP7_75t_L g1582 ( 
.A1(n_1556),
.A2(n_1355),
.A3(n_1443),
.B1(n_1464),
.B2(n_1538),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_SL g1583 ( 
.A(n_1532),
.B(n_1545),
.Y(n_1583)
);

O2A1O1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1539),
.A2(n_1549),
.B(n_1547),
.C(n_1548),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1517),
.A2(n_1543),
.B(n_1551),
.C(n_1548),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1480),
.A2(n_1503),
.B(n_1552),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1521),
.B(n_1561),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1535),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1539),
.B(n_1569),
.Y(n_1589)
);

NOR2x1_ASAP7_75t_SL g1590 ( 
.A(n_1532),
.B(n_1545),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1482),
.B(n_1494),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1512),
.Y(n_1592)
);

BUFx12f_ASAP7_75t_L g1593 ( 
.A(n_1544),
.Y(n_1593)
);

OR2x6_ASAP7_75t_L g1594 ( 
.A(n_1532),
.B(n_1525),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1541),
.A2(n_1542),
.B(n_1530),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1519),
.A2(n_1541),
.B(n_1545),
.Y(n_1596)
);

AO32x2_ASAP7_75t_L g1597 ( 
.A1(n_1556),
.A2(n_1538),
.A3(n_1550),
.B1(n_1569),
.B2(n_1555),
.Y(n_1597)
);

O2A1O1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1557),
.A2(n_1558),
.B(n_1559),
.C(n_1518),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1567),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1518),
.B(n_1559),
.C(n_1558),
.D(n_1557),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1527),
.B(n_1576),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1526),
.A2(n_1485),
.B(n_1510),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1562),
.A2(n_1529),
.B(n_1523),
.C(n_1511),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1485),
.A2(n_1516),
.B(n_1507),
.Y(n_1605)
);

AO32x2_ASAP7_75t_L g1606 ( 
.A1(n_1550),
.A2(n_1569),
.A3(n_1555),
.B1(n_1500),
.B2(n_1494),
.Y(n_1606)
);

INVxp33_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1520),
.A2(n_1514),
.B1(n_1515),
.B2(n_1529),
.C(n_1553),
.Y(n_1608)
);

A2O1A1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1563),
.A2(n_1554),
.B(n_1522),
.C(n_1497),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1518),
.A2(n_1516),
.B(n_1519),
.C(n_1575),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1573),
.B(n_1564),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1533),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1478),
.A2(n_1484),
.B1(n_1487),
.B2(n_1495),
.C(n_1492),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1576),
.B(n_1544),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1496),
.B(n_1525),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1545),
.A2(n_1486),
.B(n_1483),
.Y(n_1617)
);

OAI21xp33_ASAP7_75t_L g1618 ( 
.A1(n_1488),
.A2(n_1495),
.B(n_1492),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1491),
.B(n_1568),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1566),
.A2(n_1571),
.B(n_1546),
.C(n_1525),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1528),
.A2(n_1486),
.B(n_1483),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1535),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1537),
.Y(n_1623)
);

AO32x2_ASAP7_75t_L g1624 ( 
.A1(n_1555),
.A2(n_1540),
.A3(n_1508),
.B1(n_1528),
.B2(n_1537),
.Y(n_1624)
);

NOR2x1_ASAP7_75t_SL g1625 ( 
.A(n_1532),
.B(n_1572),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1483),
.A2(n_1486),
.B(n_1536),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1483),
.A2(n_1486),
.B(n_1536),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1501),
.A2(n_1502),
.B(n_1504),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1570),
.A2(n_1532),
.B1(n_1476),
.B2(n_1509),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1628),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1600),
.A2(n_1513),
.B1(n_1565),
.B2(n_1570),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1592),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1613),
.B(n_1506),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1628),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1597),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1588),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1581),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1624),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1624),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1589),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1610),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1624),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1591),
.B(n_1479),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1578),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1593),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1594),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1622),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1623),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1619),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1618),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1594),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1625),
.B(n_1499),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1583),
.B(n_1590),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1614),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1498),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1626),
.B(n_1627),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1587),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1607),
.B(n_1572),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1626),
.B(n_1489),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1635),
.B(n_1578),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1654),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1641),
.A2(n_1605),
.B(n_1621),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1634),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1630),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1636),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1652),
.B(n_1617),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1654),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1630),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1641),
.A2(n_1584),
.B(n_1585),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1635),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1654),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1636),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1586),
.Y(n_1674)
);

INVx5_ASAP7_75t_L g1675 ( 
.A(n_1652),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1636),
.Y(n_1676)
);

AOI33xp33_ASAP7_75t_L g1677 ( 
.A1(n_1655),
.A2(n_1598),
.A3(n_1577),
.B1(n_1580),
.B2(n_1608),
.B3(n_1611),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1647),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1644),
.A2(n_1577),
.B(n_1579),
.C(n_1629),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1650),
.B(n_1586),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1651),
.B(n_1599),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1651),
.B(n_1604),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1655),
.A2(n_1577),
.B(n_1595),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1655),
.B(n_1602),
.C(n_1605),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1652),
.B(n_1620),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1638),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1649),
.B(n_1596),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1656),
.B(n_1621),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1645),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1648),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1664),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1682),
.B(n_1658),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1674),
.B(n_1649),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1666),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1688),
.A2(n_1670),
.B1(n_1657),
.B2(n_1663),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1674),
.B(n_1637),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1683),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1683),
.B(n_1632),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1687),
.A2(n_1603),
.B1(n_1609),
.B2(n_1640),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1675),
.B(n_1652),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1670),
.A2(n_1640),
.B(n_1657),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1693),
.B(n_1601),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1686),
.B(n_1637),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1666),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1632),
.Y(n_1710)
);

AND2x4_ASAP7_75t_SL g1711 ( 
.A(n_1693),
.B(n_1689),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1664),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1665),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1672),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1682),
.B(n_1658),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1666),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1673),
.B(n_1638),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1684),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1684),
.B(n_1638),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1675),
.B(n_1646),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1673),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1639),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1673),
.B(n_1639),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1678),
.B(n_1661),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1671),
.B(n_1643),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1678),
.B(n_1639),
.Y(n_1727)
);

AND2x4_ASAP7_75t_SL g1728 ( 
.A(n_1693),
.B(n_1653),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1690),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1678),
.B(n_1639),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1690),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1676),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1679),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_1699),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1719),
.B(n_1671),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1698),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1719),
.B(n_1671),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1719),
.B(n_1662),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1728),
.B(n_1662),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1698),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1701),
.B(n_1677),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1728),
.B(n_1662),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1709),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1687),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_1708),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1709),
.Y(n_1746)
);

AOI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1703),
.A2(n_1663),
.B(n_1688),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1728),
.B(n_1668),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1705),
.B(n_1693),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1704),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1700),
.B(n_1685),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1695),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1713),
.A2(n_1693),
.B(n_1560),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1704),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1725),
.B(n_1668),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1701),
.B(n_1677),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1708),
.B(n_1685),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1695),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1717),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1717),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1725),
.B(n_1668),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1725),
.B(n_1661),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1705),
.B(n_1676),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1722),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1695),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1697),
.B(n_1676),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1697),
.B(n_1694),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1707),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1711),
.B(n_1661),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1722),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1706),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1702),
.B(n_1680),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1732),
.Y(n_1773)
);

OAI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1733),
.A2(n_1681),
.B(n_1669),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1706),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1732),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1729),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1711),
.B(n_1672),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1696),
.B(n_1672),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1745),
.B(n_1702),
.Y(n_1780)
);

NOR2x1_ASAP7_75t_SL g1781 ( 
.A(n_1744),
.B(n_1693),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1736),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1745),
.B(n_1716),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1736),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1735),
.B(n_1720),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1754),
.B(n_1704),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1531),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1751),
.B(n_1716),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1741),
.B(n_1733),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1747),
.B(n_1707),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1735),
.B(n_1737),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1740),
.Y(n_1792)
);

AND2x4_ASAP7_75t_SL g1793 ( 
.A(n_1754),
.B(n_1721),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1754),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1737),
.B(n_1720),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1740),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1754),
.B(n_1720),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1756),
.B(n_1696),
.Y(n_1799)
);

OAI222xp33_ASAP7_75t_L g1800 ( 
.A1(n_1744),
.A2(n_1730),
.B1(n_1727),
.B2(n_1723),
.C1(n_1631),
.C2(n_1657),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1769),
.B(n_1723),
.Y(n_1802)
);

OAI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1774),
.A2(n_1681),
.B(n_1713),
.C(n_1679),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1769),
.B(n_1723),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1756),
.B(n_1696),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1746),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1751),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1746),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1734),
.B(n_1715),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1759),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1759),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1734),
.B(n_1715),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1738),
.B(n_1727),
.Y(n_1814)
);

AND4x1_ASAP7_75t_L g1815 ( 
.A(n_1749),
.B(n_1615),
.C(n_1612),
.D(n_1659),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1760),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1803),
.A2(n_1744),
.B1(n_1747),
.B2(n_1774),
.Y(n_1817)
);

XOR2x2_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1781),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1781),
.B(n_1794),
.Y(n_1819)
);

AOI322xp5_ASAP7_75t_L g1820 ( 
.A1(n_1810),
.A2(n_1762),
.A3(n_1727),
.B1(n_1730),
.B2(n_1763),
.C1(n_1642),
.C2(n_1744),
.Y(n_1820)
);

OAI321xp33_ASAP7_75t_L g1821 ( 
.A1(n_1813),
.A2(n_1744),
.A3(n_1763),
.B1(n_1762),
.B2(n_1679),
.C(n_1777),
.Y(n_1821)
);

OAI322xp33_ASAP7_75t_L g1822 ( 
.A1(n_1789),
.A2(n_1768),
.A3(n_1757),
.B1(n_1753),
.B2(n_1777),
.C1(n_1726),
.C2(n_1767),
.Y(n_1822)
);

O2A1O1Ixp5_ASAP7_75t_L g1823 ( 
.A1(n_1790),
.A2(n_1766),
.B(n_1767),
.C(n_1776),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1799),
.A2(n_1768),
.B1(n_1753),
.B2(n_1757),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1808),
.Y(n_1825)
);

CKINVDCx20_ASAP7_75t_R g1826 ( 
.A(n_1794),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1806),
.B(n_1715),
.Y(n_1827)
);

AOI322xp5_ASAP7_75t_L g1828 ( 
.A1(n_1785),
.A2(n_1730),
.A3(n_1642),
.B1(n_1729),
.B2(n_1731),
.C1(n_1692),
.C2(n_1755),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1782),
.Y(n_1829)
);

AOI21xp33_ASAP7_75t_SL g1830 ( 
.A1(n_1783),
.A2(n_1476),
.B(n_1778),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1800),
.A2(n_1731),
.B(n_1766),
.C(n_1772),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1786),
.B(n_1750),
.Y(n_1832)
);

AOI322xp5_ASAP7_75t_L g1833 ( 
.A1(n_1785),
.A2(n_1642),
.A3(n_1692),
.B1(n_1755),
.B2(n_1761),
.C1(n_1665),
.C2(n_1669),
.Y(n_1833)
);

A2O1A1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1780),
.A2(n_1642),
.B(n_1691),
.C(n_1660),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1793),
.A2(n_1691),
.B(n_1663),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1782),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1793),
.A2(n_1778),
.B(n_1742),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1798),
.B(n_1750),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1791),
.B(n_1761),
.Y(n_1839)
);

CKINVDCx14_ASAP7_75t_R g1840 ( 
.A(n_1791),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1783),
.B(n_1710),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1798),
.B(n_1739),
.Y(n_1842)
);

AO32x1_ASAP7_75t_L g1843 ( 
.A1(n_1805),
.A2(n_1742),
.A3(n_1739),
.B1(n_1748),
.B2(n_1779),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1784),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1840),
.B(n_1802),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1842),
.B(n_1795),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1826),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1821),
.A2(n_1817),
.B(n_1823),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1829),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1821),
.B(n_1786),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1825),
.B(n_1802),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1824),
.A2(n_1663),
.B1(n_1804),
.B2(n_1795),
.Y(n_1852)
);

O2A1O1Ixp5_ASAP7_75t_SL g1853 ( 
.A1(n_1832),
.A2(n_1816),
.B(n_1792),
.C(n_1796),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1822),
.B(n_1786),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1818),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1839),
.B(n_1804),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1819),
.B(n_1814),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1820),
.B(n_1805),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1841),
.B(n_1814),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1843),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1843),
.Y(n_1861)
);

OAI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1827),
.A2(n_1780),
.B1(n_1788),
.B2(n_1667),
.Y(n_1862)
);

AOI21xp33_ASAP7_75t_L g1863 ( 
.A1(n_1831),
.A2(n_1844),
.B(n_1836),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_SL g1864 ( 
.A(n_1838),
.B(n_1792),
.C(n_1784),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1834),
.A2(n_1788),
.B1(n_1830),
.B2(n_1837),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1847),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1851),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1848),
.A2(n_1835),
.B(n_1797),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1847),
.Y(n_1869)
);

XNOR2x1_ASAP7_75t_L g1870 ( 
.A(n_1855),
.B(n_1571),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1859),
.B(n_1858),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1856),
.B(n_1833),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1849),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1846),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1860),
.B(n_1861),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1854),
.A2(n_1726),
.B1(n_1750),
.B2(n_1779),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1866),
.B(n_1850),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1866),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1876),
.A2(n_1863),
.B1(n_1871),
.B2(n_1872),
.C(n_1860),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1868),
.B(n_1853),
.C(n_1864),
.Y(n_1881)
);

AOI221x1_ASAP7_75t_L g1882 ( 
.A1(n_1876),
.A2(n_1861),
.B1(n_1854),
.B2(n_1850),
.C(n_1865),
.Y(n_1882)
);

NAND4xp25_ASAP7_75t_L g1883 ( 
.A(n_1877),
.B(n_1852),
.C(n_1857),
.D(n_1828),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1869),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1869),
.B(n_1815),
.Y(n_1885)
);

AOI211xp5_ASAP7_75t_L g1886 ( 
.A1(n_1875),
.A2(n_1862),
.B(n_1796),
.C(n_1816),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1874),
.Y(n_1887)
);

OAI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1881),
.A2(n_1868),
.B1(n_1870),
.B2(n_1873),
.C(n_1867),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_R g1889 ( 
.A(n_1887),
.B(n_1645),
.Y(n_1889)
);

AOI221x1_ASAP7_75t_L g1890 ( 
.A1(n_1879),
.A2(n_1811),
.B1(n_1807),
.B2(n_1797),
.C(n_1812),
.Y(n_1890)
);

OAI211xp5_ASAP7_75t_L g1891 ( 
.A1(n_1882),
.A2(n_1868),
.B(n_1843),
.C(n_1750),
.Y(n_1891)
);

OAI211xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1880),
.A2(n_1862),
.B(n_1812),
.C(n_1811),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1878),
.A2(n_1884),
.B1(n_1879),
.B2(n_1883),
.C(n_1886),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1891),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1888),
.A2(n_1885),
.B1(n_1809),
.B2(n_1807),
.C(n_1801),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1893),
.A2(n_1809),
.B(n_1750),
.C(n_1748),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1892),
.A2(n_1750),
.B1(n_1760),
.B2(n_1773),
.C(n_1770),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_L g1898 ( 
.A(n_1890),
.B(n_1758),
.C(n_1752),
.Y(n_1898)
);

OAI221xp5_ASAP7_75t_L g1899 ( 
.A1(n_1889),
.A2(n_1758),
.B1(n_1775),
.B2(n_1752),
.C(n_1771),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1898),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1896),
.B(n_1645),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1894),
.B(n_1772),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1897),
.B(n_1714),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1899),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1900),
.B(n_1895),
.C(n_1758),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1901),
.B(n_1645),
.Y(n_1906)
);

XNOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1902),
.B(n_1566),
.Y(n_1907)
);

AOI222xp33_ASAP7_75t_L g1908 ( 
.A1(n_1905),
.A2(n_1904),
.B1(n_1903),
.B2(n_1765),
.C1(n_1775),
.C2(n_1752),
.Y(n_1908)
);

AO22x2_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1906),
.B1(n_1907),
.B2(n_1765),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_SL g1910 ( 
.A1(n_1909),
.A2(n_1524),
.B1(n_1570),
.B2(n_1773),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1909),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1911),
.B(n_1765),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1910),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1912),
.A2(n_1775),
.B(n_1771),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1913),
.B(n_1771),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1724),
.B(n_1718),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1914),
.B(n_1712),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1917),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_R g1919 ( 
.A1(n_1918),
.A2(n_1582),
.B1(n_1770),
.B2(n_1764),
.C(n_1776),
.Y(n_1919)
);

AOI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1919),
.A2(n_1524),
.B(n_1560),
.C(n_1764),
.Y(n_1920)
);


endmodule