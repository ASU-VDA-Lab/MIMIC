module real_aes_4816_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_1086, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_1088, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_1087, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_1086;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_1088;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_1087;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_1021;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_960;
wire n_1081;
wire n_1084;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_1014;
wire n_366;
wire n_346;
wire n_1083;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_0), .A2(n_688), .B(n_690), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_1), .A2(n_148), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g446 ( .A(n_2), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_3), .A2(n_127), .B1(n_408), .B2(n_523), .Y(n_598) );
INVx1_ASAP7_75t_L g391 ( .A(n_4), .Y(n_391) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_5), .Y(n_309) );
AND2x4_ASAP7_75t_L g838 ( .A(n_5), .B(n_290), .Y(n_838) );
AND2x4_ASAP7_75t_L g843 ( .A(n_5), .B(n_844), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_6), .A2(n_7), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI221x1_ASAP7_75t_L g771 ( .A1(n_8), .A2(n_80), .B1(n_529), .B2(n_591), .C(n_772), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_9), .A2(n_241), .B1(n_483), .B2(n_492), .Y(n_737) );
AO22x1_ASAP7_75t_L g864 ( .A1(n_10), .A2(n_16), .B1(n_839), .B2(n_849), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_11), .A2(n_69), .B1(n_512), .B2(n_513), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_12), .A2(n_254), .B1(n_490), .B2(n_496), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_13), .A2(n_63), .B1(n_417), .B2(n_419), .Y(n_416) );
XNOR2x1_ASAP7_75t_L g579 ( .A(n_14), .B(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_14), .A2(n_213), .B1(n_842), .B2(n_845), .Y(n_841) );
INVx1_ASAP7_75t_L g804 ( .A(n_15), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_17), .A2(n_210), .B1(n_442), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_18), .A2(n_41), .B1(n_492), .B2(n_493), .Y(n_615) );
INVx1_ASAP7_75t_L g754 ( .A(n_19), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_20), .A2(n_281), .B1(n_570), .B2(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g750 ( .A(n_21), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_22), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_23), .A2(n_230), .B1(n_417), .B2(n_513), .Y(n_820) );
AO22x1_ASAP7_75t_L g649 ( .A1(n_24), .A2(n_135), .B1(n_515), .B2(n_636), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_25), .A2(n_110), .B1(n_459), .B2(n_460), .Y(n_1067) );
XNOR2xp5_ASAP7_75t_L g1079 ( .A(n_26), .B(n_1080), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_27), .A2(n_137), .B1(n_862), .B2(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_28), .A2(n_200), .B1(n_375), .B2(n_448), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_29), .A2(n_99), .B1(n_483), .B2(n_504), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_30), .A2(n_251), .B1(n_519), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_31), .A2(n_92), .B1(n_489), .B2(n_492), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_32), .A2(n_280), .B1(n_630), .B2(n_631), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_33), .A2(n_108), .B1(n_424), .B2(n_683), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_34), .A2(n_273), .B1(n_349), .B2(n_610), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_35), .A2(n_93), .B1(n_420), .B2(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_36), .A2(n_181), .B1(n_442), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_37), .A2(n_161), .B1(n_592), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g717 ( .A(n_38), .Y(n_717) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_39), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_40), .A2(n_155), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_42), .A2(n_250), .B1(n_483), .B2(n_484), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_43), .B(n_633), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_44), .A2(n_71), .B1(n_420), .B2(n_467), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_45), .A2(n_172), .B1(n_462), .B2(n_464), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_46), .A2(n_84), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_47), .A2(n_95), .B1(n_470), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_48), .A2(n_295), .B1(n_442), .B2(n_658), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_49), .B(n_219), .Y(n_307) );
INVx1_ASAP7_75t_L g345 ( .A(n_49), .Y(n_345) );
INVxp67_ASAP7_75t_L g358 ( .A(n_49), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_50), .A2(n_144), .B1(n_842), .B2(n_845), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_51), .A2(n_238), .B1(n_515), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_52), .A2(n_167), .B1(n_484), .B2(n_493), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_53), .A2(n_259), .B1(n_565), .B2(n_567), .Y(n_564) );
INVx1_ASAP7_75t_L g450 ( .A(n_54), .Y(n_450) );
INVx1_ASAP7_75t_L g508 ( .A(n_55), .Y(n_508) );
INVx1_ASAP7_75t_L g662 ( .A(n_56), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_57), .A2(n_235), .B1(n_417), .B2(n_419), .Y(n_679) );
INVx1_ASAP7_75t_L g805 ( .A(n_58), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_59), .B(n_330), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_60), .A2(n_81), .B1(n_417), .B2(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g437 ( .A(n_61), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_62), .A2(n_179), .B1(n_439), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_64), .A2(n_263), .B1(n_501), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_65), .A2(n_180), .B1(n_399), .B2(n_404), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_66), .A2(n_190), .B1(n_835), .B2(n_839), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_67), .A2(n_292), .B1(n_404), .B2(n_414), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_68), .A2(n_113), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g304 ( .A(n_70), .Y(n_304) );
INVx1_ASAP7_75t_L g837 ( .A(n_72), .Y(n_837) );
AND2x4_ASAP7_75t_L g840 ( .A(n_72), .B(n_304), .Y(n_840) );
INVx1_ASAP7_75t_SL g871 ( .A(n_72), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_73), .A2(n_203), .B1(n_448), .B2(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_74), .A2(n_279), .B1(n_459), .B2(n_460), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_75), .A2(n_142), .B1(n_486), .B2(n_487), .Y(n_613) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_76), .A2(n_138), .B1(n_549), .B2(n_551), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_77), .B(n_555), .Y(n_664) );
INVx1_ASAP7_75t_L g444 ( .A(n_78), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_79), .A2(n_201), .B1(n_849), .B2(n_893), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_82), .A2(n_224), .B1(n_399), .B2(n_404), .Y(n_681) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_83), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_85), .A2(n_123), .B1(n_462), .B2(n_653), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_86), .A2(n_236), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g696 ( .A(n_87), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_88), .B(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_89), .A2(n_96), .B1(n_600), .B2(n_760), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_90), .A2(n_91), .B1(n_408), .B2(n_414), .Y(n_823) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_94), .B(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_94), .A2(n_177), .B1(n_842), .B2(n_860), .Y(n_859) );
INVx1_ASAP7_75t_SL g770 ( .A(n_97), .Y(n_770) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_97), .B(n_797), .C(n_798), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_98), .A2(n_130), .B1(n_349), .B2(n_360), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_100), .B(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g1060 ( .A1(n_101), .A2(n_157), .B1(n_526), .B2(n_547), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_102), .A2(n_212), .B1(n_835), .B2(n_839), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_103), .A2(n_193), .B1(n_839), .B2(n_849), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_104), .A2(n_229), .B1(n_486), .B2(n_487), .Y(n_738) );
INVx1_ASAP7_75t_L g331 ( .A(n_105), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_105), .B(n_217), .Y(n_355) );
AOI33xp33_ASAP7_75t_R g640 ( .A1(n_106), .A2(n_247), .A3(n_327), .B1(n_383), .B2(n_641), .B3(n_1086), .Y(n_640) );
INVx1_ASAP7_75t_L g440 ( .A(n_107), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_109), .A2(n_205), .B1(n_512), .B2(n_513), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_111), .A2(n_153), .B1(n_460), .B2(n_522), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_112), .A2(n_262), .B1(n_512), .B2(n_572), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_114), .A2(n_121), .B1(n_496), .B2(n_502), .Y(n_731) );
INVx1_ASAP7_75t_L g727 ( .A(n_115), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_116), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_117), .A2(n_226), .B1(n_459), .B2(n_460), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_118), .A2(n_221), .B1(n_489), .B2(n_490), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_119), .A2(n_283), .B1(n_408), .B2(n_414), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_120), .A2(n_132), .B1(n_842), .B2(n_845), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_122), .A2(n_184), .B1(n_842), .B2(n_890), .Y(n_889) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_124), .A2(n_501), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g506 ( .A(n_125), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g503 ( .A1(n_126), .A2(n_504), .B(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_128), .A2(n_284), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_129), .A2(n_150), .B1(n_490), .B2(n_493), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_131), .A2(n_242), .B1(n_424), .B2(n_576), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_133), .A2(n_166), .B1(n_452), .B2(n_504), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_134), .A2(n_169), .B1(n_439), .B2(n_448), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_136), .A2(n_222), .B1(n_890), .B2(n_919), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_139), .A2(n_253), .B1(n_408), .B2(n_414), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_140), .A2(n_202), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_141), .A2(n_170), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g386 ( .A(n_143), .Y(n_386) );
XNOR2x1_ASAP7_75t_L g540 ( .A(n_144), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_145), .A2(n_186), .B1(n_544), .B2(n_545), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_146), .A2(n_160), .B1(n_486), .B2(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_147), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g809 ( .A(n_149), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_151), .A2(n_261), .B1(n_591), .B2(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_152), .B(n_694), .Y(n_1061) );
INVx1_ASAP7_75t_L g691 ( .A(n_154), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_156), .A2(n_174), .B1(n_462), .B2(n_520), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_158), .A2(n_272), .B1(n_484), .B2(n_489), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_159), .A2(n_162), .B1(n_587), .B2(n_589), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_163), .A2(n_187), .B1(n_562), .B2(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_164), .B(n_583), .Y(n_582) );
XOR2xp5_ASAP7_75t_L g603 ( .A(n_165), .B(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_165), .A2(n_269), .B1(n_845), .B2(n_870), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_168), .A2(n_268), .B1(n_526), .B2(n_631), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_171), .A2(n_215), .B1(n_325), .B2(n_1064), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_173), .A2(n_232), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_175), .A2(n_188), .B1(n_452), .B2(n_502), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_176), .A2(n_257), .B1(n_388), .B2(n_529), .C(n_531), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_178), .A2(n_183), .B1(n_399), .B2(n_404), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_182), .A2(n_231), .B1(n_835), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_185), .A2(n_196), .B1(n_375), .B2(n_448), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_189), .A2(n_220), .B1(n_442), .B2(n_628), .Y(n_627) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_191), .A2(n_554), .B(n_556), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_192), .B(n_631), .Y(n_692) );
AO221x2_ASAP7_75t_L g863 ( .A1(n_194), .A2(n_246), .B1(n_842), .B2(n_860), .C(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g1070 ( .A(n_194), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_194), .A2(n_1077), .B1(n_1079), .B2(n_1081), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_195), .A2(n_282), .B1(n_512), .B2(n_513), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_197), .A2(n_296), .B1(n_424), .B2(n_683), .Y(n_682) );
OA22x2_ASAP7_75t_L g335 ( .A1(n_198), .A2(n_219), .B1(n_330), .B2(n_334), .Y(n_335) );
INVx1_ASAP7_75t_L g370 ( .A(n_198), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_199), .A2(n_206), .B1(n_499), .B2(n_631), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_204), .A2(n_287), .B1(n_835), .B2(n_893), .Y(n_892) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_207), .Y(n_783) );
AO22x2_ASAP7_75t_L g431 ( .A1(n_208), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_208), .Y(n_432) );
AND2x2_ASAP7_75t_L g772 ( .A(n_209), .B(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_211), .A2(n_274), .B1(n_683), .B2(n_757), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_214), .A2(n_248), .B1(n_404), .B2(n_515), .Y(n_1066) );
CKINVDCx6p67_ASAP7_75t_R g800 ( .A(n_216), .Y(n_800) );
INVx1_ASAP7_75t_L g347 ( .A(n_217), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_217), .B(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_218), .A2(n_243), .B1(n_501), .B2(n_502), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g384 ( .A1(n_219), .A2(n_237), .B(n_359), .Y(n_384) );
XNOR2x1_ASAP7_75t_L g479 ( .A(n_223), .B(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_225), .A2(n_255), .B1(n_470), .B2(n_483), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_227), .B(n_375), .Y(n_606) );
INVx1_ASAP7_75t_L g702 ( .A(n_228), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_233), .A2(n_245), .B1(n_399), .B2(n_597), .Y(n_596) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_234), .A2(n_645), .B(n_665), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_234), .B(n_648), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_237), .B(n_278), .Y(n_308) );
INVx1_ASAP7_75t_L g333 ( .A(n_237), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_239), .A2(n_265), .B1(n_459), .B2(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_240), .B(n_501), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_244), .A2(n_260), .B1(n_399), .B2(n_424), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_249), .A2(n_256), .B1(n_515), .B2(n_516), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_252), .Y(n_317) );
INVx1_ASAP7_75t_L g813 ( .A(n_258), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_264), .A2(n_294), .B1(n_360), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_266), .A2(n_285), .B1(n_388), .B2(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g748 ( .A(n_267), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_270), .Y(n_752) );
INVx1_ASAP7_75t_L g557 ( .A(n_271), .Y(n_557) );
INVx1_ASAP7_75t_L g815 ( .A(n_275), .Y(n_815) );
INVx1_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
INVx1_ASAP7_75t_L g372 ( .A(n_277), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_278), .B(n_340), .Y(n_339) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_286), .A2(n_388), .B(n_661), .Y(n_660) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_288), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_289), .Y(n_743) );
INVx1_ASAP7_75t_L g844 ( .A(n_290), .Y(n_844) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_290), .Y(n_1083) );
INVx1_ASAP7_75t_L g532 ( .A(n_291), .Y(n_532) );
INVx1_ASAP7_75t_L g379 ( .A(n_293), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_310), .B(n_827), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .C(n_309), .Y(n_301) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_302), .B(n_1074), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_302), .B(n_1075), .Y(n_1078) );
AOI21xp5_ASAP7_75t_L g1084 ( .A1(n_302), .A2(n_309), .B(n_871), .Y(n_1084) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AO21x1_ASAP7_75t_L g1082 ( .A1(n_303), .A2(n_1083), .B(n_1084), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g836 ( .A(n_304), .B(n_837), .Y(n_836) );
AND3x4_ASAP7_75t_L g870 ( .A(n_304), .B(n_843), .C(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_305), .B(n_1075), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_306), .A2(n_364), .B(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g1075 ( .A(n_309), .Y(n_1075) );
XNOR2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_618), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_537), .B2(n_538), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_476), .B1(n_534), .B2(n_536), .Y(n_313) );
INVx1_ASAP7_75t_L g536 ( .A(n_314), .Y(n_536) );
OA22x2_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_429), .B1(n_473), .B2(n_474), .Y(n_314) );
INVx4_ASAP7_75t_R g315 ( .A(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g473 ( .A(n_316), .Y(n_473) );
XNOR2x1_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_397), .Y(n_318) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_371), .C(n_385), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_348), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_324), .A2(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g530 ( .A(n_326), .Y(n_530) );
INVx2_ASAP7_75t_L g585 ( .A(n_326), .Y(n_585) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_336), .Y(n_326) );
AND2x2_ASAP7_75t_L g396 ( .A(n_327), .B(n_390), .Y(n_396) );
AND2x4_ASAP7_75t_L g400 ( .A(n_327), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g425 ( .A(n_327), .B(n_412), .Y(n_425) );
AND2x2_ASAP7_75t_L g463 ( .A(n_327), .B(n_412), .Y(n_463) );
AND2x4_ASAP7_75t_L g483 ( .A(n_327), .B(n_412), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_327), .B(n_406), .Y(n_484) );
AND2x4_ASAP7_75t_L g496 ( .A(n_327), .B(n_390), .Y(n_496) );
AND2x2_ASAP7_75t_L g501 ( .A(n_327), .B(n_336), .Y(n_501) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_335), .Y(n_327) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
NAND2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g334 ( .A(n_330), .Y(n_334) );
INVx3_ASAP7_75t_L g340 ( .A(n_330), .Y(n_340) );
NAND2xp33_ASAP7_75t_L g346 ( .A(n_330), .B(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_330), .Y(n_354) );
INVx1_ASAP7_75t_L g359 ( .A(n_330), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_331), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_333), .A2(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g356 ( .A(n_335), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g377 ( .A(n_335), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g411 ( .A(n_335), .Y(n_411) );
AND2x4_ASAP7_75t_L g376 ( .A(n_336), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g382 ( .A(n_336), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g422 ( .A(n_336), .B(n_410), .Y(n_422) );
AND2x4_ASAP7_75t_L g487 ( .A(n_336), .B(n_410), .Y(n_487) );
AND2x2_ASAP7_75t_L g499 ( .A(n_336), .B(n_377), .Y(n_499) );
AND2x4_ASAP7_75t_L g502 ( .A(n_336), .B(n_383), .Y(n_502) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_342), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g352 ( .A(n_338), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g390 ( .A(n_338), .B(n_342), .Y(n_390) );
OR2x2_ASAP7_75t_L g402 ( .A(n_338), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g412 ( .A(n_338), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
NAND3xp33_ASAP7_75t_L g365 ( .A(n_341), .B(n_366), .C(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g403 ( .A(n_343), .Y(n_403) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_350), .A2(n_557), .B(n_558), .Y(n_556) );
INVx4_ASAP7_75t_L g594 ( .A(n_350), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_350), .A2(n_691), .B(n_692), .Y(n_690) );
INVx5_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g526 ( .A(n_351), .Y(n_526) );
BUFx2_ASAP7_75t_L g628 ( .A(n_351), .Y(n_628) );
BUFx4f_ASAP7_75t_L g658 ( .A(n_351), .Y(n_658) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .Y(n_351) );
AND2x2_ASAP7_75t_L g452 ( .A(n_352), .B(n_356), .Y(n_452) );
AND2x4_ASAP7_75t_L g497 ( .A(n_352), .B(n_356), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g364 ( .A(n_354), .Y(n_364) );
INVx4_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g559 ( .A(n_361), .Y(n_559) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g774 ( .A(n_362), .Y(n_774) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_363), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_367), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g383 ( .A(n_368), .B(n_384), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_379), .B2(n_380), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g445 ( .A(n_375), .Y(n_445) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_376), .Y(n_550) );
BUFx8_ASAP7_75t_SL g591 ( .A(n_376), .Y(n_591) );
BUFx3_ASAP7_75t_L g633 ( .A(n_376), .Y(n_633) );
INVx2_ASAP7_75t_L g695 ( .A(n_376), .Y(n_695) );
INVx2_ASAP7_75t_L g812 ( .A(n_376), .Y(n_812) );
AND2x4_ASAP7_75t_L g389 ( .A(n_377), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g504 ( .A(n_377), .B(n_390), .Y(n_504) );
AND2x4_ASAP7_75t_L g410 ( .A(n_378), .B(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_380), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
INVx3_ASAP7_75t_L g552 ( .A(n_382), .Y(n_552) );
AND2x4_ASAP7_75t_L g405 ( .A(n_383), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g428 ( .A(n_383), .B(n_412), .Y(n_428) );
AND2x4_ASAP7_75t_L g492 ( .A(n_383), .B(n_412), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_383), .B(n_406), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_391), .B2(n_392), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_387), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
INVx4_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
INVx1_ASAP7_75t_L g588 ( .A(n_389), .Y(n_588) );
BUFx3_ASAP7_75t_L g713 ( .A(n_389), .Y(n_713) );
AND2x4_ASAP7_75t_L g418 ( .A(n_390), .B(n_410), .Y(n_418) );
AND2x4_ASAP7_75t_L g486 ( .A(n_390), .B(n_410), .Y(n_486) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g589 ( .A(n_394), .Y(n_589) );
INVx2_ASAP7_75t_L g686 ( .A(n_394), .Y(n_686) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g807 ( .A(n_395), .Y(n_807) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_396), .Y(n_442) );
BUFx3_ASAP7_75t_L g547 ( .A(n_396), .Y(n_547) );
AND4x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_407), .C(n_416), .D(n_423), .Y(n_397) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_400), .Y(n_470) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_400), .Y(n_515) );
BUFx12f_ASAP7_75t_L g568 ( .A(n_400), .Y(n_568) );
AND2x4_ASAP7_75t_L g490 ( .A(n_401), .B(n_410), .Y(n_490) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g406 ( .A(n_402), .Y(n_406) );
INVx1_ASAP7_75t_L g413 ( .A(n_403), .Y(n_413) );
BUFx12f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx6_ASAP7_75t_L g472 ( .A(n_405), .Y(n_472) );
AND2x4_ASAP7_75t_L g415 ( .A(n_406), .B(n_410), .Y(n_415) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx12f_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_409), .Y(n_522) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
AND2x4_ASAP7_75t_L g489 ( .A(n_410), .B(n_412), .Y(n_489) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_412), .Y(n_641) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_414), .Y(n_562) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_415), .Y(n_523) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_415), .Y(n_639) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g468 ( .A(n_418), .Y(n_468) );
BUFx12f_ASAP7_75t_L g512 ( .A(n_418), .Y(n_512) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_422), .Y(n_513) );
BUFx3_ASAP7_75t_L g572 ( .A(n_422), .Y(n_572) );
BUFx5_ASAP7_75t_L g600 ( .A(n_422), .Y(n_600) );
BUFx8_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_425), .Y(n_566) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx4_ASAP7_75t_L g464 ( .A(n_427), .Y(n_464) );
INVx2_ASAP7_75t_SL g520 ( .A(n_427), .Y(n_520) );
INVx1_ASAP7_75t_L g576 ( .A(n_427), .Y(n_576) );
INVx4_ASAP7_75t_L g653 ( .A(n_427), .Y(n_653) );
INVx4_ASAP7_75t_L g683 ( .A(n_427), .Y(n_683) );
INVx8_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g475 ( .A(n_431), .Y(n_475) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_456), .Y(n_434) );
NOR3xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_443), .C(n_449), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g544 ( .A(n_439), .Y(n_544) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_443) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_454), .B(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_455), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g610 ( .A(n_455), .Y(n_610) );
INVx2_ASAP7_75t_L g631 ( .A(n_455), .Y(n_631) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_455), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_465), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .Y(n_457) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_459), .Y(n_574) );
BUFx12f_ASAP7_75t_L g757 ( .A(n_459), .Y(n_757) );
BUFx4f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_463), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
BUFx4f_ASAP7_75t_L g760 ( .A(n_467), .Y(n_760) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g516 ( .A(n_472), .Y(n_516) );
INVx1_ASAP7_75t_L g597 ( .A(n_472), .Y(n_597) );
INVx5_ASAP7_75t_L g636 ( .A(n_472), .Y(n_636) );
INVx2_ASAP7_75t_L g706 ( .A(n_472), .Y(n_706) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g535 ( .A(n_477), .Y(n_535) );
AO22x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_507), .B2(n_533), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_494), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .C(n_488), .D(n_491), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .C(n_500), .D(n_503), .Y(n_494) );
INVx2_ASAP7_75t_L g791 ( .A(n_496), .Y(n_791) );
INVx4_ASAP7_75t_L g784 ( .A(n_497), .Y(n_784) );
INVx2_ASAP7_75t_L g786 ( .A(n_502), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_504), .Y(n_789) );
INVx1_ASAP7_75t_L g533 ( .A(n_507), .Y(n_533) );
XNOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
NAND4xp75_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .C(n_524), .D(n_528), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_512), .Y(n_570) );
BUFx2_ASAP7_75t_L g563 ( .A(n_516), .Y(n_563) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
INVx1_ASAP7_75t_L g689 ( .A(n_529), .Y(n_689) );
INVx1_ASAP7_75t_L g816 ( .A(n_529), .Y(n_816) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g555 ( .A(n_530), .Y(n_555) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
XOR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_577), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_560), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .C(n_553), .Y(n_542) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_546), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g592 ( .A(n_552), .Y(n_592) );
INVx2_ASAP7_75t_L g626 ( .A(n_552), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_552), .A2(n_809), .B1(n_810), .B2(n_813), .Y(n_808) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .C(n_569), .D(n_573), .Y(n_560) );
BUFx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AO22x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_602), .B1(n_616), .B2(n_617), .Y(n_578) );
INVx2_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_595), .Y(n_580) );
NAND4xp25_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .C(n_590), .D(n_593), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g745 ( .A(n_584), .Y(n_745) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g630 ( .A(n_585), .Y(n_630) );
INVx2_ASAP7_75t_L g753 ( .A(n_587), .Y(n_753) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .C(n_599), .D(n_601), .Y(n_595) );
INVx1_ASAP7_75t_L g617 ( .A(n_602), .Y(n_617) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_611), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .C(n_608), .D(n_609), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .C(n_614), .D(n_615), .Y(n_611) );
XOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_721), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_672), .B1(n_673), .B2(n_720), .Y(n_619) );
INVx1_ASAP7_75t_L g720 ( .A(n_620), .Y(n_720) );
AO22x2_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_642), .B1(n_643), .B2(n_669), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g671 ( .A(n_622), .Y(n_671) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_634), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .C(n_629), .D(n_632), .Y(n_624) );
INVx2_ASAP7_75t_L g749 ( .A(n_633), .Y(n_749) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .C(n_638), .D(n_640), .Y(n_634) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_654), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .C(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_649), .B(n_659), .C(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_650), .B(n_655), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_659), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_663), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g1064 ( .A(n_663), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_697), .B2(n_718), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
XOR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_696), .Y(n_676) );
NOR2x1_ASAP7_75t_L g677 ( .A(n_678), .B(n_684), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .C(n_681), .D(n_682), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .C(n_693), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g719 ( .A(n_698), .Y(n_719) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
XNOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .C(n_708), .D(n_709), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .C(n_714), .D(n_715), .Y(n_710) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_762), .B2(n_826), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
XNOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_739), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
XNOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
OR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_734), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .C(n_732), .D(n_733), .Y(n_729) );
NAND4xp25_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .C(n_737), .D(n_738), .Y(n_734) );
NAND2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_755), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_747), .C(n_751), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B(n_746), .Y(n_742) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND4x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .C(n_759), .D(n_761), .Y(n_755) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_763), .Y(n_826) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_764), .A2(n_765), .B1(n_799), .B2(n_825), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_792), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_775), .C(n_779), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_771), .B2(n_1087), .Y(n_768) );
INVx1_ASAP7_75t_L g797 ( .A(n_769), .Y(n_797) );
NOR2xp67_ASAP7_75t_L g775 ( .A(n_770), .B(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_770), .A2(n_780), .B1(n_781), .B2(n_1088), .Y(n_779) );
INVx1_ASAP7_75t_L g794 ( .A(n_771), .Y(n_794) );
INVx4_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_776), .B(n_793), .C(n_796), .Y(n_792) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g798 ( .A(n_780), .Y(n_798) );
INVx1_ASAP7_75t_L g795 ( .A(n_781), .Y(n_795) );
NOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_787), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_799), .Y(n_825) );
XNOR2x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
NAND2x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_818), .Y(n_801) );
NOR3xp33_ASAP7_75t_SL g802 ( .A(n_803), .B(n_808), .C(n_814), .Y(n_802) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B(n_817), .Y(n_814) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_1048), .B1(n_1050), .B2(n_1071), .C(n_1076), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_1006), .C(n_1030), .Y(n_828) );
AOI33xp33_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_894), .A3(n_922), .B1(n_959), .B2(n_984), .B3(n_997), .Y(n_829) );
A2O1A1Ixp33_ASAP7_75t_SL g830 ( .A1(n_831), .A2(n_851), .B(n_865), .C(n_887), .Y(n_830) );
AND2x2_ASAP7_75t_L g940 ( .A(n_831), .B(n_886), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_831), .B(n_885), .Y(n_1047) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_832), .A2(n_874), .B1(n_907), .B2(n_912), .C(n_916), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_832), .B(n_930), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_832), .B(n_993), .Y(n_992) );
OR2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_846), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_833), .B(n_852), .Y(n_879) );
INVx4_ASAP7_75t_L g902 ( .A(n_833), .Y(n_902) );
OR2x2_ASAP7_75t_L g905 ( .A(n_833), .B(n_847), .Y(n_905) );
AND2x2_ASAP7_75t_L g947 ( .A(n_833), .B(n_846), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_833), .B(n_852), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_833), .B(n_853), .Y(n_1039) );
AND2x2_ASAP7_75t_L g833 ( .A(n_834), .B(n_841), .Y(n_833) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_838), .Y(n_835) );
AND2x4_ASAP7_75t_L g842 ( .A(n_836), .B(n_843), .Y(n_842) );
AND2x4_ASAP7_75t_L g849 ( .A(n_836), .B(n_838), .Y(n_849) );
AND2x2_ASAP7_75t_L g873 ( .A(n_836), .B(n_838), .Y(n_873) );
AND2x2_ASAP7_75t_L g839 ( .A(n_838), .B(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g862 ( .A(n_838), .B(n_840), .Y(n_862) );
AND2x4_ASAP7_75t_L g893 ( .A(n_838), .B(n_840), .Y(n_893) );
AND2x4_ASAP7_75t_L g845 ( .A(n_840), .B(n_843), .Y(n_845) );
AND2x4_ASAP7_75t_L g860 ( .A(n_840), .B(n_843), .Y(n_860) );
INVx3_ASAP7_75t_L g920 ( .A(n_842), .Y(n_920) );
INVx2_ASAP7_75t_SL g891 ( .A(n_845), .Y(n_891) );
INVx2_ASAP7_75t_L g874 ( .A(n_846), .Y(n_874) );
OR2x2_ASAP7_75t_L g938 ( .A(n_846), .B(n_902), .Y(n_938) );
INVxp67_ASAP7_75t_L g969 ( .A(n_846), .Y(n_969) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_846), .B(n_962), .Y(n_1022) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_847), .B(n_888), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
AND2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_856), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_852), .B(n_857), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_852), .B(n_944), .Y(n_943) );
A2O1A1Ixp33_ASAP7_75t_L g954 ( .A1(n_852), .A2(n_876), .B(n_955), .C(n_957), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g1005 ( .A(n_852), .B(n_900), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_852), .B(n_903), .Y(n_1028) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx3_ASAP7_75t_L g886 ( .A(n_853), .Y(n_886) );
INVx2_ASAP7_75t_L g910 ( .A(n_853), .Y(n_910) );
AND2x2_ASAP7_75t_L g915 ( .A(n_853), .B(n_857), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_853), .B(n_949), .Y(n_967) );
AOI321xp33_ASAP7_75t_L g997 ( .A1(n_853), .A2(n_874), .A3(n_881), .B1(n_998), .B2(n_1001), .C(n_1002), .Y(n_997) );
AND2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
AND2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_863), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_857), .B(n_877), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_857), .B(n_933), .Y(n_932) );
AND2x2_ASAP7_75t_L g980 ( .A(n_857), .B(n_882), .Y(n_980) );
AND2x2_ASAP7_75t_L g987 ( .A(n_857), .B(n_914), .Y(n_987) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_857), .B(n_867), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_857), .B(n_895), .Y(n_1014) );
A2O1A1Ixp33_ASAP7_75t_SL g1023 ( .A1(n_857), .A2(n_1024), .B(n_1028), .C(n_1029), .Y(n_1023) );
CKINVDCx6p67_ASAP7_75t_R g857 ( .A(n_858), .Y(n_857) );
AND2x2_ASAP7_75t_L g876 ( .A(n_858), .B(n_877), .Y(n_876) );
AND2x2_ASAP7_75t_L g884 ( .A(n_858), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g903 ( .A(n_858), .B(n_882), .Y(n_903) );
AND2x2_ASAP7_75t_L g923 ( .A(n_858), .B(n_924), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_858), .B(n_877), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_858), .B(n_863), .Y(n_949) );
AND2x2_ASAP7_75t_L g951 ( .A(n_858), .B(n_867), .Y(n_951) );
AND2x2_ASAP7_75t_L g964 ( .A(n_858), .B(n_933), .Y(n_964) );
AND2x2_ASAP7_75t_L g975 ( .A(n_858), .B(n_914), .Y(n_975) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_858), .B(n_868), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_858), .B(n_934), .Y(n_1017) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_861), .Y(n_858) );
AND2x2_ASAP7_75t_L g867 ( .A(n_863), .B(n_868), .Y(n_867) );
OR2x2_ASAP7_75t_L g883 ( .A(n_863), .B(n_868), .Y(n_883) );
AND2x2_ASAP7_75t_L g914 ( .A(n_863), .B(n_877), .Y(n_914) );
INVx1_ASAP7_75t_L g934 ( .A(n_863), .Y(n_934) );
OAI321xp33_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_867), .A3(n_874), .B1(n_875), .B2(n_878), .C(n_880), .Y(n_865) );
AND2x2_ASAP7_75t_L g924 ( .A(n_867), .B(n_886), .Y(n_924) );
INVx1_ASAP7_75t_L g981 ( .A(n_867), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_867), .B(n_884), .Y(n_1046) );
INVx1_ASAP7_75t_L g877 ( .A(n_868), .Y(n_877) );
AND2x2_ASAP7_75t_L g933 ( .A(n_868), .B(n_934), .Y(n_933) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .Y(n_868) );
INVx3_ASAP7_75t_SL g946 ( .A(n_874), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_874), .B(n_962), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_874), .B(n_1003), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_874), .A2(n_1001), .B1(n_1016), .B2(n_1018), .C(n_1020), .Y(n_1015) );
NAND2xp5_ASAP7_75t_SL g998 ( .A(n_875), .B(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_876), .B(n_940), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_876), .A2(n_916), .B1(n_967), .B2(n_968), .C(n_970), .Y(n_966) );
INVxp67_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_881), .B(n_925), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_881), .B(n_1035), .Y(n_1034) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_884), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR2x1_ASAP7_75t_L g895 ( .A(n_883), .B(n_885), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_885), .B(n_933), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g970 ( .A(n_885), .B(n_971), .Y(n_970) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_885), .B(n_931), .Y(n_1032) );
INVx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_886), .B(n_987), .Y(n_986) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_887), .A2(n_942), .B1(n_950), .B2(n_952), .C(n_954), .Y(n_941) );
OAI211xp5_ASAP7_75t_L g1006 ( .A1(n_887), .A2(n_1007), .B(n_1015), .C(n_1023), .Y(n_1006) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
AND2x2_ASAP7_75t_L g936 ( .A(n_888), .B(n_937), .Y(n_936) );
AND2x2_ASAP7_75t_L g953 ( .A(n_888), .B(n_908), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_888), .B(n_926), .Y(n_958) );
INVx4_ASAP7_75t_L g962 ( .A(n_888), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_888), .B(n_938), .Y(n_996) );
AND2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_892), .Y(n_888) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_896), .B1(n_903), .B2(n_904), .C(n_906), .Y(n_894) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_898), .Y(n_1013) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_900), .Y(n_1035) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g926 ( .A(n_901), .Y(n_926) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g908 ( .A(n_902), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_903), .B(n_936), .Y(n_989) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_905), .B(n_910), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_905), .B(n_962), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_910), .B(n_929), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_910), .B(n_964), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_910), .B(n_1004), .Y(n_1011) );
INVx1_ASAP7_75t_L g929 ( .A(n_911), .Y(n_929) );
INVxp67_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g1027 ( .A(n_914), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_916), .B(n_962), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_921), .Y(n_917) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_919), .Y(n_1049) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AOI211xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_925), .B(n_927), .C(n_941), .Y(n_922) );
INVx1_ASAP7_75t_L g991 ( .A(n_924), .Y(n_991) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_925), .B(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
A2O1A1Ixp33_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_930), .B(n_935), .C(n_939), .Y(n_927) );
INVx1_ASAP7_75t_L g994 ( .A(n_929), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_930), .A2(n_1043), .B1(n_1046), .B2(n_1047), .Y(n_1042) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g1026 ( .A(n_933), .Y(n_1026) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
O2A1O1Ixp33_ASAP7_75t_L g1036 ( .A1(n_940), .A2(n_1037), .B(n_1040), .C(n_1042), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_942) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g971 ( .A(n_947), .Y(n_971) );
O2A1O1Ixp33_ASAP7_75t_SL g1007 ( .A1(n_947), .A2(n_980), .B(n_1008), .C(n_1012), .Y(n_1007) );
INVxp67_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
AOI21xp33_ASAP7_75t_L g1020 ( .A1(n_950), .A2(n_1003), .B(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
AOI211xp5_ASAP7_75t_L g984 ( .A1(n_957), .A2(n_985), .B(n_988), .C(n_990), .Y(n_984) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
NOR4xp25_ASAP7_75t_L g959 ( .A(n_960), .B(n_965), .C(n_977), .D(n_978), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_963), .Y(n_960) );
INVx1_ASAP7_75t_L g1001 ( .A(n_961), .Y(n_1001) );
INVx2_ASAP7_75t_L g993 ( .A(n_962), .Y(n_993) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_962), .B(n_969), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_964), .B(n_980), .Y(n_1041) );
AOI21xp33_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_972), .B(n_976), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_967), .B(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_975), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
AOI21xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_981), .B(n_982), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVxp67_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVxp67_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B1(n_994), .B2(n_995), .Y(n_990) );
OAI221xp5_ASAP7_75t_L g1030 ( .A1(n_993), .A2(n_1031), .B1(n_1033), .B2(n_1034), .C(n_1036), .Y(n_1030) );
NOR2xp33_ASAP7_75t_L g1037 ( .A(n_993), .B(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1005), .Y(n_1003) );
INVxp67_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1014), .Y(n_1012) );
INVxp67_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_1035), .B(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVxp67_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
XOR2x2_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1070), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1058), .Y(n_1080) );
NOR2x1_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1065), .Y(n_1058) );
NAND4xp25_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .C(n_1062), .D(n_1063), .Y(n_1059) );
NAND4xp25_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .C(n_1068), .D(n_1069), .Y(n_1065) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
endmodule