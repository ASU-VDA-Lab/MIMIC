module fake_jpeg_17388_n_184 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_12),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_8),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_36),
.B(n_49),
.Y(n_77)
);

CKINVDCx9p33_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_47),
.B(n_52),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_17),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_17),
.B(n_6),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_55),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_22),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_22),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_19),
.A2(n_7),
.B(n_13),
.C(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_16),
.B1(n_33),
.B2(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_74),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_78),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_23),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_43),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_110),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_46),
.B(n_54),
.C(n_40),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_105),
.B(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_44),
.B1(n_39),
.B2(n_23),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_113),
.B1(n_98),
.B2(n_94),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_40),
.B1(n_43),
.B2(n_48),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_106),
.B1(n_108),
.B2(n_116),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_28),
.B(n_30),
.C(n_43),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_114),
.C(n_96),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_30),
.B1(n_77),
.B2(n_61),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_76),
.B(n_65),
.C(n_79),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_58),
.B(n_87),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_59),
.B1(n_79),
.B2(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_64),
.Y(n_113)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_74),
.A3(n_73),
.B1(n_86),
.B2(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_72),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_64),
.B1(n_69),
.B2(n_72),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_120),
.B(n_125),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_58),
.C(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_123),
.C(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_108),
.C(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_130),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_100),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_94),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_92),
.B(n_112),
.C(n_91),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_121),
.C(n_123),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_102),
.B(n_109),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_103),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_152),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_153),
.B(n_120),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_155),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_98),
.B1(n_134),
.B2(n_127),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_135),
.B1(n_118),
.B2(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_126),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_136),
.B1(n_133),
.B2(n_128),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_140),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_118),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_132),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_124),
.C(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_162),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_164),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_155),
.B(n_145),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_171),
.A2(n_172),
.B1(n_156),
.B2(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_176),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_161),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.C(n_170),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_157),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_158),
.B(n_160),
.C(n_165),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_179),
.B(n_174),
.C(n_144),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_146),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_182),
.Y(n_184)
);


endmodule