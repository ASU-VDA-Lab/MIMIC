module real_jpeg_4375_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_58),
.B1(n_91),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_127),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_1),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_2),
.A2(n_140),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_8),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_5),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_6),
.Y(n_123)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_53),
.B1(n_57),
.B2(n_60),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_53),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_8),
.A2(n_53),
.B1(n_147),
.B2(n_150),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_153),
.B(n_154),
.C(n_158),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_104),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_8),
.B(n_22),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_8),
.B(n_219),
.C(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_89),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_8),
.B(n_84),
.C(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_199),
.B1(n_272),
.B2(n_273),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_13),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_197),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_169),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_129),
.C(n_159),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_16),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_97),
.B2(n_98),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_55),
.B2(n_96),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_20),
.B(n_55),
.C(n_97),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_47),
.B(n_48),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_21),
.A2(n_47),
.B1(n_48),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_21),
.A2(n_47),
.B1(n_48),
.B2(n_182),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_24),
.Y(n_135)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_24),
.Y(n_141)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_31),
.Y(n_149)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_39),
.Y(n_185)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_53),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_55),
.A2(n_96),
.B1(n_180),
.B2(n_181),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_55),
.B(n_180),
.C(n_240),
.Y(n_264)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B1(n_89),
.B2(n_90),
.Y(n_55)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_56),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_64),
.A2(n_65),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_80),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22x1_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_73),
.B2(n_76),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_82),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_124),
.B2(n_128),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_99),
.A2(n_103),
.B1(n_124),
.B2(n_128),
.Y(n_173)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_129),
.A2(n_130),
.B1(n_159),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_151),
.B2(n_152),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_131),
.A2(n_132),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_132),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_211),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_132),
.B(n_229),
.C(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_139),
.B1(n_145),
.B2(n_146),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_139),
.B1(n_146),
.B2(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_133),
.B(n_146),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_133),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_146),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_159),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_167),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_160),
.A2(n_161),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_160),
.A2(n_161),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_262)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_207),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_181),
.B1(n_215),
.B2(n_223),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_223),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_193),
.B(n_196),
.Y(n_188)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_266),
.B(n_271),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_254),
.B(n_265),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_235),
.B(n_253),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_225),
.B(n_234),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_213),
.B(n_224),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_210),
.B(n_212),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_233),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_239),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_238),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_257),
.C(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_252),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_251),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_251),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_264),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);


endmodule