module fake_jpeg_22326_n_225 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_28),
.B1(n_34),
.B2(n_26),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_46),
.B1(n_15),
.B2(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_15),
.B1(n_27),
.B2(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_52),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_26),
.B1(n_21),
.B2(n_19),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_30),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_75),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_29),
.B1(n_36),
.B2(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_16),
.B1(n_15),
.B2(n_21),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_49),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_74),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_16),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_44),
.C(n_43),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.C(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_40),
.B1(n_52),
.B2(n_51),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_76),
.B1(n_96),
.B2(n_91),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_85),
.B1(n_83),
.B2(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_114),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_51),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_65),
.C(n_53),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_83),
.C(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_63),
.B1(n_53),
.B2(n_97),
.Y(n_128)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_51),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_69),
.B(n_67),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_112),
.B(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_107),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_86),
.B(n_89),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_128),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_126),
.C(n_135),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_55),
.B(n_47),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_77),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_111),
.B(n_106),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_88),
.C(n_65),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_72),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_24),
.C(n_21),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_24),
.C(n_14),
.Y(n_155)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_153),
.B(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_146),
.B(n_149),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_156),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_117),
.B1(n_99),
.B2(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_99),
.B1(n_106),
.B2(n_109),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_135),
.B(n_137),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_160),
.C(n_163),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_155),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_133),
.C(n_136),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_167),
.B(n_22),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_134),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_134),
.C(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_127),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_22),
.B(n_18),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_1),
.C(n_2),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_47),
.C(n_14),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_156),
.C(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_176),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_181),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_142),
.B1(n_140),
.B2(n_6),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_18),
.B1(n_17),
.B2(n_7),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_22),
.C(n_18),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_163),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_164),
.CI(n_157),
.CON(n_182),
.SN(n_182)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_182),
.B(n_159),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_160),
.C(n_170),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_185),
.C(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_4),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_182),
.B1(n_173),
.B2(n_174),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_180),
.B1(n_17),
.B2(n_7),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_200),
.B(n_191),
.Y(n_205)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_184),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_4),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_206),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_210),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_17),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_209),
.Y(n_212)
);

AOI211xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_192),
.B(n_5),
.C(n_7),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_4),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_198),
.A3(n_201),
.B1(n_202),
.B2(n_200),
.C1(n_10),
.C2(n_11),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_213),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_8),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_9),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_218),
.B1(n_216),
.B2(n_9),
.Y(n_221)
);

AOI31xp67_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_208),
.A3(n_211),
.B(n_11),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_212),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_220),
.A2(n_221),
.B(n_9),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_10),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_10),
.Y(n_225)
);


endmodule