module real_aes_17555_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_917, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_917;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_0), .Y(n_585) );
AND2x4_ASAP7_75t_L g913 ( .A(n_1), .B(n_914), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_2), .A2(n_5), .B1(n_177), .B2(n_178), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_3), .A2(n_67), .B1(n_895), .B2(n_896), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_3), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_4), .A2(n_20), .B1(n_128), .B2(n_130), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_6), .A2(n_52), .B1(n_202), .B2(n_211), .Y(n_210) );
BUFx3_ASAP7_75t_L g620 ( .A(n_7), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_8), .A2(n_15), .B1(n_135), .B2(n_194), .Y(n_272) );
INVx1_ASAP7_75t_L g914 ( .A(n_9), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_10), .Y(n_255) );
XOR2xp5_ASAP7_75t_L g531 ( .A(n_11), .B(n_55), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_12), .B(n_175), .Y(n_562) );
OR2x2_ASAP7_75t_L g510 ( .A(n_13), .B(n_31), .Y(n_510) );
BUFx2_ASAP7_75t_L g908 ( .A(n_13), .Y(n_908) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_14), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_16), .B(n_217), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_17), .B(n_224), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_18), .A2(n_88), .B1(n_128), .B2(n_217), .Y(n_629) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_19), .A2(n_48), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_21), .B(n_130), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_22), .Y(n_149) );
INVx4_ASAP7_75t_R g232 ( .A(n_23), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_24), .B(n_133), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_25), .Y(n_898) );
AO32x1_ASAP7_75t_L g626 ( .A1(n_26), .A2(n_141), .A3(n_142), .B1(n_601), .B2(n_627), .Y(n_626) );
AO32x2_ASAP7_75t_L g661 ( .A1(n_26), .A2(n_141), .A3(n_142), .B1(n_601), .B2(n_627), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_27), .B(n_130), .Y(n_167) );
INVx1_ASAP7_75t_L g185 ( .A(n_28), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_SL g253 ( .A1(n_29), .A2(n_132), .B(n_135), .C(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_30), .A2(n_45), .B1(n_135), .B2(n_136), .Y(n_134) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_31), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_32), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_33), .A2(n_51), .B1(n_130), .B2(n_233), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_34), .B(n_564), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_35), .A2(n_93), .B1(n_128), .B2(n_136), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_36), .B(n_595), .Y(n_598) );
INVx1_ASAP7_75t_L g164 ( .A(n_37), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_38), .B(n_135), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_39), .A2(n_70), .B1(n_136), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_40), .A2(n_105), .B1(n_905), .B2(n_915), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_41), .Y(n_195) );
INVx2_ASAP7_75t_L g522 ( .A(n_42), .Y(n_522) );
INVx1_ASAP7_75t_L g508 ( .A(n_43), .Y(n_508) );
BUFx3_ASAP7_75t_L g529 ( .A(n_43), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_44), .B(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_46), .A2(n_87), .B1(n_135), .B2(n_136), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_47), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_49), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_50), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_53), .A2(n_81), .B1(n_160), .B2(n_595), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_54), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_56), .A2(n_85), .B1(n_128), .B2(n_217), .Y(n_616) );
INVx1_ASAP7_75t_L g144 ( .A(n_57), .Y(n_144) );
AND2x4_ASAP7_75t_L g146 ( .A(n_58), .B(n_147), .Y(n_146) );
AO22x1_ASAP7_75t_SL g114 ( .A1(n_59), .A2(n_69), .B1(n_115), .B2(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_59), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_60), .A2(n_92), .B1(n_136), .B2(n_174), .Y(n_173) );
AO22x1_ASAP7_75t_L g215 ( .A1(n_61), .A2(n_76), .B1(n_159), .B2(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_62), .B(n_128), .Y(n_561) );
INVx1_ASAP7_75t_L g147 ( .A(n_63), .Y(n_147) );
AND2x2_ASAP7_75t_L g256 ( .A(n_64), .B(n_141), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_65), .B(n_141), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_66), .A2(n_138), .B(n_202), .C(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g896 ( .A(n_67), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_68), .B(n_128), .C(n_566), .Y(n_567) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_71), .B(n_202), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_72), .Y(n_249) );
OAI22x1_ASAP7_75t_SL g108 ( .A1(n_73), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
AND2x2_ASAP7_75t_L g586 ( .A(n_74), .B(n_238), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_75), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_77), .B(n_130), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_78), .A2(n_99), .B1(n_160), .B2(n_217), .Y(n_609) );
INVx2_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_80), .B(n_197), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_82), .B(n_141), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_83), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_84), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_86), .B(n_151), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_89), .B(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_90), .A2(n_103), .B1(n_136), .B2(n_233), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_91), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_94), .B(n_141), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_95), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g537 ( .A(n_95), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_96), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_97), .B(n_224), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_98), .A2(n_181), .B(n_202), .C(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g237 ( .A(n_100), .B(n_238), .Y(n_237) );
NAND2xp33_ASAP7_75t_L g200 ( .A(n_101), .B(n_175), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_102), .Y(n_550) );
AO221x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_518), .B1(n_523), .B2(n_530), .C(n_897), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_112), .B(n_511), .Y(n_107) );
OAI31xp33_ASAP7_75t_L g511 ( .A1(n_108), .A2(n_113), .A3(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g111 ( .A(n_109), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_502), .Y(n_112) );
XNOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
OAI22x1_ASAP7_75t_L g533 ( .A1(n_117), .A2(n_534), .B1(n_538), .B2(n_890), .Y(n_533) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_392), .Y(n_117) );
NOR4xp25_ASAP7_75t_L g118 ( .A(n_119), .B(n_292), .C(n_334), .D(n_366), .Y(n_118) );
OAI211xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_186), .B(n_239), .C(n_277), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_152), .Y(n_122) );
INVx2_ASAP7_75t_L g305 ( .A(n_123), .Y(n_305) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g384 ( .A(n_124), .B(n_154), .Y(n_384) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_125), .B(n_170), .Y(n_242) );
AND2x2_ASAP7_75t_L g265 ( .A(n_125), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g291 ( .A(n_125), .Y(n_291) );
OR2x2_ASAP7_75t_L g354 ( .A(n_125), .B(n_170), .Y(n_354) );
AO31x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_140), .A3(n_145), .B(n_148), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_131), .B1(n_134), .B2(n_137), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_128), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_SL g595 ( .A(n_128), .Y(n_595) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_129), .Y(n_130) );
INVx3_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
INVx1_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx1_ASAP7_75t_L g202 ( .A(n_129), .Y(n_202) );
INVx1_ASAP7_75t_L g212 ( .A(n_129), .Y(n_212) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_129), .Y(n_217) );
INVx1_ASAP7_75t_L g233 ( .A(n_129), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_130), .B(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_130), .A2(n_233), .B1(n_580), .B2(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g642 ( .A(n_130), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_131), .A2(n_173), .B1(n_176), .B2(n_180), .Y(n_172) );
OAI22x1_ASAP7_75t_L g271 ( .A1(n_131), .A2(n_180), .B1(n_272), .B2(n_273), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_131), .A2(n_598), .B(n_599), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_131), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_131), .A2(n_132), .B1(n_616), .B2(n_617), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_131), .A2(n_137), .B1(n_641), .B2(n_643), .Y(n_640) );
INVx6_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_132), .A2(n_200), .B(n_201), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_132), .B(n_215), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_132), .A2(n_209), .B(n_215), .C(n_219), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_132), .A2(n_561), .B(n_562), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_132), .A2(n_252), .B1(n_628), .B2(n_629), .Y(n_627) );
BUFx8_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx1_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
INVx4_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_136), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
INVx2_ASAP7_75t_L g564 ( .A(n_136), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_137), .A2(n_166), .B(n_167), .Y(n_165) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_137), .A2(n_210), .B(n_213), .Y(n_209) );
AOI21x1_ASAP7_75t_L g593 ( .A1(n_137), .A2(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
AOI31xp67_ASAP7_75t_L g614 ( .A1(n_140), .A2(n_145), .A3(n_615), .B(n_618), .Y(n_614) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2x1_ASAP7_75t_L g203 ( .A(n_141), .B(n_204), .Y(n_203) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g168 ( .A(n_142), .B(n_145), .Y(n_168) );
INVx2_ASAP7_75t_L g547 ( .A(n_142), .Y(n_547) );
INVx2_ASAP7_75t_SL g591 ( .A(n_142), .Y(n_591) );
BUFx3_ASAP7_75t_L g605 ( .A(n_142), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_142), .B(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_142), .B(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
OAI21x1_ASAP7_75t_L g548 ( .A1(n_145), .A2(n_549), .B(n_552), .Y(n_548) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_145), .A2(n_560), .B(n_563), .Y(n_559) );
BUFx10_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g183 ( .A(n_146), .Y(n_183) );
INVx1_ASAP7_75t_L g220 ( .A(n_146), .Y(n_220) );
BUFx10_ASAP7_75t_L g236 ( .A(n_146), .Y(n_236) );
AO31x2_ASAP7_75t_L g639 ( .A1(n_146), .A2(n_605), .A3(n_640), .B(n_644), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx2_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_150), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g238 ( .A(n_150), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_150), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_150), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI21xp33_ASAP7_75t_L g219 ( .A1(n_151), .A2(n_213), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
INVx2_ASAP7_75t_L g274 ( .A(n_151), .Y(n_274) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g288 ( .A(n_153), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g300 ( .A(n_153), .Y(n_300) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_153), .Y(n_478) );
OR2x2_ASAP7_75t_L g491 ( .A(n_153), .B(n_492), .Y(n_491) );
OR2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_169), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_154), .B(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g263 ( .A(n_154), .Y(n_263) );
AND2x2_ASAP7_75t_L g311 ( .A(n_154), .B(n_312), .Y(n_311) );
NAND2x1p5_ASAP7_75t_SL g330 ( .A(n_154), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_154), .B(n_264), .Y(n_380) );
INVx1_ASAP7_75t_L g469 ( .A(n_154), .Y(n_469) );
AND2x2_ASAP7_75t_L g498 ( .A(n_154), .B(n_170), .Y(n_498) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_165), .B(n_168), .Y(n_156) );
OAI21xp33_ASAP7_75t_SL g157 ( .A1(n_158), .A2(n_159), .B(n_161), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_160), .B(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx4f_ASAP7_75t_L g252 ( .A(n_163), .Y(n_252) );
INVx1_ASAP7_75t_L g566 ( .A(n_163), .Y(n_566) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g264 ( .A(n_170), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_170), .B(n_291), .Y(n_313) );
INVx1_ASAP7_75t_L g333 ( .A(n_170), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_170), .B(n_266), .Y(n_385) );
AO31x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .A3(n_182), .B(n_184), .Y(n_170) );
AOI21x1_ASAP7_75t_L g245 ( .A1(n_171), .A2(n_246), .B(n_256), .Y(n_245) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_175), .A2(n_232), .B1(n_233), .B2(n_234), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g549 ( .A1(n_178), .A2(n_252), .B(n_550), .C(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_179), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_180), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g582 ( .A(n_181), .Y(n_582) );
INVx1_ASAP7_75t_SL g608 ( .A(n_181), .Y(n_608) );
AO31x2_ASAP7_75t_L g604 ( .A1(n_182), .A2(n_605), .A3(n_606), .B(n_610), .Y(n_604) );
INVx2_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_SL g601 ( .A(n_183), .Y(n_601) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_205), .Y(n_187) );
OR2x2_ASAP7_75t_L g282 ( .A(n_188), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g389 ( .A(n_188), .B(n_338), .Y(n_389) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g298 ( .A(n_189), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_189), .B(n_318), .Y(n_317) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_189), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
BUFx3_ASAP7_75t_L g309 ( .A(n_190), .Y(n_309) );
AND2x2_ASAP7_75t_L g345 ( .A(n_190), .B(n_326), .Y(n_345) );
AND2x2_ASAP7_75t_L g425 ( .A(n_190), .B(n_270), .Y(n_425) );
AND2x2_ASAP7_75t_L g438 ( .A(n_190), .B(n_222), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_199), .B(n_203), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .C(n_197), .Y(n_193) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_198), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_552) );
INVx2_ASAP7_75t_L g378 ( .A(n_205), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_205), .B(n_308), .Y(n_386) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_221), .Y(n_205) );
AND2x2_ASAP7_75t_L g297 ( .A(n_206), .B(n_222), .Y(n_297) );
INVx1_ASAP7_75t_L g405 ( .A(n_206), .Y(n_405) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g258 ( .A(n_207), .B(n_222), .Y(n_258) );
AND2x2_ASAP7_75t_L g322 ( .A(n_207), .B(n_221), .Y(n_322) );
AOI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_214), .B(n_218), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_212), .B(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g600 ( .A(n_217), .Y(n_600) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_220), .A2(n_247), .B(n_253), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_220), .A2(n_578), .B(n_583), .Y(n_577) );
AND2x2_ASAP7_75t_L g280 ( .A(n_221), .B(n_270), .Y(n_280) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g269 ( .A(n_222), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g338 ( .A(n_222), .B(n_270), .Y(n_338) );
INVx1_ASAP7_75t_L g349 ( .A(n_222), .Y(n_349) );
AND2x2_ASAP7_75t_L g412 ( .A(n_222), .B(n_260), .Y(n_412) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_226), .B(n_237), .Y(n_222) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_223), .A2(n_577), .B(n_586), .Y(n_576) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_235), .Y(n_226) );
INVx1_ASAP7_75t_L g554 ( .A(n_233), .Y(n_554) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_236), .A2(n_271), .A3(n_274), .B(n_275), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_257), .B1(n_261), .B2(n_267), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_240), .A2(n_311), .B1(n_314), .B2(n_316), .Y(n_310) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
OR2x2_ASAP7_75t_L g390 ( .A(n_242), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g496 ( .A(n_242), .Y(n_496) );
INVx1_ASAP7_75t_L g355 ( .A(n_243), .Y(n_355) );
OR2x2_ASAP7_75t_L g418 ( .A(n_243), .B(n_313), .Y(n_418) );
OR2x2_ASAP7_75t_L g289 ( .A(n_244), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_244), .B(n_263), .Y(n_365) );
AND2x2_ASAP7_75t_L g382 ( .A(n_244), .B(n_309), .Y(n_382) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_244), .Y(n_399) );
INVxp67_ASAP7_75t_L g447 ( .A(n_244), .Y(n_447) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g266 ( .A(n_245), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B(n_252), .Y(n_247) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_258), .Y(n_357) );
INVx3_ASAP7_75t_L g362 ( .A(n_258), .Y(n_362) );
AND2x2_ASAP7_75t_L g375 ( .A(n_258), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g475 ( .A(n_258), .B(n_437), .Y(n_475) );
INVx1_ASAP7_75t_L g268 ( .A(n_259), .Y(n_268) );
OR2x2_ASAP7_75t_L g452 ( .A(n_259), .B(n_427), .Y(n_452) );
BUFx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g376 ( .A(n_260), .B(n_286), .Y(n_376) );
AND2x2_ASAP7_75t_L g397 ( .A(n_260), .B(n_322), .Y(n_397) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_262), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g398 ( .A(n_262), .Y(n_398) );
AND2x2_ASAP7_75t_L g440 ( .A(n_262), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g341 ( .A(n_263), .Y(n_341) );
AND2x2_ASAP7_75t_L g372 ( .A(n_263), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_263), .B(n_331), .Y(n_391) );
AND2x2_ASAP7_75t_L g340 ( .A(n_265), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g456 ( .A(n_265), .Y(n_456) );
AND2x2_ASAP7_75t_L g479 ( .A(n_265), .B(n_469), .Y(n_479) );
INVx1_ASAP7_75t_L g492 ( .A(n_265), .Y(n_492) );
INVx2_ASAP7_75t_L g331 ( .A(n_266), .Y(n_331) );
OR2x2_ASAP7_75t_L g427 ( .A(n_266), .B(n_291), .Y(n_427) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_269), .B(n_308), .Y(n_315) );
INVx2_ASAP7_75t_L g286 ( .A(n_270), .Y(n_286) );
INVx2_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_270), .B(n_284), .Y(n_348) );
INVx2_ASAP7_75t_L g558 ( .A(n_274), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_287), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_280), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g421 ( .A(n_283), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx2_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g301 ( .A(n_289), .Y(n_301) );
INVxp67_ASAP7_75t_L g472 ( .A(n_289), .Y(n_472) );
OR2x2_ASAP7_75t_L g374 ( .A(n_290), .B(n_331), .Y(n_374) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND4xp25_ASAP7_75t_L g292 ( .A(n_293), .B(n_302), .C(n_310), .D(n_319), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .C(n_301), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_295), .A2(n_489), .B(n_491), .C(n_493), .Y(n_488) );
OR2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_297), .B(n_345), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_297), .B(n_401), .C(n_403), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_297), .B(n_376), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_297), .A2(n_402), .B1(n_494), .B2(n_497), .C(n_499), .Y(n_493) );
INVx1_ASAP7_75t_L g484 ( .A(n_298), .Y(n_484) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_303), .A2(n_311), .B1(n_346), .B2(n_420), .C(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_305), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g370 ( .A(n_306), .Y(n_370) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_308), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g485 ( .A(n_308), .B(n_336), .Y(n_485) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g321 ( .A(n_309), .Y(n_321) );
AND3x1_ASAP7_75t_L g494 ( .A(n_309), .B(n_495), .C(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g364 ( .A(n_313), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g434 ( .A(n_316), .Y(n_434) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g410 ( .A(n_318), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g437 ( .A(n_318), .Y(n_437) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B(n_328), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2x1_ASAP7_75t_L g335 ( .A(n_321), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g358 ( .A(n_326), .Y(n_358) );
OR2x2_ASAP7_75t_L g337 ( .A(n_327), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g450 ( .A(n_327), .Y(n_450) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_329), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
OR2x2_ASAP7_75t_L g406 ( .A(n_330), .B(n_354), .Y(n_406) );
INVx2_ASAP7_75t_L g495 ( .A(n_330), .Y(n_495) );
INVx1_ASAP7_75t_L g369 ( .A(n_331), .Y(n_369) );
NOR4xp25_ASAP7_75t_L g499 ( .A(n_331), .B(n_362), .C(n_500), .D(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_332), .Y(n_501) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g487 ( .A(n_333), .Y(n_487) );
OAI211xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_339), .B(n_342), .C(n_350), .Y(n_334) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g474 ( .A(n_337), .Y(n_474) );
INVx2_ASAP7_75t_L g459 ( .A(n_338), .Y(n_459) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_340), .A2(n_343), .B(n_346), .Y(n_342) );
OR2x2_ASAP7_75t_L g426 ( .A(n_341), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g444 ( .A(n_341), .B(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g360 ( .A(n_345), .Y(n_360) );
AND2x4_ASAP7_75t_SL g449 ( .A(n_345), .B(n_450), .Y(n_449) );
INVx3_ASAP7_75t_R g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_348), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
AOI32xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_356), .A3(n_358), .B1(n_359), .B2(n_363), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_353), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_353), .Y(n_414) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g431 ( .A(n_354), .B(n_369), .Y(n_431) );
INVx2_ASAP7_75t_L g445 ( .A(n_354), .Y(n_445) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_362), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B(n_371), .C(n_387), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B(n_377), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_376), .B(n_463), .Y(n_462) );
OAI32xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .A3(n_381), .B1(n_383), .B2(n_386), .Y(n_377) );
INVx1_ASAP7_75t_L g463 ( .A(n_378), .Y(n_463) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g455 ( .A(n_380), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_464), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_394), .B(n_419), .C(n_432), .D(n_460), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_395), .B(n_407), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_406), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g446 ( .A(n_398), .B(n_447), .Y(n_446) );
OAI32xp33_ASAP7_75t_L g451 ( .A1(n_398), .A2(n_452), .A3(n_453), .B1(n_455), .B2(n_457), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_399), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_401), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g458 ( .A(n_404), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g490 ( .A(n_404), .Y(n_490) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g454 ( .A(n_405), .Y(n_454) );
OAI22x1_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_413), .B1(n_415), .B2(n_416), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_417), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_421), .B(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_428), .B2(n_429), .Y(n_423) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_425), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g500 ( .A(n_425), .Y(n_500) );
INVx2_ASAP7_75t_L g441 ( .A(n_427), .Y(n_441) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR3xp33_ASAP7_75t_SL g432 ( .A(n_433), .B(n_442), .C(n_451), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_439), .Y(n_433) );
NAND2xp33_ASAP7_75t_L g461 ( .A(n_435), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g497 ( .A(n_441), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g468 ( .A(n_445), .B(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_447), .Y(n_467) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_470), .C(n_482), .Y(n_464) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g473 ( .A(n_469), .Y(n_473) );
AOI222xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_474), .B1(n_475), .B2(n_476), .C1(n_479), .C2(n_480), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
O2A1O1Ixp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_486), .C(n_488), .Y(n_482) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx12f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx5_ASAP7_75t_L g514 ( .A(n_505), .Y(n_514) );
AND2x6_ASAP7_75t_SL g505 ( .A(n_506), .B(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_509), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2x1_ASAP7_75t_L g904 ( .A(n_510), .B(n_529), .Y(n_904) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_514), .B(n_517), .Y(n_516) );
OAI21xp33_ASAP7_75t_L g897 ( .A1(n_515), .A2(n_898), .B(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx8_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g526 ( .A(n_522), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_522), .B(n_902), .Y(n_901) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx6_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x6_ASAP7_75t_SL g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NOR3x1_ASAP7_75t_L g911 ( .A(n_529), .B(n_536), .C(n_912), .Y(n_911) );
XOR2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
XNOR2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_893), .Y(n_532) );
INVx4_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g892 ( .A(n_537), .Y(n_892) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_764), .Y(n_539) );
AND5x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_690), .C(n_710), .D(n_726), .E(n_746), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_650), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_569), .B(n_621), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g758 ( .A(n_544), .Y(n_758) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g744 ( .A(n_545), .Y(n_744) );
OR2x2_ASAP7_75t_L g781 ( .A(n_545), .B(n_782), .Y(n_781) );
OR2x2_ASAP7_75t_L g847 ( .A(n_545), .B(n_603), .Y(n_847) );
OR2x2_ASAP7_75t_L g856 ( .A(n_545), .B(n_675), .Y(n_856) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_557), .Y(n_545) );
BUFx2_ASAP7_75t_L g633 ( .A(n_546), .Y(n_633) );
INVx1_ASAP7_75t_L g649 ( .A(n_546), .Y(n_649) );
INVx2_ASAP7_75t_SL g708 ( .A(n_546), .Y(n_708) );
AND2x2_ASAP7_75t_L g729 ( .A(n_546), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g833 ( .A(n_546), .B(n_604), .Y(n_833) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_556), .Y(n_546) );
OA21x2_ASAP7_75t_L g673 ( .A1(n_547), .A2(n_548), .B(n_556), .Y(n_673) );
AND2x2_ASAP7_75t_L g689 ( .A(n_557), .B(n_673), .Y(n_689) );
AND2x2_ASAP7_75t_L g799 ( .A(n_557), .B(n_657), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_568), .Y(n_557) );
OAI21x1_ASAP7_75t_L g636 ( .A1(n_558), .A2(n_559), .B(n_568), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_587), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_573), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g733 ( .A(n_574), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_575), .Y(n_631) );
AND2x2_ASAP7_75t_L g663 ( .A(n_575), .B(n_639), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_575), .Y(n_667) );
INVx1_ASAP7_75t_L g705 ( .A(n_575), .Y(n_705) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g646 ( .A(n_576), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_582), .Y(n_578) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_603), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g732 ( .A(n_588), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g630 ( .A(n_589), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g659 ( .A(n_589), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g668 ( .A(n_589), .Y(n_668) );
INVx3_ASAP7_75t_L g680 ( .A(n_589), .Y(n_680) );
BUFx2_ASAP7_75t_L g718 ( .A(n_589), .Y(n_718) );
INVxp67_ASAP7_75t_L g738 ( .A(n_589), .Y(n_738) );
AND2x2_ASAP7_75t_L g761 ( .A(n_589), .B(n_661), .Y(n_761) );
INVx1_ASAP7_75t_L g775 ( .A(n_589), .Y(n_775) );
OR2x2_ASAP7_75t_L g796 ( .A(n_589), .B(n_660), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_589), .B(n_639), .Y(n_852) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B(n_602), .Y(n_590) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_597), .B(n_601), .Y(n_592) );
INVx1_ASAP7_75t_L g763 ( .A(n_603), .Y(n_763) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_612), .Y(n_603) );
AND2x2_ASAP7_75t_L g648 ( .A(n_604), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g675 ( .A(n_604), .Y(n_675) );
INVx2_ASAP7_75t_L g694 ( .A(n_604), .Y(n_694) );
AND2x2_ASAP7_75t_L g709 ( .A(n_604), .B(n_657), .Y(n_709) );
INVx1_ASAP7_75t_L g730 ( .A(n_604), .Y(n_730) );
AND2x2_ASAP7_75t_L g788 ( .A(n_604), .B(n_612), .Y(n_788) );
AND2x2_ASAP7_75t_L g798 ( .A(n_604), .B(n_673), .Y(n_798) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g635 ( .A(n_613), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g657 ( .A(n_614), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_632), .B1(n_637), .B2(n_647), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_622), .A2(n_850), .B1(n_854), .B2(n_855), .Y(n_849) );
AND2x4_ASAP7_75t_L g622 ( .A(n_623), .B(n_630), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_623), .B(n_663), .Y(n_754) );
NAND2xp5_ASAP7_75t_R g773 ( .A(n_623), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g785 ( .A(n_625), .B(n_680), .Y(n_785) );
INVx1_ASAP7_75t_L g853 ( .A(n_625), .Y(n_853) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g681 ( .A(n_626), .B(n_639), .Y(n_681) );
OR2x2_ASAP7_75t_L g722 ( .A(n_626), .B(n_639), .Y(n_722) );
INVx1_ASAP7_75t_L g734 ( .A(n_626), .Y(n_734) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_630), .Y(n_876) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
AND2x2_ASAP7_75t_L g691 ( .A(n_633), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_633), .B(n_709), .Y(n_725) );
INVx1_ASAP7_75t_L g787 ( .A(n_633), .Y(n_787) );
AND2x2_ASAP7_75t_L g647 ( .A(n_634), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_634), .B(n_729), .Y(n_878) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g695 ( .A(n_635), .Y(n_695) );
INVx1_ASAP7_75t_L g771 ( .A(n_635), .Y(n_771) );
OR2x2_ASAP7_75t_L g824 ( .A(n_635), .B(n_693), .Y(n_824) );
INVx2_ASAP7_75t_L g655 ( .A(n_636), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_637), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_637), .B(n_738), .Y(n_759) );
INVx1_ASAP7_75t_L g819 ( .A(n_637), .Y(n_819) );
OAI31xp33_ASAP7_75t_L g875 ( .A1(n_637), .A2(n_791), .A3(n_876), .B(n_877), .Y(n_875) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_646), .Y(n_637) );
AND2x4_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g741 ( .A(n_638), .B(n_661), .Y(n_741) );
INVx1_ASAP7_75t_L g776 ( .A(n_638), .Y(n_776) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g704 ( .A(n_639), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g684 ( .A(n_646), .Y(n_684) );
INVx1_ASAP7_75t_L g740 ( .A(n_646), .Y(n_740) );
OR2x2_ASAP7_75t_L g814 ( .A(n_646), .B(n_734), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_646), .B(n_680), .Y(n_872) );
AND2x4_ASAP7_75t_L g652 ( .A(n_648), .B(n_653), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_658), .B1(n_664), .B2(n_669), .C(n_678), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g751 ( .A(n_654), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g793 ( .A(n_654), .B(n_694), .Y(n_793) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g677 ( .A(n_655), .Y(n_677) );
INVx1_ASAP7_75t_L g687 ( .A(n_656), .Y(n_687) );
INVx1_ASAP7_75t_L g745 ( .A(n_656), .Y(n_745) );
AND2x2_ASAP7_75t_L g809 ( .A(n_656), .B(n_730), .Y(n_809) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g672 ( .A(n_657), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
AND2x2_ASAP7_75t_L g714 ( .A(n_659), .B(n_704), .Y(n_714) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g701 ( .A(n_661), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_662), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
BUFx2_ASAP7_75t_L g697 ( .A(n_663), .Y(n_697) );
AND2x4_ASAP7_75t_L g784 ( .A(n_663), .B(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g863 ( .A(n_663), .B(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_665), .B(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx2_ASAP7_75t_L g804 ( .A(n_666), .Y(n_804) );
INVx1_ASAP7_75t_L g720 ( .A(n_667), .Y(n_720) );
AND2x2_ASAP7_75t_L g703 ( .A(n_668), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g778 ( .A(n_668), .B(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_SL g813 ( .A(n_668), .Y(n_813) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_668), .Y(n_864) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_672), .B(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_672), .B(n_728), .Y(n_859) );
INVx1_ASAP7_75t_L g752 ( .A(n_673), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g728 ( .A(n_677), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B(n_685), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g829 ( .A(n_680), .B(n_741), .Y(n_829) );
AND2x2_ASAP7_75t_L g682 ( .A(n_681), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_SL g779 ( .A(n_681), .Y(n_779) );
INVx1_ASAP7_75t_L g712 ( .A(n_682), .Y(n_712) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
AND2x2_ASAP7_75t_L g749 ( .A(n_687), .B(n_750), .Y(n_749) );
OR2x2_ASAP7_75t_L g806 ( .A(n_687), .B(n_751), .Y(n_806) );
OR2x2_ASAP7_75t_L g888 ( .A(n_688), .B(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_696), .A3(n_698), .B1(n_702), .B2(n_706), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_692), .A2(n_797), .B1(n_829), .B2(n_863), .Y(n_862) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx2_ASAP7_75t_L g757 ( .A(n_693), .Y(n_757) );
NAND4xp25_ASAP7_75t_L g767 ( .A(n_693), .B(n_697), .C(n_768), .D(n_769), .Y(n_767) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g822 ( .A(n_694), .B(n_775), .Y(n_822) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g702 ( .A(n_699), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g882 ( .A(n_701), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g836 ( .A1(n_703), .A2(n_809), .B(n_837), .C(n_838), .Y(n_836) );
BUFx2_ASAP7_75t_L g791 ( .A(n_704), .Y(n_791) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_708), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g845 ( .A(n_708), .Y(n_845) );
INVx2_ASAP7_75t_L g782 ( .A(n_709), .Y(n_782) );
AND2x4_ASAP7_75t_L g838 ( .A(n_709), .B(n_750), .Y(n_838) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_715), .B(n_723), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
AOI322xp5_ASAP7_75t_L g816 ( .A1(n_717), .A2(n_817), .A3(n_819), .B1(n_820), .B2(n_821), .C1(n_823), .C2(n_825), .Y(n_816) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g835 ( .A(n_718), .B(n_722), .Y(n_835) );
INVx1_ASAP7_75t_L g846 ( .A(n_719), .Y(n_846) );
AND2x4_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
AND2x2_ASAP7_75t_L g840 ( .A(n_720), .B(n_761), .Y(n_840) );
AND2x2_ASAP7_75t_L g861 ( .A(n_721), .B(n_740), .Y(n_861) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g871 ( .A(n_722), .B(n_872), .Y(n_871) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI222xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_731), .B1(n_735), .B2(n_739), .C1(n_742), .C2(n_917), .Y(n_726) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_727), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx2_ASAP7_75t_L g769 ( .A(n_728), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_729), .B(n_799), .Y(n_818) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g803 ( .A(n_738), .B(n_804), .Y(n_803) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_738), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_739), .Y(n_868) );
AND2x4_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx3_ASAP7_75t_L g815 ( .A(n_741), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_742), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_753), .B(n_755), .Y(n_746) );
INVxp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_750), .B(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g837 ( .A(n_750), .Y(n_837) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI32xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .A3(n_759), .B1(n_760), .B2(n_762), .Y(n_755) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g858 ( .A(n_757), .B(n_859), .Y(n_858) );
BUFx2_ASAP7_75t_L g768 ( .A(n_761), .Y(n_768) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_841), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_800), .C(n_827), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .C(n_783), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_769), .B(n_787), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_777), .B2(n_780), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_786), .B(n_789), .Y(n_783) );
INVx1_ASAP7_75t_L g826 ( .A(n_785), .Y(n_826) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g889 ( .A(n_788), .Y(n_889) );
OAI21xp33_ASAP7_75t_SL g789 ( .A1(n_790), .A2(n_792), .B(n_794), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_L g873 ( .A(n_793), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
INVx2_ASAP7_75t_L g848 ( .A(n_795), .Y(n_848) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
AND2x2_ASAP7_75t_L g831 ( .A(n_799), .B(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_816), .Y(n_800) );
AOI22xp5_ASAP7_75t_SL g801 ( .A1(n_802), .A2(n_805), .B1(n_807), .B2(n_810), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_804), .B(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVxp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g844 ( .A(n_809), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_815), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2x1p5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NAND4xp25_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .C(n_836), .D(n_839), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_834), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_838), .B(n_840), .Y(n_839) );
NOR4xp25_ASAP7_75t_L g841 ( .A(n_842), .B(n_857), .C(n_865), .D(n_874), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_846), .B1(n_847), .B2(n_848), .C(n_849), .Y(n_842) );
INVx2_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g854 ( .A(n_847), .Y(n_854) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g883 ( .A(n_851), .Y(n_883) );
OR2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g886 ( .A(n_853), .Y(n_886) );
INVx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI21xp5_ASAP7_75t_SL g857 ( .A1(n_858), .A2(n_860), .B(n_862), .Y(n_857) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
O2A1O1Ixp33_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_868), .B(n_869), .C(n_873), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_879), .Y(n_874) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
OAI31xp33_ASAP7_75t_SL g879 ( .A1(n_880), .A2(n_883), .A3(n_884), .B(n_887), .Y(n_879) );
INVxp67_ASAP7_75t_SL g880 ( .A(n_881), .Y(n_880) );
INVxp67_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g903 ( .A(n_892), .B(n_904), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
BUFx10_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx6f_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
INVx6_ASAP7_75t_L g915 ( .A(n_906), .Y(n_915) );
AND2x6_ASAP7_75t_L g906 ( .A(n_907), .B(n_911), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
INVxp33_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_SL g912 ( .A(n_913), .Y(n_912) );
endmodule