module fake_jpeg_22183_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_18),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_28),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_30),
.B1(n_24),
.B2(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_37),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_22),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_37),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_22),
.B(n_21),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_78),
.B(n_55),
.Y(n_93)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_68),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_41),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_77),
.B1(n_85),
.B2(n_41),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_79),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_41),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_37),
.B1(n_35),
.B2(n_22),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_21),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_84),
.C(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_47),
.B1(n_24),
.B2(n_18),
.Y(n_86)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_93),
.B1(n_107),
.B2(n_77),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_96),
.C(n_59),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_112),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_52),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_47),
.B1(n_55),
.B2(n_52),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_75),
.B1(n_85),
.B2(n_60),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_52),
.B1(n_44),
.B2(n_49),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_24),
.B(n_29),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_29),
.B(n_25),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_52),
.B1(n_44),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_44),
.B1(n_35),
.B2(n_20),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_49),
.B1(n_46),
.B2(n_29),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_40),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_81),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_102),
.Y(n_169)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_72),
.B(n_66),
.C(n_80),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_103),
.B1(n_107),
.B2(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_122),
.C(n_136),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_59),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_138),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_40),
.C(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_0),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_98),
.B1(n_108),
.B2(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_28),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_100),
.B(n_94),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_0),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_40),
.C(n_74),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_73),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_20),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_96),
.Y(n_149)
);

CKINVDCx10_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_140),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_156),
.C(n_165),
.Y(n_188)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_150),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_157),
.B1(n_168),
.B2(n_32),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_130),
.Y(n_170)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_158),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_127),
.B(n_134),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_91),
.B1(n_86),
.B2(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_137),
.B1(n_128),
.B2(n_123),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_105),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_105),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_146),
.C(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_102),
.B1(n_62),
.B2(n_61),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_173),
.C(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_172),
.B(n_194),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_138),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_162),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_161),
.B1(n_159),
.B2(n_141),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_187),
.B(n_4),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_183),
.B1(n_168),
.B2(n_157),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_189),
.B(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_134),
.B1(n_89),
.B2(n_106),
.Y(n_183)
);

OAI322xp33_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_31),
.A3(n_17),
.B1(n_19),
.B2(n_26),
.C1(n_23),
.C2(n_104),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_160),
.C(n_10),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_106),
.B(n_32),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_20),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_31),
.B1(n_26),
.B2(n_19),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_8),
.B1(n_13),
.B2(n_3),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_20),
.B(n_28),
.C(n_2),
.D(n_3),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_167),
.C(n_169),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_25),
.B(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_201),
.B1(n_204),
.B2(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_150),
.B1(n_154),
.B2(n_143),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_140),
.B(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_188),
.C(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_195),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_166),
.B(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_145),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_190),
.C(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_220),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_201),
.B(n_212),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_182),
.C(n_181),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_174),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_225),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_180),
.CI(n_189),
.CON(n_225),
.SN(n_225)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_227),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

OAI322xp33_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_175),
.A3(n_192),
.B1(n_191),
.B2(n_179),
.C1(n_9),
.C2(n_11),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_230),
.CI(n_211),
.CON(n_232),
.SN(n_232)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_179),
.C(n_5),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_225),
.C(n_234),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_224),
.B1(n_198),
.B2(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_196),
.B1(n_202),
.B2(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_241),
.B1(n_244),
.B2(n_219),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_231),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_209),
.B1(n_203),
.B2(n_210),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_215),
.C(n_216),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_246),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_218),
.C(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_217),
.C(n_228),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_247),
.A2(n_250),
.B(n_239),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_253),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_230),
.C(n_210),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_225),
.B(n_200),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_239),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_4),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_6),
.C(n_12),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_237),
.B1(n_241),
.B2(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_262),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_247),
.B(n_254),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_252),
.B(n_9),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_6),
.B(n_9),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_257),
.C(n_15),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_13),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_269),
.B(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_273),
.B1(n_263),
.B2(n_266),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_270),
.B(n_255),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_273),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_276),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_13),
.Y(n_280)
);


endmodule