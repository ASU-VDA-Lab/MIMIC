module fake_netlist_1_759_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_8), .B(n_7), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_9), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_15), .B(n_0), .C(n_1), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_12), .B(n_0), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_13), .B1(n_14), .B2(n_17), .Y(n_24) );
AOI21xp5_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_16), .B(n_13), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_11), .B1(n_17), .B2(n_14), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_19), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_24), .B(n_23), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_18), .B1(n_17), .B2(n_14), .C(n_19), .Y(n_29) );
NAND4xp25_ASAP7_75t_SL g30 ( .A(n_25), .B(n_18), .C(n_22), .D(n_4), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_28), .B(n_2), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_17), .Y(n_32) );
NAND2xp5_ASAP7_75t_SL g33 ( .A(n_31), .B(n_17), .Y(n_33) );
INVx2_ASAP7_75t_SL g34 ( .A(n_32), .Y(n_34) );
NOR2xp33_ASAP7_75t_L g35 ( .A(n_31), .B(n_30), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AOI32xp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_2), .A3(n_3), .B1(n_5), .B2(n_6), .Y(n_37) );
BUFx3_ASAP7_75t_L g38 ( .A(n_33), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_36), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_38), .B1(n_17), .B2(n_37), .Y(n_40) );
AOI322xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_39), .A3(n_38), .B1(n_6), .B2(n_5), .C1(n_27), .C2(n_10), .Y(n_41) );
endmodule