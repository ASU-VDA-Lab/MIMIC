module fake_jpeg_3889_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_6),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_27),
.Y(n_50)
);

CKINVDCx9p33_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_31),
.B1(n_32),
.B2(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_33),
.B1(n_41),
.B2(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_53),
.B1(n_21),
.B2(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_16),
.B1(n_22),
.B2(n_18),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_33),
.B1(n_41),
.B2(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_63),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_34),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_24),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_33),
.B1(n_18),
.B2(n_22),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_74),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_36),
.C(n_35),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_28),
.B1(n_48),
.B2(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_60),
.C(n_68),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_100),
.B1(n_106),
.B2(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_53),
.B1(n_55),
.B2(n_46),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_26),
.B1(n_51),
.B2(n_83),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_55),
.B(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_36),
.B(n_35),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_110),
.B(n_102),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_88),
.B1(n_99),
.B2(n_94),
.C(n_84),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_38),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_58),
.B1(n_63),
.B2(n_59),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_114),
.B1(n_119),
.B2(n_123),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_64),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_122),
.C(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_26),
.B1(n_47),
.B2(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_47),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_37),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_37),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_126),
.B1(n_96),
.B2(n_117),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_47),
.B1(n_37),
.B2(n_77),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_94),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_132),
.B(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_145),
.C(n_42),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_84),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_108),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_146),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_96),
.B(n_85),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_23),
.B(n_42),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_107),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_38),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_124),
.B1(n_123),
.B2(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_147),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_114),
.B1(n_110),
.B2(n_120),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_159),
.B1(n_5),
.B2(n_7),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_155),
.B(n_156),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_145),
.C(n_6),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_51),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_5),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_163),
.B(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_107),
.B1(n_74),
.B2(n_42),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_164),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_14),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_1),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_171),
.C(n_172),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_143),
.B1(n_140),
.B2(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_144),
.B1(n_137),
.B2(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_10),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_10),
.C(n_12),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_11),
.C(n_13),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_151),
.Y(n_181)
);

OAI21x1_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_153),
.B(n_170),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_179),
.B(n_180),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_165),
.C(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_190),
.C(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_161),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_191),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_176),
.C(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_153),
.B1(n_164),
.B2(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_158),
.C(n_172),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_187),
.B1(n_180),
.B2(n_11),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_189),
.B(n_8),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_193),
.B(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_8),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_9),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_197),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_201),
.Y(n_204)
);


endmodule