module fake_jpeg_24119_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_26),
.B1(n_19),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_56),
.B1(n_30),
.B2(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_30),
.B1(n_20),
.B2(n_18),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_17),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_21),
.C(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_61),
.B1(n_51),
.B2(n_20),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_37),
.B(n_36),
.C(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_62),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_1),
.B(n_2),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_21),
.B(n_22),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_60),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_41),
.C(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_51),
.B1(n_43),
.B2(n_35),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_91),
.B1(n_68),
.B2(n_63),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_14),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_41),
.B1(n_58),
.B2(n_28),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_29),
.B(n_28),
.C(n_25),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_32),
.B1(n_69),
.B2(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_18),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_84),
.Y(n_95)
);

AOI221xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_99),
.B1(n_29),
.B2(n_28),
.C(n_40),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_1),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_106),
.B1(n_76),
.B2(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_41),
.B1(n_37),
.B2(n_40),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_3),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_86),
.B(n_91),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_114),
.B(n_120),
.C(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_75),
.B(n_81),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_118),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_89),
.C(n_80),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_108),
.C(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_45),
.Y(n_115)
);

OAI322xp33_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_110),
.A3(n_116),
.B1(n_117),
.B2(n_120),
.C1(n_99),
.C2(n_119),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_45),
.B(n_44),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_44),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_104),
.Y(n_130)
);

NOR4xp25_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_134),
.C(n_120),
.D(n_118),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_96),
.B1(n_121),
.B2(n_44),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.C(n_132),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_122),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_107),
.C(n_101),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_103),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_3),
.C(n_4),
.Y(n_143)
);

NOR4xp25_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_96),
.C(n_99),
.D(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_139),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_116),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_143),
.C(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_141),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_121),
.C(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_148),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_125),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_140),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_125),
.CI(n_5),
.CON(n_153),
.SN(n_153)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_156),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_152),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_8),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_146),
.B1(n_155),
.B2(n_154),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_159),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_148),
.C(n_8),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_6),
.B(n_8),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_10),
.C(n_11),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_166),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_167),
.B(n_164),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_10),
.Y(n_170)
);


endmodule