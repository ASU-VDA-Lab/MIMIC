module fake_jpeg_31593_n_93 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_55),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_35),
.B(n_32),
.C(n_37),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_1),
.C(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_39),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_32),
.B1(n_40),
.B2(n_14),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_49),
.B1(n_7),
.B2(n_11),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_6),
.Y(n_67)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_64),
.B(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_5),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

AO21x2_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_49),
.B(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_74),
.B1(n_9),
.B2(n_12),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_7),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_13),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_77),
.B1(n_70),
.B2(n_73),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_70),
.B1(n_68),
.B2(n_17),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_15),
.B(n_18),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_82),
.B1(n_80),
.B2(n_77),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_78),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_76),
.B1(n_20),
.B2(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_19),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_24),
.B(n_25),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_76),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_26),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_30),
.Y(n_93)
);


endmodule