module real_aes_2028_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_0), .B(n_122), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_1), .A2(n_131), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_2), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_3), .B(n_122), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_4), .B(n_138), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_5), .B(n_138), .Y(n_508) );
INVx1_ASAP7_75t_L g129 ( .A(n_6), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_7), .B(n_138), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g791 ( .A(n_8), .Y(n_791) );
NAND2xp33_ASAP7_75t_L g489 ( .A(n_9), .B(n_140), .Y(n_489) );
AND2x2_ASAP7_75t_L g158 ( .A(n_10), .B(n_147), .Y(n_158) );
AND2x2_ASAP7_75t_L g167 ( .A(n_11), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
AOI221x1_ASAP7_75t_L g530 ( .A1(n_13), .A2(n_24), .B1(n_122), .B2(n_131), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_14), .B(n_138), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_15), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g789 ( .A(n_15), .B(n_790), .C(n_792), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_16), .B(n_122), .Y(n_485) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_17), .A2(n_147), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_18), .B(n_142), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_19), .B(n_138), .Y(n_468) );
AO21x1_ASAP7_75t_L g503 ( .A1(n_20), .A2(n_122), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_21), .B(n_122), .Y(n_192) );
INVx1_ASAP7_75t_L g455 ( .A(n_22), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_23), .A2(n_92), .B1(n_122), .B2(n_231), .Y(n_230) );
NAND2x1_ASAP7_75t_L g517 ( .A(n_25), .B(n_138), .Y(n_517) );
NAND2x1_ASAP7_75t_L g478 ( .A(n_26), .B(n_140), .Y(n_478) );
OR2x2_ASAP7_75t_L g145 ( .A(n_27), .B(n_89), .Y(n_145) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_27), .A2(n_89), .B(n_144), .Y(n_148) );
OAI22x1_ASAP7_75t_R g779 ( .A1(n_28), .A2(n_780), .B1(n_781), .B2(n_784), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_28), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_29), .B(n_140), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_30), .B(n_138), .Y(n_488) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_31), .A2(n_168), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_32), .B(n_140), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_33), .A2(n_131), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_34), .B(n_138), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_35), .A2(n_131), .B(n_549), .Y(n_548) );
XNOR2x2_ASAP7_75t_SL g106 ( .A(n_36), .B(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g128 ( .A(n_37), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g132 ( .A(n_37), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g239 ( .A(n_37), .Y(n_239) );
OR2x6_ASAP7_75t_L g453 ( .A(n_38), .B(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g792 ( .A(n_38), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_39), .B(n_122), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_40), .B(n_122), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_41), .B(n_138), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_42), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_43), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_44), .B(n_140), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_45), .B(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_46), .A2(n_131), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_47), .A2(n_131), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_48), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_49), .B(n_140), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_50), .B(n_122), .Y(n_174) );
INVx1_ASAP7_75t_L g125 ( .A(n_51), .Y(n_125) );
INVx1_ASAP7_75t_L g135 ( .A(n_51), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_52), .A2(n_69), .B1(n_782), .B2(n_783), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_52), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_53), .B(n_138), .Y(n_165) );
AND2x2_ASAP7_75t_L g203 ( .A(n_54), .B(n_142), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_55), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_56), .B(n_140), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_57), .B(n_138), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_58), .B(n_140), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_59), .A2(n_131), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_60), .B(n_122), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_61), .B(n_122), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_62), .A2(n_131), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g198 ( .A(n_63), .B(n_143), .Y(n_198) );
AO21x1_ASAP7_75t_L g505 ( .A1(n_64), .A2(n_131), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_65), .B(n_122), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_66), .A2(n_83), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_67), .B(n_140), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_68), .B(n_122), .Y(n_480) );
INVx1_ASAP7_75t_L g783 ( .A(n_69), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_70), .B(n_140), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_71), .A2(n_97), .B1(n_131), .B2(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_72), .B(n_138), .Y(n_195) );
AND2x2_ASAP7_75t_L g553 ( .A(n_73), .B(n_143), .Y(n_553) );
INVx1_ASAP7_75t_L g127 ( .A(n_74), .Y(n_127) );
INVx1_ASAP7_75t_L g133 ( .A(n_74), .Y(n_133) );
AND2x2_ASAP7_75t_L g481 ( .A(n_75), .B(n_168), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_76), .B(n_140), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_77), .A2(n_131), .B(n_207), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_78), .A2(n_131), .B(n_136), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_79), .A2(n_131), .B(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g189 ( .A(n_80), .B(n_143), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_81), .B(n_142), .Y(n_228) );
INVx1_ASAP7_75t_L g456 ( .A(n_82), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_82), .B(n_455), .Y(n_788) );
INVx1_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_84), .B(n_122), .Y(n_470) );
AND2x2_ASAP7_75t_L g491 ( .A(n_85), .B(n_168), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_86), .A2(n_106), .B1(n_750), .B2(n_754), .Y(n_749) );
AND2x2_ASAP7_75t_L g146 ( .A(n_87), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g504 ( .A(n_88), .B(n_179), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_90), .B(n_140), .Y(n_469) );
AND2x2_ASAP7_75t_L g520 ( .A(n_91), .B(n_168), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_93), .B(n_138), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_94), .A2(n_131), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_95), .B(n_140), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_96), .A2(n_131), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_98), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_99), .B(n_138), .Y(n_496) );
BUFx2_ASAP7_75t_L g197 ( .A(n_100), .Y(n_197) );
BUFx2_ASAP7_75t_L g762 ( .A(n_101), .Y(n_762) );
BUFx2_ASAP7_75t_SL g771 ( .A(n_101), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_102), .A2(n_131), .B(n_487), .Y(n_486) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_785), .B(n_793), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_758), .B(n_769), .Y(n_104) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B(n_749), .Y(n_105) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_448), .B1(n_457), .B2(n_747), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_113), .A2(n_450), .B1(n_751), .B2(n_752), .Y(n_750) );
OAI22x1_ASAP7_75t_SL g776 ( .A1(n_113), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
INVx5_ASAP7_75t_L g777 ( .A(n_113), .Y(n_777) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_352), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_277), .C(n_313), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_251), .Y(n_115) );
AOI211xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_169), .B(n_199), .C(n_224), .Y(n_116) );
AND2x2_ASAP7_75t_L g342 ( .A(n_117), .B(n_201), .Y(n_342) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_149), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_118), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g375 ( .A(n_118), .B(n_257), .Y(n_375) );
AND2x2_ASAP7_75t_L g391 ( .A(n_118), .B(n_216), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_118), .B(n_401), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_118), .B(n_425), .Y(n_424) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_SL g211 ( .A(n_119), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g246 ( .A(n_119), .Y(n_246) );
AND2x2_ASAP7_75t_L g293 ( .A(n_119), .B(n_226), .Y(n_293) );
AND2x2_ASAP7_75t_L g312 ( .A(n_119), .B(n_149), .Y(n_312) );
BUFx2_ASAP7_75t_L g317 ( .A(n_119), .Y(n_317) );
AND2x2_ASAP7_75t_L g361 ( .A(n_119), .B(n_159), .Y(n_361) );
AND2x4_ASAP7_75t_L g433 ( .A(n_119), .B(n_434), .Y(n_433) );
NOR2x1_ASAP7_75t_L g445 ( .A(n_119), .B(n_215), .Y(n_445) );
OR2x6_ASAP7_75t_L g119 ( .A(n_120), .B(n_146), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_130), .B(n_142), .Y(n_120) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_128), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
AND2x6_ASAP7_75t_L g140 ( .A(n_124), .B(n_133), .Y(n_140) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g138 ( .A(n_126), .B(n_135), .Y(n_138) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx5_ASAP7_75t_L g141 ( .A(n_128), .Y(n_141) );
AND2x2_ASAP7_75t_L g134 ( .A(n_129), .B(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_129), .Y(n_234) );
AND2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
BUFx3_ASAP7_75t_L g235 ( .A(n_132), .Y(n_235) );
INVx2_ASAP7_75t_L g241 ( .A(n_133), .Y(n_241) );
AND2x4_ASAP7_75t_L g237 ( .A(n_134), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g233 ( .A(n_135), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_139), .B(n_141), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_140), .B(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_141), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_141), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_141), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_141), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_141), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_141), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_141), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_141), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_141), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_141), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_141), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_141), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_141), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_141), .A2(n_550), .B(n_551), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_142), .Y(n_151) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_142), .A2(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_142), .A2(n_493), .B(n_494), .Y(n_492) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_142), .A2(n_530), .B(n_534), .Y(n_529) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_142), .A2(n_530), .B(n_534), .Y(n_541) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x4_ASAP7_75t_L g179 ( .A(n_144), .B(n_145), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_147), .A2(n_192), .B(n_193), .Y(n_191) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_149), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g364 ( .A(n_149), .Y(n_364) );
BUFx2_ASAP7_75t_L g413 ( .A(n_149), .Y(n_413) );
INVx1_ASAP7_75t_L g435 ( .A(n_149), .Y(n_435) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_159), .Y(n_149) );
INVx3_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_150), .Y(n_401) );
AOI21x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_158), .Y(n_150) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_151), .A2(n_475), .B(n_481), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
INVx2_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_159), .B(n_212), .Y(n_216) );
INVx2_ASAP7_75t_L g301 ( .A(n_159), .Y(n_301) );
OR2x2_ASAP7_75t_L g308 ( .A(n_159), .B(n_257), .Y(n_308) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_167), .Y(n_159) );
INVx4_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
INVx3_ASAP7_75t_L g182 ( .A(n_168), .Y(n_182) );
AND2x2_ASAP7_75t_L g263 ( .A(n_169), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g297 ( .A(n_169), .B(n_260), .Y(n_297) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_180), .Y(n_169) );
AND2x2_ASAP7_75t_L g333 ( .A(n_170), .B(n_222), .Y(n_333) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g290 ( .A(n_171), .B(n_181), .Y(n_290) );
AND2x2_ASAP7_75t_L g409 ( .A(n_171), .B(n_190), .Y(n_409) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
INVx1_ASAP7_75t_L g249 ( .A(n_172), .Y(n_249) );
AND2x2_ASAP7_75t_L g305 ( .A(n_172), .B(n_181), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_172), .B(n_202), .Y(n_310) );
OR2x2_ASAP7_75t_L g373 ( .A(n_172), .B(n_190), .Y(n_373) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_172), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_179), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_179), .A2(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_SL g464 ( .A(n_179), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_179), .A2(n_485), .B(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_179), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g201 ( .A(n_180), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g250 ( .A(n_180), .Y(n_250) );
NOR2x1_ASAP7_75t_SL g180 ( .A(n_181), .B(n_190), .Y(n_180) );
AO21x1_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_181) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_223) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_182), .A2(n_514), .B(n_520), .Y(n_513) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_182), .A2(n_547), .B(n_553), .Y(n_546) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_182), .A2(n_547), .B(n_553), .Y(n_582) );
AO21x2_ASAP7_75t_L g585 ( .A1(n_182), .A2(n_514), .B(n_520), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
AND2x2_ASAP7_75t_L g218 ( .A(n_190), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_SL g276 ( .A(n_190), .Y(n_276) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_190), .B(n_202), .Y(n_286) );
OR2x2_ASAP7_75t_L g291 ( .A(n_190), .B(n_219), .Y(n_291) );
BUFx2_ASAP7_75t_L g347 ( .A(n_190), .Y(n_347) );
AND2x2_ASAP7_75t_L g383 ( .A(n_190), .B(n_262), .Y(n_383) );
AND2x2_ASAP7_75t_L g394 ( .A(n_190), .B(n_222), .Y(n_394) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_198), .Y(n_190) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_210), .B1(n_216), .B2(n_217), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_201), .A2(n_391), .B1(n_441), .B2(n_446), .Y(n_440) );
INVx4_ASAP7_75t_L g219 ( .A(n_202), .Y(n_219) );
INVx2_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_202), .Y(n_331) );
OR2x2_ASAP7_75t_L g346 ( .A(n_202), .B(n_222), .Y(n_346) );
OR2x2_ASAP7_75t_SL g372 ( .A(n_202), .B(n_373), .Y(n_372) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_211), .B(n_213), .Y(n_210) );
INVx2_ASAP7_75t_SL g253 ( .A(n_211), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_211), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g321 ( .A(n_211), .B(n_269), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_211), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_212), .Y(n_268) );
AND2x2_ASAP7_75t_L g324 ( .A(n_212), .B(n_301), .Y(n_324) );
INVx1_ASAP7_75t_L g434 ( .A(n_212), .Y(n_434) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_214), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_214), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g242 ( .A(n_215), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_216), .B(n_375), .Y(n_374) );
AOI321xp33_ASAP7_75t_L g396 ( .A1(n_217), .A2(n_298), .A3(n_366), .B1(n_397), .B2(n_398), .C(n_402), .Y(n_396) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_218), .Y(n_295) );
AND2x2_ASAP7_75t_L g320 ( .A(n_218), .B(n_249), .Y(n_320) );
AND2x2_ASAP7_75t_L g395 ( .A(n_218), .B(n_305), .Y(n_395) );
INVx1_ASAP7_75t_L g264 ( .A(n_219), .Y(n_264) );
BUFx2_ASAP7_75t_L g274 ( .A(n_219), .Y(n_274) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_219), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g319 ( .A(n_220), .Y(n_319) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
BUFx2_ASAP7_75t_L g326 ( .A(n_221), .Y(n_326) );
INVx2_ASAP7_75t_L g262 ( .A(n_222), .Y(n_262) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_222), .Y(n_285) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AOI21xp33_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_244), .B(n_247), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_225), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_242), .Y(n_226) );
INVx3_ASAP7_75t_L g269 ( .A(n_227), .Y(n_269) );
AND2x2_ASAP7_75t_L g300 ( .A(n_227), .B(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AND2x4_ASAP7_75t_L g257 ( .A(n_228), .B(n_229), .Y(n_257) );
AND2x4_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NOR2x1p5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
INVx1_ASAP7_75t_SL g425 ( .A(n_243), .Y(n_425) );
INVxp33_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_246), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g351 ( .A(n_246), .B(n_308), .Y(n_351) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
AND2x2_ASAP7_75t_L g355 ( .A(n_248), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_248), .B(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_249), .B(n_286), .Y(n_341) );
NOR4xp25_ASAP7_75t_L g436 ( .A(n_249), .B(n_280), .C(n_437), .D(n_438), .Y(n_436) );
OR2x2_ASAP7_75t_L g404 ( .A(n_250), .B(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_258), .B1(n_263), .B2(n_265), .C(n_270), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g279 ( .A(n_254), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g316 ( .A(n_255), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g336 ( .A(n_256), .Y(n_336) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx3_ASAP7_75t_L g359 ( .A(n_257), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_257), .B(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OR2x2_ASAP7_75t_L g303 ( .A(n_260), .B(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_262), .B(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx2_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_267), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g272 ( .A(n_269), .Y(n_272) );
OAI321xp33_ASAP7_75t_L g384 ( .A1(n_269), .A2(n_377), .A3(n_385), .B1(n_390), .B2(n_392), .C(n_396), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
OR2x2_ASAP7_75t_L g339 ( .A(n_272), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g439 ( .A(n_275), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_276), .B(n_319), .Y(n_318) );
NAND2xp33_ASAP7_75t_SL g419 ( .A(n_276), .B(n_290), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_292), .C(n_296), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2x1_ASAP7_75t_L g281 ( .A(n_282), .B(n_287), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g388 ( .A(n_285), .Y(n_388) );
INVx3_ASAP7_75t_L g327 ( .A(n_286), .Y(n_327) );
OR2x2_ASAP7_75t_L g430 ( .A(n_286), .B(n_304), .Y(n_430) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_288), .A2(n_372), .B1(n_374), .B2(n_376), .Y(n_371) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_SL g370 ( .A(n_291), .Y(n_370) );
OR2x2_ASAP7_75t_L g447 ( .A(n_291), .B(n_304), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_298), .B(n_302), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_300), .B(n_317), .Y(n_416) );
AND2x2_ASAP7_75t_L g422 ( .A(n_300), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g367 ( .A(n_301), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B1(n_309), .B2(n_311), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_304), .A2(n_347), .B(n_349), .C(n_351), .Y(n_348) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_307), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_307), .B(n_399), .Y(n_421) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g393 ( .A(n_310), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_312), .A2(n_344), .B(n_347), .C(n_348), .Y(n_343) );
NAND3xp33_ASAP7_75t_SL g313 ( .A(n_314), .B(n_328), .C(n_343), .Y(n_313) );
AOI222xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_320), .B2(n_321), .C1(n_322), .C2(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_317), .B(n_350), .Y(n_403) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g337 ( .A(n_324), .Y(n_337) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OR2x2_ASAP7_75t_L g442 ( .A(n_326), .B(n_359), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_327), .A2(n_418), .B1(n_420), .B2(n_422), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_334), .B1(n_338), .B2(n_341), .C(n_342), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI21xp5_ASAP7_75t_SL g402 ( .A1(n_335), .A2(n_403), .B(n_404), .Y(n_402) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g350 ( .A(n_336), .Y(n_350) );
AND2x2_ASAP7_75t_L g444 ( .A(n_336), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g428 ( .A(n_340), .Y(n_428) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g357 ( .A(n_346), .B(n_347), .Y(n_357) );
INVx1_ASAP7_75t_L g410 ( .A(n_346), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_384), .C(n_406), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B(n_360), .C(n_365), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g360 ( .A1(n_355), .A2(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI211xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B(n_371), .C(n_378), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g389 ( .A(n_372), .Y(n_389) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_373), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_375), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g437 ( .A(n_375), .Y(n_437) );
AND2x2_ASAP7_75t_L g427 ( .A(n_377), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g397 ( .A(n_379), .Y(n_397) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_393), .A2(n_427), .B1(n_429), .B2(n_431), .C(n_436), .Y(n_426) );
OAI21xp33_ASAP7_75t_SL g441 ( .A1(n_398), .A2(n_442), .B(n_443), .Y(n_441) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_417), .C(n_426), .D(n_440), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B1(n_414), .B2(n_415), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
CKINVDCx6p67_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
AND2x6_ASAP7_75t_SL g451 ( .A(n_452), .B(n_453), .Y(n_451) );
OR2x6_ASAP7_75t_SL g747 ( .A(n_452), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g757 ( .A(n_452), .B(n_453), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_452), .B(n_748), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_453), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx2_ASAP7_75t_L g751 ( .A(n_457), .Y(n_751) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_645), .Y(n_457) );
NAND3xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_557), .C(n_612), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_498), .B1(n_521), .B2(n_525), .C(n_535), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_482), .Y(n_460) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_461), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g556 ( .A(n_461), .Y(n_556) );
AND2x2_ASAP7_75t_L g601 ( .A(n_461), .B(n_538), .Y(n_601) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g589 ( .A(n_463), .Y(n_589) );
INVx1_ASAP7_75t_L g599 ( .A(n_463), .Y(n_599) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_471), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_464), .B(n_472), .Y(n_471) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_464), .A2(n_465), .B(n_471), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
OR2x2_ASAP7_75t_L g578 ( .A(n_473), .B(n_483), .Y(n_578) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_473), .B(n_524), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_473), .B(n_490), .Y(n_622) );
INVx2_ASAP7_75t_L g631 ( .A(n_473), .Y(n_631) );
AND2x2_ASAP7_75t_L g652 ( .A(n_473), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g736 ( .A(n_473), .B(n_555), .Y(n_736) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g564 ( .A(n_474), .B(n_490), .Y(n_564) );
AND2x2_ASAP7_75t_L g697 ( .A(n_474), .B(n_524), .Y(n_697) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_474), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
AND2x4_ASAP7_75t_L g651 ( .A(n_482), .B(n_652), .Y(n_651) );
AOI321xp33_ASAP7_75t_L g665 ( .A1(n_482), .A2(n_594), .A3(n_595), .B1(n_627), .B2(n_666), .C(n_669), .Y(n_665) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_490), .Y(n_482) );
BUFx3_ASAP7_75t_L g522 ( .A(n_483), .Y(n_522) );
INVx2_ASAP7_75t_L g555 ( .A(n_483), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_483), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g588 ( .A(n_483), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g621 ( .A(n_483), .Y(n_621) );
INVx5_ASAP7_75t_L g524 ( .A(n_490), .Y(n_524) );
NOR2x1_ASAP7_75t_SL g573 ( .A(n_490), .B(n_563), .Y(n_573) );
BUFx2_ASAP7_75t_L g668 ( .A(n_490), .Y(n_668) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVxp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
NOR2xp33_ASAP7_75t_SL g566 ( .A(n_500), .B(n_567), .Y(n_566) );
NOR4xp25_ASAP7_75t_L g669 ( .A(n_500), .B(n_663), .C(n_667), .D(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g707 ( .A(n_500), .Y(n_707) );
AND2x2_ASAP7_75t_L g741 ( .A(n_500), .B(n_681), .Y(n_741) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g542 ( .A(n_501), .Y(n_542) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g596 ( .A(n_502), .Y(n_596) );
OAI21x1_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_505), .B(n_509), .Y(n_502) );
INVx1_ASAP7_75t_L g510 ( .A(n_504), .Y(n_510) );
AOI33xp33_ASAP7_75t_L g737 ( .A1(n_511), .A2(n_539), .A3(n_570), .B1(n_586), .B2(n_692), .B3(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g527 ( .A(n_512), .B(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g537 ( .A(n_512), .B(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g544 ( .A(n_513), .Y(n_544) );
INVxp67_ASAP7_75t_L g625 ( .A(n_513), .Y(n_625) );
AND2x2_ASAP7_75t_L g681 ( .A(n_513), .B(n_546), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_521), .A2(n_703), .B(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
AND2x2_ASAP7_75t_L g690 ( .A(n_522), .B(n_564), .Y(n_690) );
AND3x2_ASAP7_75t_L g692 ( .A(n_522), .B(n_576), .C(n_631), .Y(n_692) );
INVx3_ASAP7_75t_SL g644 ( .A(n_523), .Y(n_644) );
INVx4_ASAP7_75t_L g538 ( .A(n_524), .Y(n_538) );
AND2x2_ASAP7_75t_L g576 ( .A(n_524), .B(n_563), .Y(n_576) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
AND2x4_ASAP7_75t_L g595 ( .A(n_528), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g658 ( .A(n_528), .B(n_546), .Y(n_658) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g628 ( .A(n_529), .Y(n_628) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_529), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_R g535 ( .A1(n_536), .A2(n_539), .B(n_543), .C(n_554), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g587 ( .A(n_538), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_538), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_538), .B(n_555), .Y(n_716) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g698 ( .A(n_540), .B(n_688), .Y(n_698) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g545 ( .A(n_541), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g567 ( .A(n_541), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g583 ( .A(n_541), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g616 ( .A(n_541), .B(n_596), .Y(n_616) );
AND2x4_ASAP7_75t_L g581 ( .A(n_542), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g605 ( .A(n_542), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g643 ( .A(n_542), .B(n_568), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g571 ( .A(n_544), .B(n_568), .Y(n_571) );
AND2x2_ASAP7_75t_L g586 ( .A(n_544), .B(n_546), .Y(n_586) );
BUFx2_ASAP7_75t_L g642 ( .A(n_544), .Y(n_642) );
AND2x2_ASAP7_75t_L g656 ( .A(n_544), .B(n_567), .Y(n_656) );
INVx2_ASAP7_75t_L g568 ( .A(n_546), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_552), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_554), .A2(n_605), .B1(n_607), .B2(n_611), .Y(n_604) );
INVx2_ASAP7_75t_SL g635 ( .A(n_554), .Y(n_635) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g610 ( .A(n_555), .B(n_563), .Y(n_610) );
INVx1_ASAP7_75t_L g717 ( .A(n_556), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_590), .C(n_604), .Y(n_557) );
OAI221xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_565), .B1(n_569), .B2(n_572), .C(n_574), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g618 ( .A(n_562), .Y(n_618) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_562), .Y(n_746) );
INVx1_ASAP7_75t_L g709 ( .A(n_564), .Y(n_709) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_564), .B(n_588), .Y(n_719) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_568), .B(n_596), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
OR2x2_ASAP7_75t_L g602 ( .A(n_570), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g680 ( .A(n_570), .Y(n_680) );
AND2x2_ASAP7_75t_L g615 ( .A(n_571), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g661 ( .A(n_573), .B(n_621), .Y(n_661) );
AND2x2_ASAP7_75t_L g738 ( .A(n_573), .B(n_736), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_579), .B1(n_586), .B2(n_587), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g597 ( .A(n_578), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx2_ASAP7_75t_L g603 ( .A(n_581), .Y(n_603) );
AND2x4_ASAP7_75t_L g627 ( .A(n_581), .B(n_628), .Y(n_627) );
OAI21xp33_ASAP7_75t_SL g657 ( .A1(n_581), .A2(n_658), .B(n_659), .Y(n_657) );
AND2x2_ASAP7_75t_L g684 ( .A(n_581), .B(n_642), .Y(n_684) );
INVx2_ASAP7_75t_L g606 ( .A(n_582), .Y(n_606) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_582), .Y(n_639) );
INVx1_ASAP7_75t_SL g663 ( .A(n_583), .Y(n_663) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g594 ( .A(n_585), .Y(n_594) );
AND2x4_ASAP7_75t_SL g688 ( .A(n_585), .B(n_606), .Y(n_688) );
AND2x2_ASAP7_75t_L g685 ( .A(n_588), .B(n_631), .Y(n_685) );
AND2x2_ASAP7_75t_L g711 ( .A(n_588), .B(n_697), .Y(n_711) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_589), .Y(n_633) );
INVx1_ASAP7_75t_L g653 ( .A(n_589), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_597), .B1(n_600), .B2(n_602), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_595), .B(n_606), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_595), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g734 ( .A(n_595), .Y(n_734) );
INVx2_ASAP7_75t_SL g659 ( .A(n_597), .Y(n_659) );
AND2x2_ASAP7_75t_L g671 ( .A(n_599), .B(n_631), .Y(n_671) );
INVx2_ASAP7_75t_L g677 ( .A(n_599), .Y(n_677) );
INVxp33_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g636 ( .A(n_602), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_605), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g727 ( .A(n_605), .Y(n_727) );
INVx1_ASAP7_75t_L g655 ( .A(n_607), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_608), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g666 ( .A(n_610), .B(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_610), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_634), .C(n_637), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B1(n_619), .B2(n_623), .C(n_626), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g732 ( .A(n_617), .Y(n_732) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g701 ( .A(n_618), .B(n_667), .Y(n_701) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g632 ( .A(n_621), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g703 ( .A(n_623), .Y(n_703) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g700 ( .A(n_624), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_625), .Y(n_706) );
OR2x2_ASAP7_75t_L g729 ( .A(n_625), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_SL g638 ( .A(n_628), .Y(n_638) );
AND2x2_ASAP7_75t_L g708 ( .A(n_628), .B(n_688), .Y(n_708) );
AND2x2_ASAP7_75t_SL g740 ( .A(n_628), .B(n_641), .Y(n_740) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g745 ( .A(n_631), .Y(n_745) );
INVx1_ASAP7_75t_L g695 ( .A(n_633), .Y(n_695) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_640), .C(n_644), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_638), .B(n_688), .Y(n_712) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_641), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g649 ( .A(n_643), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g730 ( .A(n_643), .Y(n_730) );
NAND4xp75_ASAP7_75t_L g645 ( .A(n_646), .B(n_702), .C(n_718), .D(n_739), .Y(n_645) );
NOR3x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_664), .C(n_686), .Y(n_646) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_648), .B(n_654), .C(n_657), .D(n_660), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g699 ( .A(n_650), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g724 ( .A(n_651), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_SL g713 ( .A(n_656), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_672), .Y(n_664) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_668), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_678), .B(n_682), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI322xp33_ASAP7_75t_L g704 ( .A1(n_676), .A2(n_705), .A3(n_709), .B1(n_710), .B2(n_712), .C1(n_713), .C2(n_714), .Y(n_704) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_677), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_680), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_681), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_691), .C(n_693), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_698), .B1(n_699), .B2(n_701), .Y(n_693) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_708), .Y(n_705) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_711), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g721 ( .A(n_716), .B(n_722), .Y(n_721) );
O2A1O1Ixp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B(n_725), .C(n_728), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI221xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_731), .B1(n_733), .B2(n_735), .C(n_737), .Y(n_728) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
CKINVDCx11_ASAP7_75t_R g753 ( .A(n_747), .Y(n_753) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_763), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI21xp33_ASAP7_75t_SL g772 ( .A1(n_764), .A2(n_773), .B(n_776), .Y(n_772) );
NOR2xp33_ASAP7_75t_SL g764 ( .A(n_765), .B(n_768), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
BUFx3_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
BUFx2_ASAP7_75t_R g775 ( .A(n_767), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx3_ASAP7_75t_SL g796 ( .A(n_787), .Y(n_796) );
AND2x2_ASAP7_75t_SL g787 ( .A(n_788), .B(n_789), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
endmodule