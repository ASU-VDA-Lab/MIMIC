module fake_jpeg_12333_n_386 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_54),
.Y(n_165)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_61),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_57),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_58),
.Y(n_170)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_21),
.B(n_9),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_63),
.B(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_10),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_102),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_68),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_69),
.B(n_85),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_72),
.Y(n_133)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_94),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_15),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_11),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_89),
.B(n_95),
.Y(n_166)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_17),
.B(n_14),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_108),
.Y(n_128)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_106),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_49),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_49),
.Y(n_116)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_32),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_62),
.B1(n_40),
.B2(n_44),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_127),
.A2(n_134),
.B1(n_137),
.B2(n_142),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_50),
.B1(n_17),
.B2(n_85),
.Y(n_130)
);

OA22x2_ASAP7_75t_SL g203 ( 
.A1(n_130),
.A2(n_161),
.B1(n_151),
.B2(n_127),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_40),
.B1(n_50),
.B2(n_41),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_138),
.B1(n_58),
.B2(n_79),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_40),
.B1(n_46),
.B2(n_41),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_140),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_72),
.A2(n_28),
.B1(n_46),
.B2(n_34),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_64),
.B1(n_69),
.B2(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_33),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_28),
.B1(n_34),
.B2(n_33),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_54),
.A2(n_48),
.B1(n_43),
.B2(n_35),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_143),
.A2(n_151),
.B1(n_167),
.B2(n_152),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_48),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_153),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_77),
.A2(n_43),
.B1(n_35),
.B2(n_24),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_24),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_87),
.B(n_14),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_80),
.B(n_82),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_92),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_39),
.B(n_1),
.C(n_3),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_100),
.A2(n_39),
.B1(n_1),
.B2(n_3),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_164),
.A2(n_133),
.B1(n_122),
.B2(n_155),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_57),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_167)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_101),
.C(n_71),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_172),
.B(n_191),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_175),
.A2(n_196),
.B1(n_203),
.B2(n_211),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_0),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_180),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_179),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_3),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_115),
.B(n_4),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_181),
.B(n_214),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_7),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_202),
.Y(n_239)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_143),
.A2(n_60),
.B1(n_78),
.B2(n_81),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_205),
.B1(n_220),
.B2(n_144),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_7),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_7),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_201),
.Y(n_250)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_110),
.A2(n_131),
.B1(n_121),
.B2(n_142),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_110),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_116),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_128),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_125),
.B(n_137),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_206),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_134),
.A2(n_111),
.B1(n_112),
.B2(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_111),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_207),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_212),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_158),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_207),
.Y(n_256)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_145),
.A2(n_170),
.B1(n_168),
.B2(n_146),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_210),
.B1(n_206),
.B2(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_132),
.B(n_118),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_133),
.A2(n_122),
.B(n_119),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_221),
.B(n_169),
.Y(n_234)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_117),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_147),
.B1(n_119),
.B2(n_152),
.Y(n_224)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_170),
.B1(n_162),
.B2(n_147),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_154),
.B(n_139),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_241),
.B1(n_246),
.B2(n_238),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_234),
.A2(n_259),
.B(n_250),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_197),
.A2(n_169),
.B1(n_139),
.B2(n_144),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_236),
.A2(n_256),
.B1(n_233),
.B2(n_224),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_171),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_184),
.B1(n_180),
.B2(n_188),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_175),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_197),
.A2(n_204),
.B(n_173),
.C(n_176),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_254),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_251),
.B1(n_245),
.B2(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_191),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_182),
.B(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_258),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_177),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_203),
.A2(n_189),
.B1(n_172),
.B2(n_185),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_194),
.A2(n_221),
.B(n_216),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_201),
.B(n_195),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_239),
.B(n_198),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_261),
.B(n_266),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_287),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_265),
.B1(n_277),
.B2(n_279),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_233),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_272),
.B1(n_275),
.B2(n_240),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_192),
.B1(n_241),
.B2(n_259),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_260),
.B(n_245),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_225),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_225),
.B(n_258),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_223),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_249),
.A2(n_252),
.B1(n_237),
.B2(n_255),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_250),
.C(n_249),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_257),
.C(n_244),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_256),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_288),
.B(n_290),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_231),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_231),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_226),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_288),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_293),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_298),
.B1(n_309),
.B2(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_257),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_303),
.Y(n_315)
);

OAI22x1_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_227),
.B1(n_244),
.B2(n_240),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_301),
.C(n_289),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_242),
.C(n_227),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_240),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_265),
.B1(n_263),
.B2(n_279),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_263),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_272),
.A2(n_235),
.B1(n_242),
.B2(n_269),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_268),
.C(n_273),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_316),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_267),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_280),
.C(n_282),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_318),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_287),
.C(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_324),
.B1(n_328),
.B2(n_306),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_270),
.C(n_268),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_326),
.C(n_327),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_270),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_308),
.Y(n_325)
);

INVx11_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_271),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_262),
.C(n_261),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_275),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_310),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_281),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_292),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_333),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_292),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_339),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_343),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_323),
.B(n_310),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_311),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_327),
.Y(n_352)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_309),
.A3(n_291),
.B1(n_299),
.B2(n_298),
.C1(n_311),
.C2(n_308),
.Y(n_342)
);

OAI322xp33_ASAP7_75t_L g356 ( 
.A1(n_342),
.A2(n_275),
.A3(n_284),
.B1(n_307),
.B2(n_304),
.C1(n_278),
.C2(n_276),
.Y(n_356)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_341),
.A2(n_330),
.B(n_328),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_346),
.A2(n_348),
.B(n_294),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_336),
.A2(n_321),
.B(n_329),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_322),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_353),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_345),
.C(n_338),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_286),
.Y(n_353)
);

AOI31xp67_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_332),
.A3(n_299),
.B(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_356),
.A2(n_264),
.B1(n_283),
.B2(n_285),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_334),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_344),
.B1(n_307),
.B2(n_294),
.Y(n_359)
);

AO22x1_ASAP7_75t_L g358 ( 
.A1(n_350),
.A2(n_344),
.B1(n_343),
.B2(n_333),
.Y(n_358)
);

A2O1A1Ixp33_ASAP7_75t_SL g373 ( 
.A1(n_358),
.A2(n_366),
.B(n_347),
.C(n_235),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_359),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_362),
.B(n_364),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_351),
.B1(n_348),
.B2(n_346),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_345),
.B1(n_338),
.B2(n_335),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_339),
.C(n_294),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_365),
.B(n_355),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_360),
.B(n_352),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_371),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_373),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_SL g372 ( 
.A1(n_363),
.A2(n_354),
.B(n_347),
.C(n_235),
.Y(n_372)
);

AOI31xp33_ASAP7_75t_L g377 ( 
.A1(n_372),
.A2(n_358),
.A3(n_366),
.B(n_359),
.Y(n_377)
);

NOR2x1_ASAP7_75t_L g375 ( 
.A(n_373),
.B(n_361),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_374),
.Y(n_380)
);

AOI21xp33_ASAP7_75t_L g376 ( 
.A1(n_368),
.A2(n_361),
.B(n_364),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_365),
.C(n_369),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_358),
.C(n_362),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_380),
.B(n_381),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_378),
.B(n_375),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_383),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_374),
.Y(n_386)
);


endmodule