module fake_jpeg_14891_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_49),
.Y(n_93)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_28),
.B1(n_35),
.B2(n_32),
.Y(n_99)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_15),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_25),
.Y(n_92)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_61),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_27),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_18),
.B(n_8),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_34),
.C(n_33),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_100),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_80),
.B(n_101),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_81),
.Y(n_107)
);

NAND2xp67_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_27),
.Y(n_73)
);

OR2x4_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_39),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_23),
.B1(n_29),
.B2(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_21),
.B1(n_35),
.B2(n_32),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_44),
.B1(n_36),
.B2(n_28),
.Y(n_106)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_12),
.B(n_13),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_74),
.Y(n_105)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_34),
.C(n_33),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_56),
.B1(n_46),
.B2(n_31),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_105),
.B(n_85),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_18),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_18),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_36),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_125),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_18),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_11),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_11),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_127),
.B(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_12),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_131),
.Y(n_139)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_91),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_69),
.Y(n_130)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_13),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_13),
.B1(n_39),
.B2(n_70),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_85),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_78),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_146),
.C(n_69),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_78),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_132),
.B1(n_120),
.B2(n_118),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_68),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_68),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_153),
.B(n_158),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_159),
.B(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_67),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_81),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_114),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_88),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_105),
.B(n_69),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_181),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_104),
.B1(n_135),
.B2(n_105),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_104),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_172),
.C(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_179),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_134),
.B1(n_106),
.B2(n_111),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_124),
.Y(n_172)
);

NAND2xp67_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_130),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_140),
.C(n_137),
.Y(n_197)
);

OAI22x1_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_103),
.B1(n_75),
.B2(n_76),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_108),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_136),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_108),
.B(n_128),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_158),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_SL g185 ( 
.A1(n_178),
.A2(n_139),
.A3(n_171),
.B1(n_181),
.B2(n_163),
.C1(n_170),
.C2(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_196),
.Y(n_206)
);

BUFx4f_ASAP7_75t_SL g187 ( 
.A(n_174),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_153),
.B1(n_141),
.B2(n_148),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_199),
.B1(n_183),
.B2(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_197),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_160),
.C(n_138),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_176),
.C(n_169),
.Y(n_205)
);

NOR4xp25_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_138),
.C(n_156),
.D(n_144),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_184),
.B(n_165),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_180),
.B(n_173),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_148),
.B1(n_144),
.B2(n_162),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_204),
.B1(n_196),
.B2(n_194),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_166),
.B1(n_180),
.B2(n_183),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_209),
.B(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_174),
.C(n_151),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_198),
.C(n_186),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_220),
.Y(n_227)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_190),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_219),
.A2(n_213),
.B(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_195),
.B1(n_193),
.B2(n_187),
.Y(n_220)
);

OAI321xp33_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_188),
.A3(n_139),
.B1(n_187),
.B2(n_161),
.C(n_162),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_207),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_210),
.C(n_205),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_225),
.B1(n_157),
.B2(n_145),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_228),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_202),
.C(n_161),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_226),
.A2(n_215),
.B(n_202),
.C(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_219),
.B(n_145),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.C(n_72),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_227),
.A3(n_222),
.B1(n_152),
.B2(n_128),
.C1(n_115),
.C2(n_86),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_235),
.B(n_237),
.C(n_133),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_115),
.A3(n_133),
.B1(n_79),
.B2(n_72),
.C1(n_75),
.C2(n_122),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_236),
.A2(n_230),
.B(n_233),
.C(n_116),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_116),
.C(n_122),
.Y(n_241)
);


endmodule