module fake_jpeg_17790_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_25),
.B1(n_22),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_52),
.B1(n_66),
.B2(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_56),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_25),
.B1(n_22),
.B2(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_25),
.B1(n_22),
.B2(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_64),
.B1(n_65),
.B2(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_25),
.B1(n_30),
.B2(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_24),
.B1(n_21),
.B2(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_31),
.B1(n_33),
.B2(n_18),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_34),
.C(n_28),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_45),
.B(n_41),
.C(n_40),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_97),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_74),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_79),
.B(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_26),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_94),
.C(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_26),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_98),
.B(n_20),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_95),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_60),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_41),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_19),
.B(n_24),
.C(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_19),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_29),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_105),
.B1(n_58),
.B2(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_17),
.B1(n_32),
.B2(n_16),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_58),
.B1(n_20),
.B2(n_16),
.Y(n_109)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_109),
.B1(n_123),
.B2(n_126),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_40),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_112),
.A2(n_119),
.B(n_135),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_40),
.B(n_44),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_124),
.B(n_28),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_115),
.B(n_86),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_35),
.B1(n_17),
.B2(n_32),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_32),
.B1(n_35),
.B2(n_20),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_35),
.B1(n_20),
.B2(n_29),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_74),
.B1(n_72),
.B2(n_90),
.Y(n_147)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_49),
.C(n_48),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_76),
.C(n_96),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_44),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_121),
.C(n_115),
.Y(n_177)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_159),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_88),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_148),
.B1(n_122),
.B2(n_120),
.Y(n_175)
);

AO21x2_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_92),
.B(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_92),
.B1(n_83),
.B2(n_85),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_149),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_79),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_98),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_162),
.B(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_82),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_76),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_84),
.B1(n_101),
.B2(n_77),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_84),
.B1(n_77),
.B2(n_106),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_94),
.B1(n_87),
.B2(n_86),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

AO221x1_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_74),
.B1(n_102),
.B2(n_81),
.C(n_49),
.Y(n_158)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_160),
.B(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_49),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_113),
.B(n_48),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_133),
.C(n_118),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_11),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_168),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_114),
.A3(n_134),
.B1(n_119),
.B2(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_137),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_114),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_177),
.C(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_135),
.B(n_120),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_176),
.B(n_189),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_191),
.B1(n_193),
.B2(n_200),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_121),
.B(n_125),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_129),
.C(n_122),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_81),
.B1(n_35),
.B2(n_116),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_194),
.B1(n_159),
.B2(n_157),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_28),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_35),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_200),
.B(n_158),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_148),
.A2(n_116),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_149),
.A2(n_116),
.B1(n_2),
.B2(n_4),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_8),
.C(n_14),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_8),
.C(n_13),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_166),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_173),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_162),
.B1(n_142),
.B2(n_154),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_226),
.B1(n_227),
.B2(n_199),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_210),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_230),
.B(n_196),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_143),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_137),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_177),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_191),
.B1(n_194),
.B2(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_229),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_174),
.A2(n_145),
.B(n_144),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_184),
.B(n_188),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_167),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_167),
.B1(n_5),
.B2(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_15),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_189),
.B(n_176),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_234),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_236),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_250),
.B(n_212),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_172),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_219),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_178),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_208),
.B(n_187),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_245),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_178),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_197),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_249),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_204),
.B(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_192),
.C(n_185),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_192),
.C(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_268),
.B(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_203),
.B1(n_218),
.B2(n_207),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_266),
.B1(n_269),
.B2(n_274),
.Y(n_289)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_238),
.B1(n_253),
.B2(n_237),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_213),
.B(n_225),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_233),
.A2(n_206),
.B1(n_215),
.B2(n_226),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_228),
.B(n_227),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_209),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_236),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_282),
.C(n_286),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_273),
.B1(n_266),
.B2(n_269),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_284),
.B1(n_263),
.B2(n_261),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_252),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_210),
.B1(n_209),
.B2(n_231),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_261),
.B(n_242),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_234),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_287),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_293),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_257),
.B1(n_259),
.B2(n_232),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_267),
.B1(n_259),
.B2(n_249),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_295),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_285),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_300),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_248),
.C(n_217),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_299),
.C(n_280),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_2),
.C(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_15),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_302),
.B(n_304),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_278),
.A2(n_15),
.B(n_6),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_287),
.B(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_312),
.C(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_308),
.B(n_292),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_286),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_7),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_7),
.B(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_298),
.B(n_292),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_7),
.Y(n_312)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_319),
.C(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_320),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_307),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_310),
.B1(n_315),
.B2(n_312),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_315),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_306),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_319),
.B(n_322),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_324),
.B(n_328),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_326),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);


endmodule