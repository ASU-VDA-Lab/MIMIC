module fake_jpeg_1115_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_10),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_59),
.Y(n_113)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_7),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_25),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_20),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_73),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_77),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_22),
.B1(n_21),
.B2(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_76),
.A2(n_90),
.B1(n_101),
.B2(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_81),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_33),
.B1(n_29),
.B2(n_38),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_107),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_28),
.B1(n_33),
.B2(n_24),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_34),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_94),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_37),
.B1(n_30),
.B2(n_38),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_51),
.B1(n_61),
.B2(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_111),
.B1(n_112),
.B2(n_12),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_54),
.B(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_96),
.B(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_35),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_35),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_15),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_29),
.B1(n_39),
.B2(n_32),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_65),
.B1(n_23),
.B2(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_43),
.B1(n_32),
.B2(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_43),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_45),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_62),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_119),
.B(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_135),
.Y(n_162)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_149),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_147),
.B1(n_149),
.B2(n_156),
.Y(n_160)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_151),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_91),
.A2(n_15),
.B1(n_16),
.B2(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_145),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_107),
.A2(n_16),
.B1(n_80),
.B2(n_111),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_113),
.B(n_87),
.C(n_118),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_105),
.B(n_102),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_101),
.B1(n_90),
.B2(n_100),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_164),
.A2(n_169),
.B1(n_191),
.B2(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_84),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_176),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_106),
.C(n_80),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_172),
.C(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_76),
.B1(n_98),
.B2(n_116),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_106),
.C(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_187),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_116),
.B1(n_102),
.B2(n_117),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_175),
.A2(n_143),
.B1(n_154),
.B2(n_155),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_71),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_98),
.B1(n_117),
.B2(n_153),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_138),
.B1(n_123),
.B2(n_121),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_131),
.C(n_120),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_129),
.Y(n_204)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_135),
.Y(n_182)
);

NAND2x1p5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_126),
.B(n_122),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_125),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_152),
.C(n_158),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_182),
.C(n_168),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_128),
.A2(n_139),
.B1(n_140),
.B2(n_119),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_132),
.B(n_137),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_145),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_151),
.B1(n_142),
.B2(n_134),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_196),
.B(n_212),
.Y(n_254)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_214),
.B(n_186),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_221),
.B1(n_159),
.B2(n_225),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_204),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_211),
.C(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_182),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_187),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_164),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_169),
.A2(n_161),
.B(n_190),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_224),
.B(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_174),
.C(n_166),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_177),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_160),
.B1(n_186),
.B2(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_159),
.B(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_228),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_181),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_204),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_191),
.B1(n_178),
.B2(n_187),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_223),
.B1(n_203),
.B2(n_199),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_243),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_159),
.B(n_227),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_204),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_211),
.B1(n_205),
.B2(n_199),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_220),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_207),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_229),
.B1(n_213),
.B2(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_235),
.B1(n_243),
.B2(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_214),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_215),
.C(n_206),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_272),
.C(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_219),
.B1(n_222),
.B2(n_217),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_224),
.B(n_198),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_276),
.B(n_241),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_273),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_253),
.B(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_236),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_240),
.C(n_251),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_255),
.C(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_239),
.C(n_231),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_238),
.C(n_246),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_238),
.C(n_246),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_248),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_291),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_232),
.A3(n_240),
.B1(n_233),
.B2(n_234),
.C1(n_251),
.C2(n_242),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_276),
.B1(n_266),
.B2(n_261),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_275),
.C(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_275),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_258),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_258),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_299),
.B(n_305),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_279),
.A2(n_261),
.B1(n_271),
.B2(n_274),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_279),
.B1(n_265),
.B2(n_262),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_284),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_293),
.C(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_310),
.B(n_318),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_257),
.B(n_273),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_300),
.B(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_233),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_307),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_297),
.B(n_281),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_317),
.B(n_282),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_327),
.B(n_310),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_303),
.C(n_302),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_324),
.B(n_325),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_323),
.A2(n_314),
.B1(n_270),
.B2(n_259),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_263),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_315),
.B(n_308),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_328),
.A2(n_329),
.B(n_326),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_308),
.B(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_322),
.B(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_330),
.C(n_316),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_331),
.B(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_338),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_337),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_339),
.Y(n_343)
);


endmodule