module fake_netlist_6_2366_n_1816 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1816);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1816;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_41),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_40),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_58),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_51),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_26),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_1),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_38),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_59),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_36),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_45),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_72),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_32),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_6),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_71),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_60),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_40),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_127),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_28),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_123),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_87),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_111),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_112),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_10),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_126),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_25),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_66),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_85),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_51),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_22),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_24),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_13),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_0),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_31),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_82),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_102),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_30),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_107),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_62),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_139),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_47),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_34),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_81),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_133),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_113),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_54),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_150),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_74),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_109),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_9),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_19),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_132),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_4),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_70),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_18),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_106),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_131),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_15),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_104),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_38),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_52),
.Y(n_261)
);

BUFx8_ASAP7_75t_SL g262 ( 
.A(n_53),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_147),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_37),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_152),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_33),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_73),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_101),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_92),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_110),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_156),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_44),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_144),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_69),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_151),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_20),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_100),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_45),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_96),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_124),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_42),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_158),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_159),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_64),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_68),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_22),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_52),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_11),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_136),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_93),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_84),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_129),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_76),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_19),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_25),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_79),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_137),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_142),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_20),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_94),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_37),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_12),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_34),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_119),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_134),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_77),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_57),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_33),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_215),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_215),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_262),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_215),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_169),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_215),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_164),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_215),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_215),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_234),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_215),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_166),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_166),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_161),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_166),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_166),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_173),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_161),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_162),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_290),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_190),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_221),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_312),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_162),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_197),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_221),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_221),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_167),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_167),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_217),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_198),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_173),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_171),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_206),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_185),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_189),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_206),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_309),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_219),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_200),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_202),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_203),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_208),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_232),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_196),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_245),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_268),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_247),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_248),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_252),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_254),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_196),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_205),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_211),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_299),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_271),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_299),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_261),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_264),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_178),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_171),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_265),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_271),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_212),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_276),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_271),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_172),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_289),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_348),
.B(n_207),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_383),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_328),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_207),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_168),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_326),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_346),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_192),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_351),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_192),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_236),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_353),
.B(n_224),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_358),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_335),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_336),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_375),
.B(n_209),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_334),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_320),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_168),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_337),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_345),
.B(n_242),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_L g442 ( 
.A1(n_324),
.A2(n_228),
.B1(n_313),
.B2(n_183),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_321),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_368),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_224),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_342),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_343),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_354),
.B(n_314),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_344),
.B(n_175),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_344),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_340),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_321),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_340),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_349),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_354),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_369),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_323),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_323),
.A2(n_295),
.B(n_292),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_349),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_370),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_347),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_325),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_347),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_325),
.B(n_314),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_381),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_350),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_327),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_327),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_470),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_440),
.B(n_375),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_400),
.B(n_382),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_399),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_400),
.B(n_393),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_339),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_408),
.B(n_371),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_470),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_440),
.B(n_322),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_331),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_409),
.B(n_363),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_419),
.B(n_331),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_410),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_461),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_402),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_418),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_339),
.Y(n_503)
);

INVxp33_ASAP7_75t_SL g504 ( 
.A(n_444),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_461),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_415),
.B(n_359),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_398),
.B(n_222),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_405),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_427),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_429),
.B(n_163),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_411),
.B(n_165),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_398),
.A2(n_297),
.B1(n_305),
.B2(n_330),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_458),
.B(n_225),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_445),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_461),
.A2(n_330),
.B1(n_357),
.B2(n_244),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_421),
.B(n_359),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_411),
.B(n_417),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_443),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_411),
.B(n_417),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_427),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_443),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_458),
.B(n_230),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_459),
.B(n_444),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_455),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_463),
.B(n_189),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_445),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_463),
.B(n_357),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_455),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_417),
.B(n_231),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_429),
.A2(n_278),
.B1(n_277),
.B2(n_279),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

AND2x2_ASAP7_75t_SL g543 ( 
.A(n_461),
.B(n_185),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_461),
.A2(n_185),
.B1(n_244),
.B2(n_275),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_446),
.B(n_238),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_461),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_435),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_446),
.B(n_240),
.Y(n_550)
);

INVx8_ASAP7_75t_L g551 ( 
.A(n_467),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_451),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_465),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_446),
.B(n_436),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_436),
.B(n_452),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_431),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_471),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g565 ( 
.A(n_467),
.B(n_372),
.C(n_367),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_468),
.B(n_233),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_452),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_468),
.A2(n_233),
.B1(n_307),
.B2(n_274),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_435),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_406),
.B(n_241),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_471),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_430),
.B(n_274),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_471),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_430),
.B(n_307),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_418),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_454),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_403),
.Y(n_579)
);

OA22x2_ASAP7_75t_L g580 ( 
.A1(n_406),
.A2(n_450),
.B1(n_420),
.B2(n_372),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_403),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_467),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_418),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_454),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_448),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_435),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_442),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_412),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_437),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_430),
.B(n_175),
.Y(n_592)
);

INVxp33_ASAP7_75t_L g593 ( 
.A(n_406),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_412),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_406),
.B(n_181),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_406),
.B(n_181),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_413),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_454),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_467),
.A2(n_185),
.B1(n_201),
.B2(n_244),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_413),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_414),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_438),
.Y(n_603)
);

BUFx4f_ASAP7_75t_L g604 ( 
.A(n_420),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_437),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_414),
.B(n_423),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_420),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_454),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_401),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_438),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_401),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_438),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_423),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_454),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_426),
.B(n_201),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_437),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_420),
.A2(n_174),
.B(n_170),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_437),
.B(n_209),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_426),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_420),
.A2(n_201),
.B1(n_275),
.B2(n_244),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_532),
.B(n_428),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_567),
.B(n_447),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_478),
.B(n_367),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_497),
.A2(n_450),
.B1(n_193),
.B2(n_301),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_567),
.B(n_447),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_527),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_527),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_544),
.B(n_246),
.Y(n_629)
);

AND2x4_ASAP7_75t_SL g630 ( 
.A(n_564),
.B(n_448),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_527),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_580),
.Y(n_632)
);

O2A1O1Ixp5_ASAP7_75t_L g633 ( 
.A1(n_560),
.A2(n_450),
.B(n_176),
.C(n_263),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_520),
.Y(n_634)
);

BUFx12f_ASAP7_75t_SL g635 ( 
.A(n_514),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_580),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_R g637 ( 
.A(n_495),
.B(n_449),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_497),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_520),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_558),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_580),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_479),
.B(n_249),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_600),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_497),
.B(n_188),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_520),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_525),
.B(n_438),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_503),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_543),
.B(n_447),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_543),
.B(n_447),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_474),
.A2(n_447),
.B1(n_255),
.B2(n_310),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_543),
.B(n_201),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_506),
.B(n_275),
.Y(n_654)
);

AND2x6_ASAP7_75t_SL g655 ( 
.A(n_514),
.B(n_374),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_522),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_607),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_494),
.B(n_438),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_479),
.B(n_251),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_486),
.B(n_438),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_522),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_551),
.B(n_256),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_472),
.B(n_438),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_579),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_522),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_477),
.A2(n_308),
.B1(n_306),
.B2(n_302),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_184),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_506),
.A2(n_450),
.B1(n_191),
.B2(n_298),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_492),
.Y(n_669)
);

BUFx4_ASAP7_75t_L g670 ( 
.A(n_504),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_506),
.B(n_275),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_472),
.B(n_438),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_512),
.B(n_431),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_547),
.B(n_194),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_512),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_551),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_547),
.A2(n_450),
.B1(n_281),
.B2(n_259),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_528),
.B(n_208),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_516),
.B(n_565),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_482),
.B(n_439),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_582),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_521),
.B(n_531),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_482),
.B(n_439),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_582),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_535),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_508),
.B(n_439),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_473),
.B(n_507),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_547),
.A2(n_199),
.B1(n_287),
.B2(n_204),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_604),
.B(n_439),
.Y(n_690)
);

INVx8_ASAP7_75t_L g691 ( 
.A(n_514),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_561),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_565),
.A2(n_374),
.B(n_397),
.C(n_394),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_535),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_524),
.B(n_184),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_536),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_528),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_480),
.B(n_516),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_516),
.B(n_439),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_516),
.B(n_439),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_604),
.B(n_439),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_553),
.B(n_208),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_536),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_536),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_595),
.A2(n_376),
.B(n_397),
.C(n_394),
.Y(n_706)
);

NAND2x1_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_610),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_596),
.A2(n_378),
.B(n_390),
.C(n_387),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_571),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_541),
.A2(n_376),
.B(n_378),
.C(n_379),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_584),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_571),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_604),
.A2(n_216),
.B1(n_227),
.B2(n_229),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_568),
.B(n_379),
.C(n_377),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_572),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_583),
.B(n_439),
.Y(n_716)
);

AO221x1_ASAP7_75t_L g717 ( 
.A1(n_478),
.A2(n_239),
.B1(n_386),
.B2(n_377),
.C(n_390),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_583),
.B(n_464),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_540),
.B(n_464),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_583),
.B(n_464),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_590),
.B(n_386),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_546),
.B(n_464),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_587),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_571),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_550),
.B(n_186),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_592),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_514),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_594),
.B(n_464),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_597),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_597),
.B(n_601),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_601),
.B(n_464),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_514),
.A2(n_187),
.B1(n_183),
.B2(n_182),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_583),
.B(n_464),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_551),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_602),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_602),
.B(n_464),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_541),
.B(n_466),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_484),
.B(n_186),
.Y(n_739)
);

BUFx6f_ASAP7_75t_SL g740 ( 
.A(n_587),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_613),
.B(n_466),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_551),
.B(n_267),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_519),
.B(n_304),
.C(n_266),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_609),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_523),
.B(n_566),
.C(n_534),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_617),
.A2(n_177),
.B1(n_318),
.B2(n_187),
.Y(n_746)
);

BUFx10_ASAP7_75t_L g747 ( 
.A(n_619),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_619),
.B(n_609),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_614),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_614),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_487),
.A2(n_387),
.B(n_392),
.C(n_457),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_609),
.B(n_466),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_611),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_611),
.B(n_466),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_611),
.B(n_466),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_481),
.B(n_466),
.Y(n_757)
);

AND2x6_ASAP7_75t_SL g758 ( 
.A(n_589),
.B(n_392),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_578),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_481),
.B(n_466),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_481),
.B(n_466),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_481),
.B(n_483),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_591),
.B(n_355),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_591),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_483),
.B(n_496),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_618),
.B(n_589),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_574),
.B(n_235),
.C(n_226),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_487),
.A2(n_434),
.B(n_462),
.C(n_457),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_501),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_483),
.B(n_456),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_483),
.B(n_456),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_614),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_578),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_586),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_496),
.B(n_456),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_599),
.A2(n_253),
.B1(n_316),
.B2(n_243),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_496),
.B(n_456),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_576),
.B(n_243),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_496),
.B(n_456),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_586),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_491),
.A2(n_517),
.B(n_542),
.C(n_537),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_605),
.B(n_220),
.C(n_213),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_617),
.A2(n_273),
.B1(n_300),
.B2(n_294),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_501),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_620),
.B(n_270),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_683),
.B(n_605),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_627),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_683),
.B(n_616),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_692),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_626),
.B(n_616),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_626),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_638),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_628),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_640),
.B(n_569),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_631),
.Y(n_795)
);

INVx6_ASAP7_75t_L g796 ( 
.A(n_747),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_653),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_751),
.B(n_569),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_657),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_773),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_673),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_698),
.B(n_569),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_637),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_617),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_648),
.B(n_569),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_632),
.B(n_581),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_646),
.A2(n_610),
.B(n_554),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_664),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_695),
.B(n_214),
.C(n_210),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_679),
.B(n_675),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_774),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_691),
.B(n_623),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_766),
.A2(n_689),
.B1(n_641),
.B2(n_636),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_643),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_654),
.A2(n_499),
.B(n_491),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_726),
.B(n_688),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_697),
.B(n_469),
.Y(n_818)
);

NOR2x1p5_ASAP7_75t_L g819 ( 
.A(n_764),
.B(n_172),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_695),
.B(n_581),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_630),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_725),
.B(n_581),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_721),
.B(n_355),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_725),
.B(n_581),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_677),
.B(n_603),
.Y(n_825)
);

AND2x2_ASAP7_75t_SL g826 ( 
.A(n_766),
.B(n_615),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_744),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_688),
.B(n_603),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_682),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_637),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_677),
.Y(n_831)
);

AND2x4_ASAP7_75t_SL g832 ( 
.A(n_623),
.B(n_209),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_744),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_703),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_689),
.A2(n_668),
.B1(n_678),
.B2(n_624),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_735),
.B(n_603),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_685),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_784),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_654),
.A2(n_500),
.B(n_499),
.Y(n_839)
);

AND2x6_ASAP7_75t_L g840 ( 
.A(n_680),
.B(n_603),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_677),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_669),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_677),
.Y(n_843)
);

NOR2x1p5_ASAP7_75t_L g844 ( 
.A(n_723),
.B(n_179),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_624),
.A2(n_537),
.B1(n_500),
.B2(n_513),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_680),
.B(n_612),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_745),
.B(n_612),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_700),
.B(n_711),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_622),
.B(n_501),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_634),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_784),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_622),
.B(n_513),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_668),
.B(n_501),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_778),
.B(n_727),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_678),
.A2(n_610),
.B1(n_554),
.B2(n_562),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_639),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_645),
.Y(n_857)
);

INVx3_ASAP7_75t_SL g858 ( 
.A(n_623),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_670),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_719),
.A2(n_610),
.B(n_554),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_656),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_721),
.B(n_356),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_729),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_739),
.A2(n_533),
.B1(n_515),
.B2(n_517),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_778),
.B(n_515),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_738),
.B(n_526),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_759),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_784),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_661),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_747),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_730),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_754),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_748),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_SL g874 ( 
.A(n_635),
.B(n_282),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_739),
.B(n_237),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_665),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_748),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_621),
.B(n_526),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_667),
.B(n_237),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_667),
.B(n_529),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_784),
.B(n_734),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_734),
.B(n_501),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_676),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_727),
.Y(n_884)
);

BUFx4f_ASAP7_75t_L g885 ( 
.A(n_691),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_763),
.B(n_356),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_767),
.B(n_529),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_660),
.B(n_533),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_699),
.B(n_577),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_644),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_686),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_740),
.Y(n_892)
);

AND2x6_ASAP7_75t_L g893 ( 
.A(n_658),
.B(n_539),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_652),
.B(n_539),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_694),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_696),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_644),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_652),
.B(n_542),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_663),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_642),
.A2(n_557),
.B1(n_552),
.B2(n_555),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_672),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_671),
.B(n_552),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_763),
.B(n_361),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_681),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_684),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_704),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_728),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_701),
.B(n_577),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_671),
.B(n_555),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_758),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_706),
.B(n_557),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_706),
.B(n_562),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_SL g913 ( 
.A(n_732),
.B(n_180),
.C(n_182),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_783),
.B(n_577),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_732),
.A2(n_563),
.B1(n_258),
.B2(n_237),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_714),
.B(n_258),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_649),
.B(n_577),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_731),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_736),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_708),
.A2(n_563),
.B(n_511),
.C(n_575),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_659),
.A2(n_608),
.B1(n_598),
.B2(n_575),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_708),
.B(n_511),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_763),
.B(n_258),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_717),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_644),
.A2(n_674),
.B1(n_649),
.B2(n_650),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_769),
.B(n_518),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_743),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_705),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_691),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_716),
.B(n_718),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_709),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_737),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_625),
.B(n_518),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_644),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_722),
.B(n_687),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_655),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_644),
.B(n_530),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_674),
.B(n_530),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_674),
.A2(n_608),
.B1(n_598),
.B2(n_570),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_746),
.B(n_651),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_768),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_712),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_740),
.Y(n_943)
);

OAI22xp33_ASAP7_75t_L g944 ( 
.A1(n_650),
.A2(n_318),
.B1(n_313),
.B2(n_284),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_782),
.B(n_361),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_724),
.Y(n_946)
);

OR2x2_ASAP7_75t_SL g947 ( 
.A(n_746),
.B(n_364),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_674),
.B(n_545),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_674),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_749),
.B(n_577),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_750),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_772),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_707),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_741),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_666),
.B(n_218),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_625),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_762),
.B(n_545),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_765),
.B(n_549),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_776),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_690),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_777),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_781),
.B(n_549),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_753),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_755),
.B(n_585),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_737),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_SL g966 ( 
.A1(n_713),
.A2(n_303),
.B1(n_250),
.B2(n_257),
.Y(n_966)
);

NAND2x1p5_ASAP7_75t_L g967 ( 
.A(n_716),
.B(n_718),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_781),
.B(n_556),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_741),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_756),
.B(n_585),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_835),
.A2(n_693),
.B1(n_720),
.B2(n_733),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_817),
.B(n_690),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_842),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_817),
.B(n_693),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_871),
.B(n_770),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_821),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_875),
.A2(n_296),
.B(n_260),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_789),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_814),
.B(n_771),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_940),
.A2(n_633),
.B(n_629),
.C(n_710),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_854),
.B(n_702),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_854),
.A2(n_715),
.B(n_752),
.C(n_702),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_SL g983 ( 
.A(n_956),
.B(n_223),
.C(n_319),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_847),
.A2(n_775),
.B(n_761),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_L g985 ( 
.A1(n_879),
.A2(n_280),
.B(n_283),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_792),
.B(n_865),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_944),
.A2(n_785),
.B(n_662),
.C(n_742),
.Y(n_987)
);

AOI21xp33_ASAP7_75t_L g988 ( 
.A1(n_944),
.A2(n_760),
.B(n_720),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_891),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_929),
.B(n_733),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_801),
.B(n_364),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_841),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_935),
.A2(n_757),
.B(n_777),
.Y(n_993)
);

AO21x2_ASAP7_75t_L g994 ( 
.A1(n_917),
.A2(n_849),
.B(n_914),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_887),
.A2(n_779),
.B(n_757),
.C(n_573),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_853),
.A2(n_585),
.B(n_588),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_792),
.B(n_556),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_810),
.B(n_253),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_812),
.B(n_365),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_853),
.A2(n_585),
.B(n_588),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_860),
.A2(n_585),
.B(n_588),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_887),
.A2(n_559),
.B(n_317),
.C(n_315),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_913),
.A2(n_282),
.B1(n_315),
.B2(n_316),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_865),
.A2(n_559),
.B(n_317),
.C(n_288),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_L g1005 ( 
.A(n_858),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_888),
.A2(n_588),
.B(n_548),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_808),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_789),
.B(n_285),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_834),
.A2(n_428),
.B(n_432),
.C(n_434),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_SL g1010 ( 
.A(n_831),
.B(n_272),
.Y(n_1010)
);

AOI221x1_ASAP7_75t_L g1011 ( 
.A1(n_933),
.A2(n_462),
.B1(n_453),
.B2(n_441),
.C(n_432),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_828),
.B(n_485),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_826),
.A2(n_282),
.B1(n_293),
.B2(n_291),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_828),
.B(n_485),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_834),
.B(n_286),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_807),
.A2(n_476),
.B(n_475),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_959),
.B(n_830),
.Y(n_1017)
);

OAI22x1_ASAP7_75t_L g1018 ( 
.A1(n_910),
.A2(n_311),
.B1(n_366),
.B2(n_365),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_791),
.B(n_488),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_791),
.B(n_488),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_818),
.B(n_366),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_841),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_814),
.B(n_489),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_SL g1024 ( 
.A1(n_933),
.A2(n_489),
.B(n_490),
.C(n_510),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_826),
.A2(n_927),
.B1(n_924),
.B2(n_787),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_841),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_884),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_884),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_823),
.B(n_441),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_831),
.B(n_490),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_848),
.B(n_502),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_829),
.B(n_502),
.Y(n_1032)
);

AND2x6_ASAP7_75t_L g1033 ( 
.A(n_925),
.B(n_475),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_822),
.A2(n_588),
.B(n_548),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_951),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_831),
.B(n_505),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_890),
.B(n_475),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_786),
.A2(n_453),
.B(n_509),
.C(n_505),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_837),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_831),
.B(n_510),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_928),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_955),
.B(n_509),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_874),
.B(n_347),
.C(n_352),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_803),
.B(n_0),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_928),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_SL g1046 ( 
.A(n_821),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_809),
.A2(n_352),
.B(n_384),
.C(n_391),
.Y(n_1047)
);

HAxp5_ASAP7_75t_L g1048 ( 
.A(n_844),
.B(n_1),
.CON(n_1048),
.SN(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_892),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_843),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_804),
.A2(n_498),
.B1(n_493),
.B2(n_476),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_886),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_863),
.B(n_498),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_797),
.B(n_493),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_812),
.B(n_476),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_843),
.B(n_493),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_793),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_824),
.A2(n_588),
.B(n_548),
.Y(n_1058)
);

CKINVDCx6p67_ASAP7_75t_R g1059 ( 
.A(n_858),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_943),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_786),
.A2(n_788),
.B(n_916),
.C(n_941),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_873),
.A2(n_352),
.B(n_384),
.C(n_391),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_843),
.A2(n_548),
.B(n_418),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_788),
.A2(n_384),
.B(n_391),
.C(n_395),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_812),
.B(n_115),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_870),
.B(n_2),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_SL g1067 ( 
.A1(n_847),
.A2(n_395),
.B(n_424),
.C(n_422),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_843),
.A2(n_548),
.B(n_418),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_799),
.B(n_548),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_946),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_868),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_795),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_820),
.A2(n_418),
.B(n_424),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_965),
.B(n_425),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_823),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_932),
.B(n_395),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_946),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_915),
.A2(n_425),
.B(n_424),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_932),
.B(n_425),
.Y(n_1079)
);

CKINVDCx8_ASAP7_75t_R g1080 ( 
.A(n_936),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_947),
.A2(n_425),
.B1(n_424),
.B2(n_422),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_862),
.B(n_2),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_960),
.B(n_418),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_923),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_859),
.A2(n_915),
.B1(n_966),
.B2(n_796),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_914),
.A2(n_418),
.B(n_424),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_899),
.B(n_425),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_868),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_862),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_867),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_872),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_901),
.B(n_422),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_960),
.B(n_422),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_904),
.B(n_422),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_886),
.Y(n_1095)
);

BUFx4f_ASAP7_75t_L g1096 ( 
.A(n_796),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_796),
.B(n_3),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_885),
.B(n_154),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_855),
.A2(n_416),
.B(n_401),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_815),
.B(n_3),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_877),
.A2(n_416),
.B(n_401),
.C(n_13),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_905),
.B(n_416),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_960),
.B(n_416),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_903),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_907),
.B(n_416),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_918),
.B(n_401),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_961),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_945),
.B(n_5),
.C(n_7),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_945),
.B(n_7),
.C(n_14),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_960),
.B(n_885),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_880),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_949),
.A2(n_148),
.B(n_141),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_794),
.A2(n_138),
.B(n_130),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_850),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_SL g1115 ( 
.A(n_890),
.B(n_21),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_949),
.B(n_114),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_819),
.B(n_105),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_805),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_949),
.A2(n_99),
.B(n_90),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_980),
.A2(n_802),
.B(n_794),
.Y(n_1120)
);

AO21x1_ASAP7_75t_L g1121 ( 
.A1(n_981),
.A2(n_849),
.B(n_930),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1016),
.A2(n_970),
.B(n_964),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1086),
.A2(n_970),
.B(n_964),
.Y(n_1123)
);

AOI221x1_ASAP7_75t_L g1124 ( 
.A1(n_982),
.A2(n_816),
.B1(n_839),
.B2(n_922),
.C(n_912),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_973),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1007),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1048),
.B(n_832),
.Y(n_1127)
);

AOI31xp67_ASAP7_75t_L g1128 ( 
.A1(n_972),
.A2(n_802),
.A3(n_864),
.B(n_900),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1011),
.A2(n_911),
.A3(n_968),
.B(n_962),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1001),
.A2(n_920),
.B(n_908),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1012),
.A2(n_827),
.B(n_833),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1014),
.A2(n_833),
.B(n_882),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1017),
.B(n_832),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_989),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1028),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_987),
.A2(n_882),
.B(n_851),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1111),
.A2(n_806),
.B1(n_790),
.B2(n_919),
.C(n_866),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_988),
.A2(n_825),
.B(n_881),
.Y(n_1138)
);

AOI221x1_ASAP7_75t_L g1139 ( 
.A1(n_971),
.A2(n_937),
.B1(n_938),
.B2(n_948),
.C(n_878),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_974),
.B(n_798),
.Y(n_1140)
);

AO32x2_ASAP7_75t_L g1141 ( 
.A1(n_971),
.A2(n_893),
.A3(n_852),
.B1(n_967),
.B2(n_930),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_996),
.A2(n_889),
.B(n_908),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1039),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1118),
.B(n_963),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1034),
.A2(n_881),
.B(n_889),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_978),
.B(n_790),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1113),
.A2(n_890),
.B(n_897),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1000),
.A2(n_958),
.B(n_957),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1104),
.B(n_806),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1096),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1118),
.B(n_963),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1061),
.B(n_846),
.C(n_921),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_993),
.A2(n_851),
.B(n_926),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_975),
.B(n_969),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1025),
.B(n_961),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_975),
.B(n_840),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_983),
.A2(n_846),
.B(n_967),
.C(n_836),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1058),
.A2(n_825),
.B(n_950),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1101),
.A2(n_902),
.A3(n_909),
.B(n_894),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_979),
.A2(n_1072),
.B1(n_1057),
.B2(n_1090),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1042),
.B(n_840),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1091),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_1065),
.B(n_1055),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1107),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1099),
.A2(n_950),
.B(n_939),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_984),
.A2(n_898),
.B(n_845),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1029),
.B(n_811),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1050),
.Y(n_1168)
);

OAI21xp33_ASAP7_75t_L g1169 ( 
.A1(n_1008),
.A2(n_954),
.B(n_813),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_988),
.A2(n_893),
.B(n_845),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1031),
.A2(n_953),
.B(n_868),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_991),
.B(n_840),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_994),
.A2(n_953),
.B(n_890),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_SL g1174 ( 
.A(n_1050),
.B(n_897),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1052),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1096),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1114),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_SL g1178 ( 
.A1(n_1023),
.A2(n_800),
.B(n_883),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_984),
.A2(n_952),
.B(n_838),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1032),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1110),
.B(n_838),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1035),
.B(n_840),
.Y(n_1182)
);

AO32x2_ASAP7_75t_L g1183 ( 
.A1(n_1085),
.A2(n_893),
.A3(n_852),
.B1(n_934),
.B2(n_897),
.Y(n_1183)
);

O2A1O1Ixp5_ASAP7_75t_SL g1184 ( 
.A1(n_1083),
.A2(n_852),
.B(n_893),
.C(n_27),
.Y(n_1184)
);

CKINVDCx16_ASAP7_75t_R g1185 ( 
.A(n_1046),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1054),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1073),
.A2(n_895),
.B(n_942),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_992),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1006),
.A2(n_857),
.B(n_856),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1079),
.A2(n_896),
.B(n_861),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_992),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1076),
.B(n_852),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1076),
.B(n_852),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1079),
.A2(n_869),
.B(n_931),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_977),
.A2(n_934),
.B(n_897),
.C(n_906),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1087),
.A2(n_1092),
.B(n_1094),
.Y(n_1196)
);

AO21x2_ASAP7_75t_L g1197 ( 
.A1(n_994),
.A2(n_876),
.B(n_893),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1013),
.A2(n_934),
.B(n_953),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_997),
.A2(n_953),
.B(n_934),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1075),
.B(n_23),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1089),
.B(n_23),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_992),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1084),
.B(n_24),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_985),
.A2(n_27),
.B(n_29),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1004),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1021),
.B(n_35),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1108),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1095),
.B(n_39),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1065),
.B(n_43),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_995),
.A2(n_55),
.B(n_88),
.Y(n_1210)
);

CKINVDCx11_ASAP7_75t_R g1211 ( 
.A(n_1080),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_976),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1062),
.A2(n_65),
.B(n_56),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_SL g1214 ( 
.A1(n_1117),
.A2(n_46),
.B(n_47),
.Y(n_1214)
);

OA22x2_ASAP7_75t_L g1215 ( 
.A1(n_1018),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_990),
.B(n_48),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1027),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_990),
.B(n_49),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1005),
.Y(n_1219)
);

NOR4xp25_ASAP7_75t_L g1220 ( 
.A(n_1109),
.B(n_50),
.C(n_53),
.D(n_1003),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1005),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1055),
.A2(n_1100),
.B1(n_1002),
.B2(n_1051),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1053),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1059),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1082),
.B(n_1070),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1087),
.A2(n_1102),
.B(n_1094),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1092),
.A2(n_1102),
.B(n_1105),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1049),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1041),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1081),
.A2(n_1105),
.A3(n_1047),
.B(n_1106),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1045),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1009),
.A2(n_1043),
.B(n_1115),
.C(n_1015),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1077),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1060),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1044),
.A2(n_998),
.B(n_1066),
.C(n_1097),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1055),
.B(n_999),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1024),
.A2(n_1116),
.B(n_1056),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1030),
.A2(n_1040),
.B(n_1036),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1078),
.A2(n_1038),
.B(n_1112),
.C(n_1119),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1069),
.A2(n_1074),
.B(n_1103),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1093),
.A2(n_1019),
.B(n_1020),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1067),
.Y(n_1242)
);

AO21x1_ASAP7_75t_L g1243 ( 
.A1(n_1081),
.A2(n_1064),
.B(n_999),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1098),
.B(n_1026),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1046),
.B(n_1022),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1033),
.A2(n_1037),
.B(n_1010),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1026),
.A2(n_1071),
.B(n_1088),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1088),
.A2(n_944),
.B1(n_766),
.B2(n_940),
.C(n_947),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1026),
.A2(n_1088),
.B(n_1033),
.C(n_1037),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1037),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1033),
.A2(n_835),
.B1(n_986),
.B2(n_689),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1011),
.A2(n_971),
.A3(n_982),
.B(n_980),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1016),
.A2(n_1086),
.B(n_1001),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_986),
.B(n_817),
.Y(n_1254)
);

AOI221x1_ASAP7_75t_L g1255 ( 
.A1(n_982),
.A2(n_766),
.B1(n_971),
.B2(n_1101),
.C(n_988),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_986),
.B(n_817),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_986),
.B(n_817),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1007),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_980),
.A2(n_971),
.B(n_982),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_L g1260 ( 
.A(n_973),
.B(n_842),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1016),
.A2(n_1086),
.B(n_1001),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1021),
.B(n_692),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1048),
.B(n_817),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_SL g1264 ( 
.A1(n_972),
.A2(n_835),
.B(n_649),
.C(n_650),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1061),
.A2(n_766),
.B(n_688),
.C(n_835),
.Y(n_1265)
);

AND3x4_ASAP7_75t_L g1266 ( 
.A(n_976),
.B(n_821),
.C(n_1117),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1262),
.B(n_1135),
.Y(n_1267)
);

AOI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1235),
.A2(n_1265),
.B(n_1248),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1175),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1164),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1150),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1134),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1176),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1176),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1122),
.A2(n_1153),
.B(n_1242),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1255),
.A2(n_1259),
.B(n_1137),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1148),
.A2(n_1145),
.B(n_1142),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1143),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1205),
.A2(n_1204),
.B(n_1259),
.C(n_1232),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1257),
.A2(n_1163),
.B1(n_1263),
.B2(n_1266),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1135),
.B(n_1217),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1204),
.A2(n_1209),
.B(n_1210),
.C(n_1251),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1210),
.A2(n_1251),
.B(n_1248),
.C(n_1170),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1162),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1189),
.A2(n_1158),
.B(n_1190),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1215),
.A2(n_1127),
.B1(n_1133),
.B2(n_1222),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1170),
.A2(n_1213),
.B(n_1152),
.C(n_1169),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1187),
.A2(n_1123),
.B(n_1173),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1165),
.A2(n_1227),
.B(n_1194),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1215),
.A2(n_1207),
.B1(n_1206),
.B2(n_1203),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1167),
.B(n_1233),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1211),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1137),
.A2(n_1120),
.B(n_1124),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1144),
.B(n_1151),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1258),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1120),
.A2(n_1139),
.B(n_1152),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1188),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1147),
.A2(n_1239),
.B(n_1199),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1264),
.A2(n_1132),
.B(n_1131),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1222),
.A2(n_1213),
.B1(n_1218),
.B2(n_1216),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1178),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1179),
.A2(n_1226),
.B(n_1196),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1160),
.A2(n_1220),
.A3(n_1141),
.B1(n_1252),
.B2(n_1183),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1136),
.A2(n_1121),
.B(n_1166),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1163),
.B(n_1236),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1177),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1188),
.B(n_1202),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1188),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1125),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1246),
.A2(n_1240),
.B(n_1171),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1192),
.A2(n_1193),
.B(n_1237),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1149),
.B(n_1225),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1216),
.B(n_1208),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1155),
.B(n_1140),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1243),
.A2(n_1160),
.A3(n_1195),
.B(n_1192),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1185),
.A2(n_1161),
.B1(n_1176),
.B2(n_1221),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1157),
.A2(n_1140),
.B(n_1156),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1198),
.A2(n_1154),
.B(n_1180),
.C(n_1186),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1229),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1231),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1212),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1146),
.B(n_1154),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1249),
.B(n_1182),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1184),
.A2(n_1241),
.B(n_1238),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1168),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1223),
.Y(n_1328)
);

AOI21xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1219),
.A2(n_1228),
.B(n_1234),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1260),
.A2(n_1172),
.B1(n_1200),
.B2(n_1201),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1181),
.A2(n_1214),
.B(n_1168),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1245),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1141),
.A2(n_1252),
.B(n_1128),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1224),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1191),
.A2(n_1244),
.B(n_1247),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1197),
.A2(n_1141),
.B(n_1252),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1220),
.A2(n_1250),
.B1(n_1202),
.B2(n_1188),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1202),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1138),
.A2(n_1129),
.B(n_1183),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1202),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1183),
.A2(n_1129),
.B1(n_1174),
.B2(n_1159),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1129),
.A2(n_726),
.B1(n_647),
.B2(n_766),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1230),
.A2(n_1255),
.B(n_1259),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1230),
.A2(n_1261),
.B(n_1253),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1230),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1188),
.Y(n_1346)
);

OR2x6_ASAP7_75t_L g1347 ( 
.A(n_1147),
.B(n_1163),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1126),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1176),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1259),
.A2(n_766),
.B1(n_940),
.B2(n_913),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1265),
.A2(n_695),
.B(n_688),
.Y(n_1351)
);

AOI21xp33_ASAP7_75t_L g1352 ( 
.A1(n_1235),
.A2(n_688),
.B(n_695),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1259),
.A2(n_835),
.B(n_986),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1217),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1265),
.A2(n_695),
.B(n_688),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1126),
.Y(n_1358)
);

NOR2xp67_ASAP7_75t_L g1359 ( 
.A(n_1125),
.B(n_973),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1235),
.A2(n_1265),
.B(n_766),
.C(n_726),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1126),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1126),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1235),
.B(n_875),
.C(n_492),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1211),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1126),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1126),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1126),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1255),
.A2(n_1259),
.B(n_1011),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1262),
.B(n_1135),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1217),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1130),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1263),
.B(n_647),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1126),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1176),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1176),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1259),
.A2(n_766),
.B1(n_940),
.B2(n_913),
.Y(n_1381)
);

OR2x6_ASAP7_75t_L g1382 ( 
.A(n_1147),
.B(n_1163),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1126),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1211),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1259),
.A2(n_835),
.B(n_766),
.C(n_1265),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1176),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1259),
.A2(n_766),
.B1(n_940),
.B2(n_913),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1176),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1164),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1215),
.A2(n_835),
.B1(n_766),
.B2(n_1259),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1176),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1263),
.B(n_1167),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1392),
.B(n_1314),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1325),
.A2(n_1363),
.B(n_1271),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1351),
.A2(n_1356),
.B(n_1300),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1267),
.B(n_1374),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1385),
.A2(n_1360),
.B(n_1364),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1350),
.A2(n_1381),
.B1(n_1387),
.B2(n_1292),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1315),
.B(n_1293),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1283),
.B(n_1355),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1296),
.B(n_1307),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1350),
.A2(n_1387),
.B1(n_1381),
.B2(n_1292),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1296),
.B(n_1307),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1377),
.A2(n_1302),
.B1(n_1288),
.B2(n_1330),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1281),
.A2(n_1385),
.B(n_1352),
.C(n_1354),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1277),
.A2(n_1301),
.B(n_1291),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1276),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1377),
.B(n_1324),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1324),
.B(n_1316),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1318),
.B(n_1282),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1355),
.B(n_1375),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1375),
.B(n_1269),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1289),
.A2(n_1347),
.B(n_1382),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1316),
.B(n_1272),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1337),
.A2(n_1284),
.B(n_1390),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1289),
.A2(n_1390),
.B(n_1285),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1328),
.B(n_1308),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1277),
.A2(n_1326),
.B(n_1285),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1332),
.A2(n_1382),
.B1(n_1347),
.B2(n_1334),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1280),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1323),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1313),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1313),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1268),
.A2(n_1342),
.B(n_1337),
.C(n_1320),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1286),
.B(n_1297),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1348),
.B(n_1358),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1320),
.A2(n_1347),
.B(n_1382),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1276),
.Y(n_1428)
);

O2A1O1Ixp5_ASAP7_75t_L g1429 ( 
.A1(n_1341),
.A2(n_1319),
.B(n_1303),
.C(n_1336),
.Y(n_1429)
);

O2A1O1Ixp5_ASAP7_75t_L g1430 ( 
.A1(n_1303),
.A2(n_1389),
.B(n_1383),
.C(n_1368),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1287),
.A2(n_1279),
.B(n_1304),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1294),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1274),
.B(n_1389),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1334),
.A2(n_1273),
.B1(n_1345),
.B2(n_1391),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1279),
.A2(n_1344),
.B(n_1357),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1361),
.A2(n_1378),
.B(n_1367),
.C(n_1370),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1353),
.A2(n_1357),
.B(n_1373),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1379),
.A2(n_1391),
.B1(n_1380),
.B2(n_1275),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1362),
.A2(n_1329),
.B(n_1322),
.C(n_1321),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1340),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1331),
.A2(n_1340),
.B(n_1335),
.C(n_1278),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1313),
.B(n_1343),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1343),
.B(n_1317),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1349),
.B(n_1388),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1353),
.A2(n_1373),
.B(n_1366),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1294),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1349),
.B(n_1388),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1386),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1327),
.B(n_1278),
.Y(n_1449)
);

CKINVDCx14_ASAP7_75t_R g1450 ( 
.A(n_1384),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1386),
.B(n_1359),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1311),
.B(n_1380),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1343),
.B(n_1298),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1339),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1372),
.A2(n_1298),
.B(n_1295),
.C(n_1309),
.Y(n_1455)
);

NOR2xp67_ASAP7_75t_L g1456 ( 
.A(n_1311),
.B(n_1365),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_L g1457 ( 
.A(n_1365),
.B(n_1340),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1335),
.B(n_1305),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1338),
.A2(n_1340),
.B1(n_1384),
.B2(n_1309),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1317),
.B(n_1295),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1366),
.A2(n_1290),
.B(n_1270),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1305),
.B(n_1338),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1317),
.B(n_1339),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1305),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1305),
.B(n_1299),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1339),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1299),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1295),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1310),
.A2(n_1346),
.B1(n_1306),
.B2(n_1333),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1312),
.A2(n_1346),
.B(n_1310),
.C(n_1376),
.Y(n_1471)
);

NOR2xp67_ASAP7_75t_L g1472 ( 
.A(n_1310),
.B(n_1346),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1369),
.A2(n_1259),
.B(n_835),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_SL g1474 ( 
.A1(n_1371),
.A2(n_835),
.B(n_1265),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1350),
.A2(n_1387),
.B1(n_1381),
.B2(n_1292),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1267),
.B(n_1374),
.Y(n_1476)
);

INVxp33_ASAP7_75t_L g1477 ( 
.A(n_1293),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1296),
.B(n_1271),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1276),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1267),
.B(n_1374),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1392),
.B(n_1314),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1351),
.A2(n_1259),
.B(n_835),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1351),
.A2(n_1259),
.B(n_835),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1392),
.B(n_1314),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1409),
.B(n_1478),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1465),
.B(n_1458),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1413),
.B(n_1427),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1395),
.B(n_1474),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1414),
.B(n_1400),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1454),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1482),
.B(n_1483),
.Y(n_1491)
);

AOI211xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1397),
.A2(n_1398),
.B(n_1402),
.C(n_1475),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1404),
.A2(n_1416),
.B1(n_1410),
.B2(n_1408),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1473),
.B(n_1424),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1411),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1412),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1462),
.B(n_1401),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1403),
.B(n_1464),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1466),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1420),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1443),
.B(n_1442),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1449),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1441),
.A2(n_1469),
.B(n_1405),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1484),
.B(n_1393),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1430),
.Y(n_1505)
);

AOI21xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1419),
.A2(n_1459),
.B(n_1451),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1430),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1481),
.B(n_1477),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1422),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1396),
.B(n_1476),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1460),
.B(n_1453),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1480),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1422),
.Y(n_1514)
);

AO21x2_ASAP7_75t_L g1515 ( 
.A1(n_1441),
.A2(n_1405),
.B(n_1455),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_1429),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1423),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1470),
.A2(n_1423),
.B(n_1437),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1425),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1436),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1426),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1463),
.B(n_1418),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1417),
.B(n_1433),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1471),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1431),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1452),
.B(n_1457),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1418),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1435),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1407),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1435),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1516),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1486),
.B(n_1406),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1434),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1499),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1509),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1493),
.A2(n_1399),
.B1(n_1450),
.B2(n_1415),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1509),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1502),
.B(n_1439),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1501),
.B(n_1461),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1501),
.B(n_1461),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1490),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1516),
.Y(n_1543)
);

NAND5xp2_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1491),
.C(n_1520),
.D(n_1485),
.E(n_1415),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1487),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1502),
.B(n_1421),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1524),
.Y(n_1547)
);

OAI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1492),
.A2(n_1456),
.B1(n_1438),
.B2(n_1468),
.C(n_1472),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1512),
.B(n_1437),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1503),
.B(n_1437),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1503),
.B(n_1445),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1525),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1467),
.Y(n_1553)
);

AOI21xp33_ASAP7_75t_L g1554 ( 
.A1(n_1491),
.A2(n_1394),
.B(n_1450),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1428),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1547),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1534),
.B(n_1494),
.C(n_1520),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1533),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1531),
.B(n_1498),
.Y(n_1559)
);

NAND4xp25_ASAP7_75t_SL g1560 ( 
.A(n_1537),
.B(n_1506),
.C(n_1432),
.D(n_1446),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1550),
.A2(n_1530),
.B(n_1527),
.Y(n_1561)
);

NOR4xp25_ASAP7_75t_SL g1562 ( 
.A(n_1554),
.B(n_1524),
.C(n_1526),
.D(n_1505),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1539),
.A2(n_1518),
.B(n_1505),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1546),
.B(n_1495),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1533),
.Y(n_1565)
);

NAND4xp25_ASAP7_75t_L g1566 ( 
.A(n_1544),
.B(n_1495),
.C(n_1510),
.D(n_1489),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1546),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1544),
.B(n_1513),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1555),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_SL g1570 ( 
.A(n_1550),
.B(n_1507),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1534),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1537),
.A2(n_1487),
.B1(n_1548),
.B2(n_1488),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1531),
.B(n_1496),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1498),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1535),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1548),
.A2(n_1487),
.B1(n_1488),
.B2(n_1494),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1554),
.A2(n_1539),
.B(n_1488),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1555),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1542),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1497),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1555),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1552),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1542),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1547),
.A2(n_1488),
.B1(n_1494),
.B2(n_1487),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1545),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1514),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1547),
.A2(n_1507),
.B(n_1508),
.C(n_1487),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1536),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1547),
.A2(n_1521),
.B1(n_1519),
.B2(n_1508),
.C(n_1500),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1553),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1532),
.B(n_1497),
.Y(n_1594)
);

INVxp67_ASAP7_75t_SL g1595 ( 
.A(n_1538),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1536),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1538),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1594),
.B(n_1559),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1589),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1594),
.B(n_1532),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1556),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1504),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1556),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1565),
.Y(n_1606)
);

INVx4_ASAP7_75t_SL g1607 ( 
.A(n_1565),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1587),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1561),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

INVx4_ASAP7_75t_L g1612 ( 
.A(n_1587),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1576),
.Y(n_1614)
);

INVx4_ASAP7_75t_SL g1615 ( 
.A(n_1597),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1580),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1580),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1557),
.A2(n_1488),
.B(n_1494),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1585),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1585),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1569),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1561),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1559),
.B(n_1532),
.Y(n_1623)
);

NOR2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1557),
.B(n_1545),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1563),
.A2(n_1551),
.B(n_1550),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_SL g1626 ( 
.A(n_1571),
.B(n_1523),
.C(n_1521),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1579),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1561),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1563),
.A2(n_1518),
.B(n_1528),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1583),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1590),
.A2(n_1551),
.B(n_1578),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1587),
.B(n_1545),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1573),
.B(n_1540),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1573),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1582),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1582),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1633),
.B(n_1570),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1584),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1615),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1634),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1593),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1626),
.B(n_1568),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1624),
.B(n_1581),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1630),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1603),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1615),
.B(n_1584),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1624),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1603),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1608),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1606),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1564),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1627),
.B(n_1553),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1618),
.A2(n_1560),
.B(n_1577),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1606),
.Y(n_1658)
);

AND2x2_ASAP7_75t_SL g1659 ( 
.A(n_1631),
.B(n_1545),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1604),
.B(n_1592),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1602),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1633),
.B(n_1570),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1608),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1635),
.B(n_1553),
.Y(n_1664)
);

OAI33xp33_ASAP7_75t_L g1665 ( 
.A1(n_1609),
.A2(n_1566),
.A3(n_1572),
.B1(n_1541),
.B2(n_1540),
.B3(n_1588),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1636),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1623),
.B(n_1581),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1609),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1623),
.B(n_1584),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1611),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1610),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1636),
.B(n_1567),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1615),
.B(n_1562),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1611),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_R g1675 ( 
.A(n_1612),
.B(n_1407),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_L g1677 ( 
.A(n_1612),
.B(n_1597),
.Y(n_1677)
);

NAND2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1602),
.B(n_1545),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1601),
.B(n_1596),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1614),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1655),
.B(n_1648),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1675),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1643),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1661),
.B(n_1614),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1663),
.B(n_1612),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1639),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1646),
.B(n_1618),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1632),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1645),
.B(n_1664),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1656),
.B(n_1605),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1642),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1649),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1652),
.Y(n_1693)
);

OAI222xp33_ASAP7_75t_L g1694 ( 
.A1(n_1660),
.A2(n_1494),
.B1(n_1586),
.B2(n_1605),
.C1(n_1612),
.C2(n_1632),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1651),
.A2(n_1601),
.B(n_1600),
.Y(n_1695)
);

OR2x2_ASAP7_75t_SL g1696 ( 
.A(n_1672),
.B(n_1631),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1654),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1658),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1632),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1668),
.Y(n_1700)
);

NAND2x1_ASAP7_75t_L g1701 ( 
.A(n_1677),
.B(n_1600),
.Y(n_1701)
);

NOR2x1p5_ASAP7_75t_SL g1702 ( 
.A(n_1637),
.B(n_1662),
.Y(n_1702)
);

NAND2xp67_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1610),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1670),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1657),
.B(n_1631),
.C(n_1625),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1665),
.B(n_1504),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1657),
.A2(n_1631),
.B(n_1625),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1675),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1640),
.B(n_1570),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1638),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1659),
.B(n_1625),
.C(n_1632),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1653),
.B(n_1616),
.Y(n_1712)
);

NOR2xp67_ASAP7_75t_L g1713 ( 
.A(n_1643),
.B(n_1600),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1659),
.A2(n_1673),
.B1(n_1515),
.B2(n_1640),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1641),
.B(n_1667),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1710),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1705),
.A2(n_1515),
.B1(n_1625),
.B2(n_1678),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1638),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1686),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1687),
.A2(n_1515),
.B1(n_1678),
.B2(n_1666),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1708),
.B(n_1706),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1706),
.B(n_1641),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1681),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.B(n_1666),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1715),
.B(n_1676),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1689),
.B(n_1674),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1684),
.B(n_1712),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1638),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1685),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1692),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1685),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1693),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1683),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1687),
.A2(n_1515),
.B1(n_1676),
.B2(n_1667),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1710),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1697),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1703),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1695),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1698),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1684),
.B(n_1637),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1722),
.A2(n_1707),
.B1(n_1699),
.B2(n_1688),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1739),
.B(n_1707),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1714),
.B1(n_1711),
.B2(n_1701),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1717),
.A2(n_1694),
.B1(n_1680),
.B2(n_1704),
.C(n_1700),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1716),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1725),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1725),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1726),
.B(n_1679),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1730),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1733),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1729),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1733),
.Y(n_1753)
);

OAI222xp33_ASAP7_75t_L g1754 ( 
.A1(n_1735),
.A2(n_1709),
.B1(n_1696),
.B2(n_1662),
.C1(n_1694),
.C2(n_1680),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1738),
.A2(n_1724),
.B(n_1732),
.C(n_1723),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1737),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1737),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1729),
.B(n_1650),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_1702),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1727),
.Y(n_1760)
);

INVxp67_ASAP7_75t_L g1761 ( 
.A(n_1718),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1728),
.B(n_1727),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1752),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1750),
.B(n_1734),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1752),
.B(n_1718),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1747),
.B(n_1728),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1761),
.B(n_1734),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1736),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1758),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1755),
.B(n_1718),
.Y(n_1770)
);

NAND3xp33_ASAP7_75t_L g1771 ( 
.A(n_1743),
.B(n_1745),
.C(n_1744),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1741),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1736),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1771),
.B(n_1743),
.C(n_1759),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1770),
.B(n_1759),
.C(n_1742),
.Y(n_1775)
);

AND4x1_ASAP7_75t_L g1776 ( 
.A(n_1764),
.B(n_1758),
.C(n_1721),
.D(n_1757),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1772),
.A2(n_1754),
.B(n_1765),
.C(n_1767),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1766),
.A2(n_1749),
.B(n_1746),
.Y(n_1778)
);

AOI21xp33_ASAP7_75t_SL g1779 ( 
.A1(n_1763),
.A2(n_1759),
.B(n_1746),
.Y(n_1779)
);

NOR3xp33_ASAP7_75t_L g1780 ( 
.A(n_1768),
.B(n_1756),
.C(n_1753),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1769),
.B(n_1719),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1773),
.B(n_1751),
.Y(n_1782)
);

AOI321xp33_ASAP7_75t_L g1783 ( 
.A1(n_1777),
.A2(n_1720),
.A3(n_1740),
.B1(n_1731),
.B2(n_1741),
.C(n_1729),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1781),
.Y(n_1784)
);

OR3x2_ASAP7_75t_L g1785 ( 
.A(n_1776),
.B(n_1617),
.C(n_1616),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1774),
.A2(n_1712),
.B1(n_1671),
.B2(n_1628),
.C(n_1622),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1782),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1787),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1784),
.B(n_1778),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1783),
.B(n_1775),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1785),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1786),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1787),
.B(n_1779),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1790),
.A2(n_1622),
.B1(n_1610),
.B2(n_1628),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1789),
.B(n_1780),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_L g1796 ( 
.A(n_1793),
.B(n_1671),
.C(n_1628),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1793),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1792),
.A2(n_1622),
.B1(n_1650),
.B2(n_1669),
.C(n_1679),
.Y(n_1798)
);

NOR3xp33_ASAP7_75t_L g1799 ( 
.A(n_1795),
.B(n_1788),
.C(n_1791),
.Y(n_1799)
);

AND2x2_ASAP7_75t_SL g1800 ( 
.A(n_1796),
.B(n_1798),
.Y(n_1800)
);

NOR3xp33_ASAP7_75t_L g1801 ( 
.A(n_1797),
.B(n_1650),
.C(n_1511),
.Y(n_1801)
);

AND3x2_ASAP7_75t_L g1802 ( 
.A(n_1799),
.B(n_1794),
.C(n_1669),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1802),
.B(n_1800),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1803),
.Y(n_1804)
);

INVxp33_ASAP7_75t_SL g1805 ( 
.A(n_1803),
.Y(n_1805)
);

NOR3xp33_ASAP7_75t_SL g1806 ( 
.A(n_1805),
.B(n_1801),
.C(n_1613),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1804),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1806),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1613),
.B(n_1629),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1808),
.A2(n_1600),
.B1(n_1620),
.B2(n_1619),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1809),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1811),
.A2(n_1620),
.B(n_1619),
.Y(n_1812)
);

OAI21x1_ASAP7_75t_SL g1813 ( 
.A1(n_1812),
.A2(n_1810),
.B(n_1529),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1813),
.A2(n_1479),
.B1(n_1448),
.B2(n_1617),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1607),
.B1(n_1595),
.B2(n_1479),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1448),
.B(n_1444),
.C(n_1447),
.Y(n_1816)
);


endmodule