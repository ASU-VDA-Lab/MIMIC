module fake_jpeg_20758_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

OAI211xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_16),
.B(n_26),
.C(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_38),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_54),
.B1(n_33),
.B2(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_40),
.B1(n_33),
.B2(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_60),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_15),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_27),
.B1(n_31),
.B2(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_71),
.B1(n_17),
.B2(n_21),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_27),
.B1(n_18),
.B2(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_73),
.B1(n_23),
.B2(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_40),
.B1(n_33),
.B2(n_26),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_32),
.B(n_35),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_44),
.B(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_23),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_49),
.B(n_54),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_80),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_84),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_49),
.B(n_46),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_44),
.C(n_20),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_20),
.C(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_96),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_69),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_16),
.C(n_10),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_92),
.C(n_94),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_19),
.B(n_22),
.C(n_23),
.D(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_94),
.B1(n_63),
.B2(n_57),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_14),
.A3(n_12),
.B1(n_8),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_14),
.C(n_1),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_63),
.B1(n_66),
.B2(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_83),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_3),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_84),
.C(n_85),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_120),
.C(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_96),
.C(n_92),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_96),
.B(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_98),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_57),
.B(n_75),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_126),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_97),
.Y(n_132)
);

AOI21x1_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_22),
.B(n_6),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_105),
.C(n_99),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_122),
.B(n_118),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_150),
.B(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_118),
.B1(n_125),
.B2(n_119),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_124),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_119),
.B(n_129),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_131),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_154),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_124),
.B(n_146),
.C(n_127),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_102),
.B(n_125),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_135),
.B(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_163),
.B(n_164),
.C(n_159),
.D(n_126),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_144),
.Y(n_161)
);

AOI31xp33_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_121),
.A3(n_120),
.B(n_111),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_145),
.B1(n_147),
.B2(n_150),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_166),
.B1(n_160),
.B2(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_138),
.C(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_107),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_168),
.B(n_7),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_107),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_169),
.C(n_7),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);


endmodule