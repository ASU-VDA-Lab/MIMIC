module fake_jpeg_25798_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_53),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_17),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_55),
.C(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_40),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_21),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_41),
.B1(n_24),
.B2(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_18),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_77),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_25),
.B(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_28),
.B1(n_23),
.B2(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_23),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_19),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_29),
.C(n_28),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_49),
.B1(n_58),
.B2(n_54),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_82),
.B1(n_87),
.B2(n_29),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_49),
.B1(n_45),
.B2(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_33),
.C(n_32),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_93),
.C(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_70),
.B1(n_62),
.B2(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_54),
.B1(n_35),
.B2(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_38),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_33),
.C(n_32),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_95),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_77),
.B(n_68),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_101),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_106),
.B1(n_81),
.B2(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_90),
.B1(n_84),
.B2(n_88),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_68),
.B(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_110),
.B(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_84),
.C(n_91),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_37),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_100),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_136),
.C(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_127),
.B1(n_0),
.B2(n_1),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_88),
.B(n_31),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_124),
.CI(n_123),
.CON(n_133),
.SN(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_135),
.A2(n_119),
.B(n_31),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_139),
.C(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_117),
.C(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_127),
.B(n_126),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_15),
.B1(n_95),
.B2(n_7),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_15),
.B1(n_5),
.B2(n_9),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_145),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_137),
.B(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_151),
.Y(n_154)
);

AO221x1_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_148),
.B(n_138),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_156),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_4),
.B(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_160),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_149),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_158),
.B(n_11),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_13),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_13),
.B(n_163),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_1),
.B(n_2),
.Y(n_167)
);

XNOR2x2_ASAP7_75t_SL g168 ( 
.A(n_167),
.B(n_165),
.Y(n_168)
);


endmodule