module fake_jpeg_2274_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_60),
.Y(n_68)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_55),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_50),
.B1(n_56),
.B2(n_53),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_86),
.B1(n_67),
.B2(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_64),
.B1(n_65),
.B2(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_67),
.B1(n_59),
.B2(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_61),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_81),
.C(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_97),
.C(n_52),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_51),
.B1(n_50),
.B2(n_56),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_103),
.B1(n_60),
.B2(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_57),
.B(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_5),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_82),
.B1(n_55),
.B2(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_82),
.B1(n_60),
.B2(n_54),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_58),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_47),
.C(n_46),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_45),
.C(n_44),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_33),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_5),
.C(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_6),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_36),
.B(n_34),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_38),
.B(n_37),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_141),
.B(n_29),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_126),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_138),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_114),
.B(n_118),
.C(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_7),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_7),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_32),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_144),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_8),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_142),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_31),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_159),
.B1(n_127),
.B2(n_143),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_12),
.B(n_13),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_148),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_24),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_23),
.C(n_16),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_160),
.C(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_17),
.C(n_18),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_143),
.B1(n_130),
.B2(n_124),
.C(n_137),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_169),
.B1(n_168),
.B2(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_152),
.B(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_168),
.B1(n_130),
.B2(n_162),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_172),
.B(n_150),
.Y(n_181)
);

OAI221xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_177),
.B1(n_158),
.B2(n_174),
.C(n_179),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_180),
.B(n_146),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_155),
.B(n_140),
.Y(n_184)
);

NOR2x1p5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_150),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_166),
.C(n_160),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_134),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_18),
.Y(n_188)
);


endmodule