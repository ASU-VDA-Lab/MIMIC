module fake_netlist_1_8328_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2x1p5_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
OAI21xp5_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
NAND3xp33_ASAP7_75t_L g8 ( .A(n_6), .B(n_4), .C(n_1), .Y(n_8) );
NOR2x1_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .Y(n_9) );
AOI211xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_7), .B(n_8), .C(n_2), .Y(n_10) );
O2A1O1Ixp33_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_0), .B(n_1), .C(n_2), .Y(n_11) );
AOI22xp33_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_11), .B(n_0), .Y(n_13) );
endmodule