module fake_jpeg_10964_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx24_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_0),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_22),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_20),
.A2(n_26),
.B(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_14),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_9),
.B1(n_12),
.B2(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_3),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_13),
.B1(n_11),
.B2(n_8),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_17),
.B(n_8),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_20),
.B(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_32),
.C(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_33),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_34),
.B(n_38),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_39),
.B1(n_36),
.B2(n_21),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_37),
.C(n_34),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_47),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_45),
.B1(n_42),
.B2(n_12),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_37),
.Y(n_49)
);

XNOR2x1_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_28),
.B(n_50),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_49),
.B(n_17),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_51),
.B(n_5),
.C(n_9),
.Y(n_57)
);


endmodule