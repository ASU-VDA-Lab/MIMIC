module fake_jpeg_19008_n_252 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_46),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_19),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_56),
.B1(n_62),
.B2(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_30),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_45),
.C(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_34),
.B1(n_18),
.B2(n_23),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_30),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_24),
.B1(n_27),
.B2(n_35),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_35),
.B1(n_27),
.B2(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_35),
.B1(n_27),
.B2(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_25),
.B1(n_17),
.B2(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_71),
.B1(n_73),
.B2(n_20),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_25),
.B1(n_17),
.B2(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_21),
.B1(n_19),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_80),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_40),
.Y(n_80)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_45),
.C(n_44),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_29),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_92),
.Y(n_126)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_45),
.B(n_41),
.C(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_105),
.Y(n_119)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_60),
.B(n_54),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_106),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_59),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_74),
.B1(n_75),
.B2(n_20),
.Y(n_133)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_63),
.B(n_68),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_115),
.B(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_15),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_66),
.B1(n_74),
.B2(n_58),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_133),
.B1(n_90),
.B2(n_101),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_80),
.B(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_66),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_59),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_87),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_138),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_83),
.B1(n_87),
.B2(n_84),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_137),
.B1(n_117),
.B2(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_131),
.B1(n_110),
.B2(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_94),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_83),
.B1(n_104),
.B2(n_100),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_159),
.B1(n_29),
.B2(n_31),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_149),
.B1(n_120),
.B2(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_158),
.B(n_26),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_113),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_101),
.B1(n_88),
.B2(n_96),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_134),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_119),
.B(n_117),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_143),
.B(n_135),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_92),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_124),
.B(n_118),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_160),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_168),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_144),
.B1(n_136),
.B2(n_141),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_26),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_82),
.B1(n_112),
.B2(n_109),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_105),
.C(n_106),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_156),
.C(n_155),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_122),
.B1(n_26),
.B2(n_3),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_178),
.B1(n_160),
.B2(n_3),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_26),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_177),
.B1(n_180),
.B2(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_158),
.B1(n_146),
.B2(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_194),
.B1(n_173),
.B2(n_164),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_140),
.B(n_138),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_15),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_7),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.C(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_159),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_163),
.B1(n_169),
.B2(n_162),
.Y(n_194)
);

OAI322xp33_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_154),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_162),
.B1(n_161),
.B2(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_5),
.C(n_6),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_204),
.B1(n_206),
.B2(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_191),
.C(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_183),
.C(n_179),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_179),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

NAND4xp25_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_220),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_200),
.B1(n_184),
.B2(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_226),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_185),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_212),
.B(n_204),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_196),
.B(n_188),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_203),
.B1(n_211),
.B2(n_216),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_203),
.C(n_208),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_161),
.C(n_11),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_224),
.C(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_207),
.C(n_206),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_170),
.B(n_174),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_170),
.B1(n_174),
.B2(n_161),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_10),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_244),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_231),
.B1(n_228),
.B2(n_12),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_238),
.C(n_243),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_246),
.C(n_10),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_228),
.C(n_235),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_242),
.C(n_11),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_248),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_249),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_12),
.Y(n_252)
);


endmodule