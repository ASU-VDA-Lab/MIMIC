module fake_jpeg_25264_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_19),
.C(n_31),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_39),
.C(n_44),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_17),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_61),
.B(n_68),
.C(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_19),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_22),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_24),
.B1(n_20),
.B2(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_62),
.B1(n_36),
.B2(n_26),
.Y(n_91)
);

AOI32xp33_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_18),
.A3(n_30),
.B1(n_27),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_24),
.B1(n_30),
.B2(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_17),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_31),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_85),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_70),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_23),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_79),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_36),
.B1(n_26),
.B2(n_44),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_92),
.B1(n_98),
.B2(n_47),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_52),
.B(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_84),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_90),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_99),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_58),
.B(n_14),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_36),
.B1(n_44),
.B2(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_17),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_97),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_31),
.B1(n_34),
.B2(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_39),
.C(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_16),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_39),
.B1(n_37),
.B2(n_34),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_43),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_43),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_43),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_88),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_112),
.B(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_47),
.B1(n_49),
.B2(n_2),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_123),
.B1(n_100),
.B2(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_43),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_0),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_127),
.B(n_105),
.C(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_110),
.B(n_117),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_86),
.B1(n_87),
.B2(n_85),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_136),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_138)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_70),
.B1(n_72),
.B2(n_98),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_70),
.C(n_96),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_144),
.C(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_101),
.B1(n_79),
.B2(n_80),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_148),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_74),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_82),
.C(n_15),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_167),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

AOI21x1_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_144),
.B(n_131),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_174),
.B(n_175),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_2),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_116),
.A3(n_112),
.B1(n_119),
.B2(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_173),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_111),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_129),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_103),
.B(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_137),
.B1(n_141),
.B2(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_184),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_170),
.CI(n_163),
.CON(n_179),
.SN(n_179)
);

OAI322xp33_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_158),
.A3(n_165),
.B1(n_166),
.B2(n_174),
.C1(n_156),
.C2(n_168),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_104),
.B(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_3),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_138),
.B1(n_114),
.B2(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_155),
.B1(n_169),
.B2(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_149),
.B1(n_130),
.B2(n_134),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_161),
.B(n_173),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_153),
.C(n_15),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_191),
.C(n_158),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_160),
.C(n_167),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_1),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_194),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_202),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_198),
.A2(n_204),
.B1(n_209),
.B2(n_194),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_193),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_207),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_206),
.B(n_178),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_159),
.C(n_161),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_205),
.C(n_184),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_179),
.C(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_179),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_213),
.B(n_215),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_187),
.C(n_188),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_219),
.C(n_220),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_208),
.A2(n_190),
.B(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND4xp25_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_200),
.C(n_195),
.D(n_207),
.Y(n_229)
);

OAI321xp33_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_192),
.A3(n_203),
.B1(n_211),
.B2(n_219),
.C(n_12),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_8),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_210),
.C(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_227),
.C(n_9),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_214),
.B(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_226),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_8),
.B(n_9),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_239),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_234),
.B1(n_10),
.B2(n_12),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_238),
.C(n_9),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_240),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_246),
.B1(n_242),
.B2(n_10),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_10),
.Y(n_248)
);


endmodule