module fake_jpeg_27258_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_70),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_0),
.Y(n_81)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_52),
.B(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_83),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_57),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_53),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_61),
.B1(n_62),
.B2(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_94),
.B1(n_46),
.B2(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_2),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_61),
.B1(n_51),
.B2(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_100),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_60),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_102),
.B(n_107),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_48),
.B(n_16),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_50),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_77),
.B1(n_63),
.B2(n_20),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_91),
.B1(n_96),
.B2(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_19),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_14),
.B(n_34),
.Y(n_125)
);

INVxp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_119),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_124),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_111),
.B1(n_90),
.B2(n_4),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_18),
.B(n_36),
.C(n_35),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_129),
.C(n_8),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_13),
.C(n_31),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.C(n_6),
.Y(n_132)
);

XOR2x2_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_131),
.B(n_130),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_126),
.B(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_127),
.B(n_123),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_3),
.Y(n_140)
);

INVxp33_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_22),
.B(n_29),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_7),
.Y(n_143)
);


endmodule