module real_jpeg_10595_n_12 (n_290, n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_289, n_3, n_10, n_9, n_12);

input n_290;
input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_289;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_181;
wire n_102;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_8),
.B(n_27),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_4),
.A2(n_40),
.B(n_63),
.C(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_40),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_8),
.B(n_65),
.Y(n_99)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_8),
.A2(n_18),
.B1(n_19),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_8),
.A2(n_51),
.B1(n_64),
.B2(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_8),
.B(n_37),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_8),
.A2(n_26),
.B(n_39),
.C(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_28),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_9),
.A2(n_20),
.B1(n_64),
.B2(n_65),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_9),
.A2(n_20),
.B1(n_40),
.B2(n_42),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_11),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_30),
.B1(n_40),
.B2(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_30),
.B1(n_64),
.B2(n_65),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_282),
.B(n_285),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_72),
.B(n_281),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_15),
.B(n_31),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_15),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_17),
.A2(n_25),
.B(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_19),
.A2(n_23),
.B(n_51),
.C(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_22),
.A2(n_25),
.B1(n_50),
.B2(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_22),
.B(n_25),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_38),
.B(n_39),
.C(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_28),
.A2(n_49),
.B(n_58),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_29),
.B(n_239),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_32),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_32),
.B(n_279),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_47),
.CI(n_52),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_37),
.B1(n_44),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_36),
.B(n_130),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_37),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_37),
.A2(n_44),
.B1(n_128),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_38),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_40),
.A2(n_43),
.B(n_51),
.Y(n_134)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_42),
.A2(n_51),
.B(n_68),
.C(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_45),
.B(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_50),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_51),
.B(n_63),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.C(n_60),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_53),
.A2(n_60),
.B1(n_259),
.B2(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_54),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_55),
.A2(n_56),
.B1(n_144),
.B2(n_150),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_55),
.B(n_144),
.C(n_187),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_55),
.A2(n_56),
.B1(n_127),
.B2(n_131),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_55),
.B(n_127),
.C(n_216),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_55),
.A2(n_56),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_60),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_62),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_63),
.A2(n_69),
.B1(n_93),
.B2(n_96),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_63),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_222),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_64),
.B(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_278),
.B(n_280),
.Y(n_72)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_251),
.A3(n_271),
.B1(n_276),
.B2(n_277),
.C(n_289),
.Y(n_73)
);

AOI321xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_206),
.A3(n_226),
.B1(n_245),
.B2(n_250),
.C(n_290),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_175),
.C(n_203),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_155),
.B(n_174),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_140),
.B(n_154),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_122),
.B(n_139),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_111),
.B(n_121),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_101),
.B(n_110),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_90),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_82),
.A2(n_103),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_144),
.C(n_149),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_86),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_85),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_85),
.A2(n_137),
.B1(n_182),
.B2(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_87),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_88),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_98),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_100),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_127),
.C(n_138),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_91),
.A2(n_100),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_100),
.B(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B(n_109),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_107),
.B(n_108),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_114),
.B1(n_115),
.B2(n_120),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_116),
.C(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_108),
.A2(n_120),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_108),
.B(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_119),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_119),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_194),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_143),
.C(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_132),
.B2(n_138),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_131),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_161),
.C(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_129),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_136),
.B(n_196),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_142),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_151),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_150),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_150),
.B(n_232),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_167),
.C(n_173),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_164),
.A2(n_165),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_164),
.A2(n_165),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_164),
.A2(n_165),
.B1(n_265),
.B2(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_164),
.B(n_259),
.C(n_260),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_164),
.B(n_269),
.C(n_270),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_165),
.B(n_198),
.C(n_200),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_176),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_188),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_177),
.B(n_188),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_184),
.CI(n_185),
.CON(n_177),
.SN(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_202),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_197),
.C(n_202),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_207),
.A2(n_246),
.B(n_249),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_208),
.B(n_209),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_225),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_217),
.B2(n_218),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_218),
.C(n_225),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_220),
.B1(n_237),
.B2(n_240),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_221),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_235),
.B(n_237),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_228),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_243),
.B2(n_244),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_231),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_242),
.C(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_253),
.C(n_261),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_253),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_263),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_263),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_262),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);


endmodule