module fake_aes_3479_n_542 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_542);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_542;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g69 ( .A(n_2), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_49), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_43), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_2), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_46), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_15), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_22), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_41), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_35), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_17), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_42), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_45), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_14), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_24), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_3), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_55), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_21), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_33), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_63), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_18), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_40), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_5), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_53), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_65), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_50), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_30), .Y(n_100) );
OR2x2_ASAP7_75t_L g101 ( .A(n_19), .B(n_16), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_29), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_16), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_70), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_105), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_84), .B(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_105), .Y(n_110) );
XOR2xp5_ASAP7_75t_L g111 ( .A(n_82), .B(n_77), .Y(n_111) );
AND2x6_ASAP7_75t_L g112 ( .A(n_99), .B(n_28), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_83), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_85), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_96), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_100), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_99), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_96), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_76), .B(n_0), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_76), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_69), .B(n_1), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_90), .B(n_31), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_69), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_117), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_122), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_130), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_106), .B(n_91), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_112), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_134), .A2(n_104), .B1(n_78), .B2(n_88), .Y(n_146) );
INVx5_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_130), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
AO22x2_ASAP7_75t_L g150 ( .A1(n_111), .A2(n_101), .B1(n_103), .B2(n_90), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_131), .Y(n_151) );
AO22x2_ASAP7_75t_L g152 ( .A1(n_111), .A2(n_101), .B1(n_103), .B2(n_91), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_106), .B(n_89), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_109), .B(n_113), .Y(n_156) );
CKINVDCx6p67_ASAP7_75t_R g157 ( .A(n_133), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_109), .B(n_94), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_113), .B(n_87), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_114), .B(n_97), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_114), .B(n_74), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_115), .A2(n_104), .B1(n_72), .B2(n_78), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_115), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
NAND3xp33_ASAP7_75t_L g166 ( .A(n_118), .B(n_93), .C(n_94), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_163), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_149), .B(n_126), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_137), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_149), .B(n_128), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_143), .B(n_118), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_143), .A2(n_132), .B1(n_121), .B2(n_119), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_140), .A2(n_122), .B1(n_128), .B2(n_132), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_140), .B(n_119), .Y(n_177) );
INVxp33_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
OR2x2_ASAP7_75t_L g180 ( .A(n_154), .B(n_116), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_154), .B(n_116), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_156), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_155), .B(n_121), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_156), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_136), .Y(n_187) );
NOR2xp33_ASAP7_75t_SL g188 ( .A(n_149), .B(n_133), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_149), .B(n_102), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_156), .A2(n_133), .B1(n_110), .B2(n_123), .Y(n_194) );
INVxp67_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_147), .B(n_98), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_150), .A2(n_133), .B1(n_127), .B2(n_129), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_161), .B(n_123), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_162), .B(n_124), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_141), .B(n_110), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_162), .B(n_124), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_142), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_160), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_188), .A2(n_147), .B(n_142), .Y(n_207) );
INVx8_ASAP7_75t_L g208 ( .A(n_199), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_191), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_191), .B(n_142), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_199), .A2(n_152), .B1(n_150), .B2(n_160), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_205), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_202), .Y(n_213) );
INVx8_ASAP7_75t_L g214 ( .A(n_199), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_187), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_204), .A2(n_152), .B1(n_150), .B2(n_160), .Y(n_216) );
INVx3_ASAP7_75t_SL g217 ( .A(n_169), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_202), .B(n_150), .Y(n_218) );
BUFx2_ASAP7_75t_SL g219 ( .A(n_183), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_195), .B(n_152), .Y(n_220) );
NAND2x2_ASAP7_75t_L g221 ( .A(n_180), .B(n_152), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_205), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_171), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_167), .B(n_158), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_167), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_172), .B(n_146), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_172), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_198), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_201), .Y(n_229) );
AOI21x1_ASAP7_75t_L g230 ( .A1(n_170), .A2(n_158), .B(n_165), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_204), .B(n_159), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_178), .B(n_124), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_204), .B(n_152), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_180), .B(n_124), .Y(n_234) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_183), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_185), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_182), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_173), .B(n_157), .Y(n_238) );
CKINVDCx11_ASAP7_75t_R g239 ( .A(n_169), .Y(n_239) );
AND3x1_ASAP7_75t_SL g240 ( .A(n_181), .B(n_72), .C(n_88), .Y(n_240) );
BUFx12f_ASAP7_75t_L g241 ( .A(n_181), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_212), .Y(n_242) );
OAI222xp33_ASAP7_75t_L g243 ( .A1(n_218), .A2(n_192), .B1(n_197), .B2(n_176), .C1(n_95), .C2(n_92), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
OAI222xp33_ASAP7_75t_L g246 ( .A1(n_218), .A2(n_92), .B1(n_95), .B2(n_174), .C1(n_89), .C2(n_177), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_225), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_218), .A2(n_193), .B1(n_160), .B2(n_157), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_211), .A2(n_129), .B1(n_127), .B2(n_166), .C(n_125), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_207), .A2(n_168), .B(n_194), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_236), .B(n_157), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_239), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_218), .A2(n_160), .B1(n_203), .B2(n_206), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_216), .A2(n_127), .B1(n_129), .B2(n_125), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_221), .A2(n_166), .B1(n_110), .B2(n_125), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_221), .A2(n_220), .B1(n_233), .B2(n_241), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_213), .B(n_175), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_212), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g261 ( .A1(n_217), .A2(n_110), .B1(n_206), .B2(n_203), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_236), .B(n_164), .Y(n_262) );
AND2x6_ASAP7_75t_L g263 ( .A(n_213), .B(n_175), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_224), .B(n_179), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
OAI21xp5_ASAP7_75t_SL g266 ( .A1(n_233), .A2(n_220), .B(n_224), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_266), .A2(n_265), .B1(n_245), .B2(n_247), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_262), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g269 ( .A1(n_266), .A2(n_226), .B1(n_234), .B2(n_237), .C(n_232), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_262), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_246), .A2(n_234), .B(n_232), .C(n_227), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_240), .B1(n_224), .B2(n_208), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_246), .A2(n_237), .B1(n_231), .B2(n_223), .C(n_224), .Y(n_273) );
OAI221xp5_ASAP7_75t_L g274 ( .A1(n_257), .A2(n_223), .B1(n_229), .B2(n_217), .C(n_228), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_245), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_247), .A2(n_217), .B1(n_241), .B2(n_208), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_250), .A2(n_230), .B(n_120), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_256), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_254), .Y(n_283) );
OAI221xp5_ASAP7_75t_L g284 ( .A1(n_248), .A2(n_229), .B1(n_228), .B2(n_238), .C(n_120), .Y(n_284) );
AOI22xp33_ASAP7_75t_SL g285 ( .A1(n_256), .A2(n_214), .B1(n_208), .B2(n_231), .Y(n_285) );
AOI22xp33_ASAP7_75t_SL g286 ( .A1(n_251), .A2(n_214), .B1(n_208), .B2(n_254), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_255), .B(n_208), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_251), .B(n_231), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_274), .B(n_276), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_275), .B(n_259), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_269), .A2(n_214), .B1(n_133), .B2(n_238), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_267), .B(n_214), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_269), .A2(n_214), .B1(n_133), .B2(n_249), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_274), .A2(n_133), .B1(n_249), .B2(n_263), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_273), .A2(n_253), .B1(n_120), .B2(n_250), .C(n_93), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_272), .A2(n_97), .B1(n_131), .B2(n_80), .C(n_79), .Y(n_296) );
OAI22xp33_ASAP7_75t_L g297 ( .A1(n_267), .A2(n_243), .B1(n_252), .B2(n_258), .Y(n_297) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_272), .A2(n_131), .B(n_230), .C(n_215), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g299 ( .A1(n_287), .A2(n_243), .B1(n_258), .B2(n_259), .Y(n_299) );
AOI222xp33_ASAP7_75t_L g300 ( .A1(n_279), .A2(n_263), .B1(n_261), .B2(n_160), .C1(n_112), .C2(n_131), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_275), .B(n_259), .Y(n_301) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_270), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_278), .A2(n_260), .B(n_244), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_275), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
OAI33xp33_ASAP7_75t_L g307 ( .A1(n_271), .A2(n_148), .A3(n_139), .B1(n_144), .B2(n_153), .B3(n_165), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_286), .A2(n_263), .B1(n_160), .B2(n_215), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_278), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_283), .B(n_259), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_283), .B(n_242), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_279), .B(n_242), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_284), .A2(n_258), .B(n_260), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_311), .B(n_281), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_304), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_304), .B(n_306), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_306), .B(n_268), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_305), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_305), .Y(n_320) );
OAI22xp5_ASAP7_75t_SL g321 ( .A1(n_289), .A2(n_285), .B1(n_287), .B2(n_280), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_311), .Y(n_322) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_309), .B(n_281), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_305), .B(n_282), .Y(n_324) );
OAI33xp33_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_282), .A3(n_144), .B1(n_148), .B2(n_153), .B3(n_139), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_297), .A2(n_288), .B1(n_270), .B2(n_280), .C(n_138), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_308), .B(n_288), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_308), .B(n_281), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_311), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_292), .A2(n_263), .B1(n_112), .B2(n_278), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_308), .B(n_278), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_1), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_299), .A2(n_263), .B1(n_112), .B2(n_244), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_296), .A2(n_138), .B1(n_136), .B2(n_145), .C(n_151), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_299), .A2(n_164), .B(n_189), .C(n_244), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_302), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_310), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_290), .B(n_242), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_3), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_290), .B(n_260), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
NOR2x1_ASAP7_75t_L g343 ( .A(n_298), .B(n_219), .Y(n_343) );
OAI31xp33_ASAP7_75t_SL g344 ( .A1(n_296), .A2(n_4), .A3(n_5), .B(n_6), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
OAI33xp33_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_4), .A3(n_6), .B1(n_7), .B2(n_9), .B3(n_10), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_290), .B(n_7), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_291), .A2(n_151), .B1(n_145), .B2(n_164), .C(n_138), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_301), .B(n_9), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_303), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
OAI31xp33_ASAP7_75t_L g353 ( .A1(n_295), .A2(n_179), .A3(n_184), .B(n_186), .Y(n_353) );
AND2x4_ASAP7_75t_SL g354 ( .A(n_326), .B(n_301), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_338), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_338), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_313), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_322), .B(n_313), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_318), .B(n_313), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_318), .B(n_302), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_345), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_352), .B(n_293), .Y(n_363) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_344), .A2(n_309), .B(n_295), .C(n_294), .Y(n_364) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_347), .B(n_307), .C(n_298), .Y(n_365) );
NAND4xp25_ASAP7_75t_SL g366 ( .A(n_337), .B(n_300), .C(n_314), .D(n_12), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_316), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_352), .B(n_314), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_317), .B(n_303), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_340), .B(n_303), .Y(n_372) );
OAI21xp33_ASAP7_75t_SL g373 ( .A1(n_326), .A2(n_300), .B(n_307), .Y(n_373) );
AND3x2_ASAP7_75t_L g374 ( .A(n_336), .B(n_10), .C(n_11), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_340), .B(n_11), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_348), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_333), .B(n_12), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_333), .B(n_209), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_348), .B(n_13), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_330), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_342), .B(n_14), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_350), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_339), .B(n_15), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
AOI211x1_ASAP7_75t_SL g387 ( .A1(n_328), .A2(n_17), .B(n_18), .C(n_19), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_346), .B(n_66), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_346), .B(n_20), .Y(n_389) );
AND2x6_ASAP7_75t_L g390 ( .A(n_343), .B(n_209), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_350), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_320), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_324), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_319), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_329), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_325), .B(n_145), .C(n_151), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_315), .B(n_20), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_321), .B(n_21), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_339), .B(n_341), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_323), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_341), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_315), .B(n_23), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_332), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_334), .B(n_27), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_392), .B(n_315), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_355), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_368), .B(n_315), .Y(n_408) );
NAND4xp75_ASAP7_75t_L g409 ( .A(n_398), .B(n_327), .C(n_343), .D(n_353), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_398), .B(n_336), .C(n_331), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_366), .B(n_321), .C(n_335), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_400), .B(n_351), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_378), .B(n_332), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_384), .B(n_323), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_373), .A2(n_351), .B(n_323), .C(n_349), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_391), .A2(n_138), .B1(n_187), .B2(n_200), .C(n_142), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_395), .B(n_263), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_365), .B(n_222), .C(n_212), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_393), .B(n_263), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_399), .B(n_32), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_376), .B(n_263), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g423 ( .A(n_383), .B(n_389), .C(n_364), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_382), .B(n_34), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_403), .A2(n_200), .B(n_142), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g426 ( .A(n_400), .B(n_36), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_379), .A2(n_209), .B1(n_219), .B2(n_184), .C(n_186), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_355), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_357), .B(n_37), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_359), .B(n_39), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_358), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_364), .B(n_196), .C(n_190), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_357), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_370), .B(n_44), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_360), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_372), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_354), .B(n_47), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_369), .B(n_48), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_381), .B(n_51), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_371), .B(n_52), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_394), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_385), .B(n_54), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_371), .B(n_56), .Y(n_446) );
INVx6_ASAP7_75t_L g447 ( .A(n_377), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_371), .B(n_57), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_354), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_356), .B(n_58), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_363), .B(n_60), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_356), .B(n_61), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_375), .B(n_62), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
OAI32xp33_ASAP7_75t_L g455 ( .A1(n_449), .A2(n_377), .A3(n_397), .B1(n_400), .B2(n_380), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_435), .B(n_361), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_436), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_438), .B(n_374), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_439), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_428), .B(n_361), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_419), .B(n_404), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_429), .B(n_362), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
OR2x6_ASAP7_75t_L g466 ( .A(n_447), .B(n_380), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_444), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_447), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_433), .B(n_362), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_413), .B(n_388), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_405), .B(n_388), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_414), .B(n_388), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_411), .A2(n_374), .B1(n_365), .B2(n_402), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_430), .B(n_390), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_447), .Y(n_477) );
NOR2xp33_ASAP7_75t_SL g478 ( .A(n_440), .B(n_390), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_416), .A2(n_396), .B(n_387), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_418), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_421), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_409), .B(n_390), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_423), .B(n_390), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_452), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_452), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_416), .B(n_390), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_410), .A2(n_396), .B1(n_209), .B2(n_222), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_431), .A2(n_112), .B1(n_210), .B2(n_212), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_423), .A2(n_142), .B1(n_190), .B2(n_235), .C(n_222), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_411), .B(n_222), .C(n_147), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_453), .A2(n_112), .B1(n_210), .B2(n_222), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_446), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_448), .Y(n_496) );
AOI211xp5_ASAP7_75t_L g497 ( .A1(n_426), .A2(n_64), .B(n_68), .C(n_112), .Y(n_497) );
NAND3xp33_ASAP7_75t_SL g498 ( .A(n_442), .B(n_210), .C(n_147), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_412), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_412), .B(n_210), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_412), .B(n_210), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_448), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_441), .B(n_210), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_445), .A2(n_147), .B1(n_205), .B2(n_451), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_450), .Y(n_507) );
AOI211xp5_ASAP7_75t_L g508 ( .A1(n_432), .A2(n_147), .B(n_205), .C(n_427), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_424), .Y(n_509) );
OAI31xp33_ASAP7_75t_L g510 ( .A1(n_425), .A2(n_147), .A3(n_205), .B(n_434), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_460), .A2(n_479), .B1(n_461), .B2(n_457), .C(n_468), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_458), .Y(n_512) );
AOI321xp33_ASAP7_75t_L g513 ( .A1(n_475), .A2(n_460), .A3(n_482), .B1(n_488), .B2(n_483), .C(n_455), .Y(n_513) );
OAI32xp33_ASAP7_75t_L g514 ( .A1(n_488), .A2(n_482), .A3(n_477), .B1(n_469), .B2(n_499), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_473), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_478), .A2(n_499), .B(n_466), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_SL g517 ( .A1(n_509), .A2(n_504), .B(n_497), .C(n_508), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_467), .B(n_459), .Y(n_518) );
NOR2x1p5_ASAP7_75t_L g519 ( .A(n_492), .B(n_472), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_466), .A2(n_463), .B(n_481), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_456), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_509), .A2(n_489), .B(n_510), .C(n_473), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_484), .A2(n_456), .B1(n_480), .B2(n_485), .C(n_470), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_514), .A2(n_470), .B1(n_462), .B2(n_464), .C(n_507), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_516), .A2(n_466), .B1(n_471), .B2(n_474), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_518), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_522), .A2(n_506), .B(n_503), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_520), .A2(n_502), .B1(n_494), .B2(n_496), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_511), .A2(n_498), .B(n_476), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_513), .B(n_491), .C(n_434), .Y(n_530) );
NOR4xp25_ASAP7_75t_L g531 ( .A(n_530), .B(n_518), .C(n_512), .D(n_523), .Y(n_531) );
NOR5xp2_ASAP7_75t_L g532 ( .A(n_527), .B(n_517), .C(n_519), .D(n_503), .E(n_495), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_525), .A2(n_521), .B1(n_515), .B2(n_487), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_529), .B(n_476), .Y(n_534) );
NAND3x1_ASAP7_75t_L g535 ( .A(n_532), .B(n_524), .C(n_526), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_534), .A2(n_528), .B1(n_486), .B2(n_470), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_535), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g538 ( .A1(n_536), .A2(n_531), .B1(n_533), .B2(n_465), .C(n_454), .Y(n_538) );
NOR3xp33_ASAP7_75t_SL g539 ( .A(n_537), .B(n_417), .C(n_505), .Y(n_539) );
AOI222xp33_ASAP7_75t_SL g540 ( .A1(n_539), .A2(n_538), .B1(n_454), .B2(n_465), .C1(n_490), .C2(n_493), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g541 ( .A(n_540), .B(n_464), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_541), .A2(n_500), .B(n_501), .Y(n_542) );
endmodule