module fake_netlist_6_146_n_1381 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1381);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1381;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_1368;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_10),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_204),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_47),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_171),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_13),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_161),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_117),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_31),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_229),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_182),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_19),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_103),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_147),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_74),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_26),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_222),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_279),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_86),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_278),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_99),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_215),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_169),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_137),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_350),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_330),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_4),
.B(n_295),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_86),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_353),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_116),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_254),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_277),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_76),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_271),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_203),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_135),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_56),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_162),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_142),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_139),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_157),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_5),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_173),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_246),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_294),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_25),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_130),
.Y(n_431)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_175),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_184),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_248),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_302),
.B(n_211),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_220),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_92),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_67),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_158),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_247),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_202),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_293),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_336),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_2),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_115),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_122),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_165),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_331),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_326),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_28),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_319),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_356),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_250),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_15),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_138),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_5),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_29),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_269),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_314),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_273),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_299),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_275),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_16),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_32),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_136),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_301),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_333),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_327),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_45),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_124),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_197),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_33),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_195),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_186),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_149),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_47),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_216),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_205),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_258),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_292),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_113),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_223),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_259),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_316),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_20),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_196),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_263),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_36),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_360),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_123),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_305),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_99),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_357),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_213),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_201),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_192),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_272),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_112),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_239),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_168),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_44),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_174),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_317),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_361),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_9),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_88),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_340),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_152),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_200),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_318),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_2),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_183),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_179),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_321),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_134),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_181),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_9),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_84),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_90),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_87),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_90),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_63),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_371),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_210),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_34),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_27),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_238),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_219),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_106),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_240),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_354),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_312),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_343),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_266),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_224),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_148),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_32),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_315),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_297),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_73),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_26),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_73),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_337),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_280),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_303),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_42),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_17),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_281),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_226),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_145),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_389),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_477),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_413),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_502),
.B(n_0),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_420),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_401),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_389),
.Y(n_559)
);

OA22x2_ASAP7_75t_SL g560 ( 
.A1(n_383),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_486),
.A2(n_437),
.B1(n_527),
.B2(n_416),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_421),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_421),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_379),
.A2(n_6),
.B(n_7),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_422),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_422),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_447),
.B(n_8),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_380),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_10),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_420),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_422),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_405),
.B(n_11),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_422),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_542),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_389),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_405),
.B(n_12),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_469),
.B(n_14),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_392),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_378),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_480),
.B(n_14),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_389),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_476),
.B(n_15),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_438),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_16),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_380),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_389),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_17),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_389),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_432),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_476),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_493),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_513),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_396),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_406),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_411),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_444),
.Y(n_601)
);

BUFx12f_ASAP7_75t_L g602 ( 
.A(n_376),
.Y(n_602)
);

OAI22x1_ASAP7_75t_R g603 ( 
.A1(n_382),
.A2(n_386),
.B1(n_393),
.B2(n_388),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_432),
.Y(n_604)
);

OA21x2_ASAP7_75t_L g605 ( 
.A1(n_381),
.A2(n_18),
.B(n_19),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_526),
.A2(n_464),
.B1(n_465),
.B2(n_457),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_473),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_469),
.B(n_18),
.Y(n_608)
);

AOI22x1_ASAP7_75t_SL g609 ( 
.A1(n_398),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_526),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_610)
);

OA21x2_ASAP7_75t_L g611 ( 
.A1(n_384),
.A2(n_23),
.B(n_24),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_432),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_441),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_489),
.Y(n_614)
);

BUFx8_ASAP7_75t_SL g615 ( 
.A(n_387),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_495),
.B(n_467),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_499),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_377),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_519),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_546),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_432),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_533),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_400),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_443),
.B(n_30),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_390),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_391),
.B(n_394),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_541),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_603),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_556),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_584),
.B(n_409),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_616),
.B(n_481),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_556),
.Y(n_635)
);

CKINVDCx6p67_ASAP7_75t_R g636 ( 
.A(n_595),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_587),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_618),
.B(n_481),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_562),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_562),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_557),
.Y(n_642)
);

INVx8_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_598),
.Y(n_644)
);

NOR2x1p5_ASAP7_75t_L g645 ( 
.A(n_557),
.B(n_435),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_582),
.B(n_608),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_582),
.B(n_546),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_598),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_563),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_564),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_616),
.B(n_508),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_566),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_594),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_567),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_572),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_579),
.B(n_423),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_572),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_555),
.A2(n_570),
.B1(n_571),
.B2(n_628),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_572),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_577),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_577),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_598),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_591),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_587),
.B(n_428),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_578),
.B(n_430),
.C(n_426),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_599),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_593),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_597),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_597),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_637),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_596),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_632),
.A2(n_410),
.B1(n_434),
.B2(n_385),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_646),
.B(n_628),
.Y(n_681)
);

AO22x2_ASAP7_75t_L g682 ( 
.A1(n_660),
.A2(n_621),
.B1(n_560),
.B2(n_609),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_647),
.B(n_552),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_656),
.B(n_596),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_645),
.B(n_662),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_644),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_631),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_653),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_669),
.A2(n_554),
.B1(n_571),
.B2(n_625),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_634),
.B(n_559),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_633),
.B(n_574),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_656),
.B(n_558),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_638),
.B(n_573),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_633),
.B(n_613),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_666),
.B(n_613),
.Y(n_695)
);

AND2x6_ASAP7_75t_SL g696 ( 
.A(n_630),
.B(n_626),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_634),
.B(n_576),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_643),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_670),
.B(n_602),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_635),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_639),
.B(n_583),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_652),
.B(n_615),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_632),
.B(n_569),
.Y(n_703)
);

NOR2xp67_ASAP7_75t_L g704 ( 
.A(n_649),
.B(n_553),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_636),
.A2(n_610),
.B1(n_575),
.B2(n_621),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_673),
.B(n_626),
.Y(n_706)
);

AND2x4_ASAP7_75t_SL g707 ( 
.A(n_636),
.B(n_561),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_639),
.B(n_568),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_657),
.B(n_624),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_651),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_661),
.B(n_586),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_651),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_651),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_664),
.B(n_597),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_665),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_665),
.A2(n_560),
.B1(n_589),
.B2(n_543),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_668),
.B(n_589),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_640),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_648),
.B(n_442),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_671),
.A2(n_452),
.B1(n_472),
.B2(n_471),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_641),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_641),
.B(n_397),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_515),
.B1(n_505),
.B2(n_606),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_650),
.B(n_588),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_650),
.B(n_590),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_672),
.A2(n_606),
.B1(n_622),
.B2(n_617),
.C(n_575),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_654),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_654),
.B(n_592),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_675),
.B(n_627),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_677),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_681),
.A2(n_443),
.B(n_483),
.C(n_622),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_678),
.B(n_561),
.Y(n_734)
);

AND2x2_ASAP7_75t_SL g735 ( 
.A(n_707),
.B(n_610),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_693),
.B(n_655),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_686),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_679),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_684),
.B(n_553),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_703),
.B(n_440),
.Y(n_740)
);

BUFx12f_ASAP7_75t_L g741 ( 
.A(n_696),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_691),
.A2(n_659),
.B(n_658),
.Y(n_742)
);

OAI21xp5_ASAP7_75t_L g743 ( 
.A1(n_683),
.A2(n_605),
.B(n_565),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_683),
.B(n_658),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_681),
.B(n_483),
.Y(n_746)
);

OR2x6_ASAP7_75t_SL g747 ( 
.A(n_689),
.B(n_705),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_718),
.A2(n_605),
.B(n_565),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_685),
.B(n_611),
.C(n_402),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_680),
.B(n_611),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_722),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_690),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_706),
.B(n_403),
.C(n_395),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_708),
.B(n_659),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_711),
.A2(n_667),
.B(n_663),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_690),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_728),
.B(n_674),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_697),
.Y(n_758)
);

AOI21x1_ASAP7_75t_L g759 ( 
.A1(n_701),
.A2(n_677),
.B(n_676),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_732),
.Y(n_760)
);

BUFx4f_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_695),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_719),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_687),
.B(n_688),
.Y(n_764)
);

AOI22x1_ASAP7_75t_L g765 ( 
.A1(n_717),
.A2(n_612),
.B1(n_623),
.B2(n_604),
.Y(n_765)
);

INVx11_ASAP7_75t_L g766 ( 
.A(n_699),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_725),
.A2(n_415),
.B(n_414),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_689),
.A2(n_600),
.B(n_601),
.C(n_580),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_725),
.A2(n_729),
.B(n_726),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_720),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_721),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_726),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_716),
.B(n_424),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_692),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_705),
.B(n_494),
.C(n_468),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_730),
.B(n_425),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_700),
.B(n_427),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_723),
.A2(n_619),
.B(n_620),
.C(n_607),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_724),
.A2(n_702),
.B1(n_727),
.B2(n_682),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_710),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_712),
.B(n_713),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_682),
.A2(n_528),
.B1(n_549),
.B2(n_517),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_714),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_709),
.B(n_431),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_731),
.B(n_445),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_704),
.B(n_629),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_698),
.B(n_399),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_683),
.A2(n_451),
.B(n_449),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_693),
.B(n_455),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_694),
.A2(n_478),
.B(n_461),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_694),
.A2(n_500),
.B(n_488),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_703),
.B(n_404),
.Y(n_792)
);

BUFx12f_ASAP7_75t_L g793 ( 
.A(n_678),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_681),
.A2(n_503),
.B(n_509),
.C(n_501),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_693),
.B(n_516),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_693),
.B(n_118),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_703),
.B(n_529),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_678),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_693),
.B(n_531),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_694),
.A2(n_535),
.B(n_534),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_694),
.A2(n_540),
.B(n_539),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_694),
.A2(n_550),
.B(n_545),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_690),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_693),
.B(n_407),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_683),
.A2(n_412),
.B(n_408),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_694),
.A2(n_418),
.B(n_417),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_693),
.B(n_419),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_693),
.A2(n_614),
.B(n_433),
.C(n_436),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_693),
.B(n_429),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_693),
.A2(n_614),
.B1(n_454),
.B2(n_458),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_693),
.B(n_439),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_693),
.B(n_446),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_693),
.A2(n_453),
.B(n_456),
.C(n_448),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_703),
.B(n_450),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_715),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_678),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_694),
.A2(n_460),
.B(n_459),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_686),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_693),
.A2(n_463),
.B(n_466),
.C(n_462),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_693),
.B(n_474),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_683),
.A2(n_479),
.B(n_475),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_678),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_693),
.B(n_484),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_822),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_743),
.A2(n_769),
.B(n_749),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_743),
.A2(n_490),
.B(n_487),
.Y(n_826)
);

OAI22x1_ASAP7_75t_L g827 ( 
.A1(n_771),
.A2(n_482),
.B1(n_506),
.B2(n_470),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_746),
.B(n_491),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_796),
.A2(n_496),
.B1(n_497),
.B2(n_492),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_737),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_738),
.B(n_585),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_762),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_744),
.A2(n_504),
.B(n_498),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_755),
.A2(n_585),
.B(n_581),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_754),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_752),
.A2(n_514),
.B(n_510),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_759),
.A2(n_581),
.B(n_120),
.Y(n_837)
);

OAI21x1_ASAP7_75t_SL g838 ( 
.A1(n_765),
.A2(n_121),
.B(n_119),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_762),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_737),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_816),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_749),
.A2(n_525),
.B(n_524),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_756),
.A2(n_536),
.B(n_532),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_804),
.B(n_537),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_738),
.B(n_512),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_764),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_758),
.A2(n_551),
.B(n_544),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_789),
.A2(n_522),
.B1(n_523),
.B2(n_521),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_807),
.B(n_530),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_788),
.A2(n_547),
.B(n_538),
.C(n_36),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_809),
.B(n_34),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_734),
.B(n_35),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_811),
.B(n_35),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_780),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_748),
.A2(n_126),
.B(n_125),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_750),
.A2(n_775),
.B1(n_779),
.B2(n_821),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_793),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_SL g858 ( 
.A1(n_782),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.C(n_40),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_747),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_812),
.B(n_37),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_795),
.A2(n_128),
.B1(n_129),
.B2(n_127),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_742),
.A2(n_375),
.B(n_132),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_739),
.B(n_38),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_815),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_820),
.B(n_39),
.Y(n_865)
);

NAND3xp33_ASAP7_75t_L g866 ( 
.A(n_821),
.B(n_40),
.C(n_41),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_772),
.A2(n_133),
.B(n_131),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_760),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_799),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_823),
.B(n_43),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_741),
.B(n_44),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_803),
.A2(n_141),
.B(n_140),
.Y(n_872)
);

OAI22x1_ASAP7_75t_L g873 ( 
.A1(n_770),
.A2(n_774),
.B1(n_735),
.B2(n_740),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_781),
.A2(n_144),
.B(n_143),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_774),
.B(n_45),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_780),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_736),
.B(n_46),
.Y(n_877)
);

INVxp67_ASAP7_75t_SL g878 ( 
.A(n_737),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_745),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_783),
.B(n_48),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_761),
.B(n_146),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_805),
.B(n_48),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_810),
.B(n_49),
.Y(n_883)
);

AOI221x1_ASAP7_75t_L g884 ( 
.A1(n_808),
.A2(n_153),
.B1(n_154),
.B2(n_151),
.C(n_150),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_797),
.B(n_49),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_813),
.A2(n_156),
.B(n_155),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_733),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_761),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_792),
.A2(n_160),
.B(n_159),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_785),
.B(n_50),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_819),
.A2(n_164),
.B(n_163),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_757),
.Y(n_892)
);

AO31x2_ASAP7_75t_L g893 ( 
.A1(n_790),
.A2(n_53),
.A3(n_51),
.B(n_52),
.Y(n_893)
);

OA21x2_ASAP7_75t_L g894 ( 
.A1(n_784),
.A2(n_167),
.B(n_166),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_753),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_895)
);

NAND3x1_ASAP7_75t_L g896 ( 
.A(n_776),
.B(n_54),
.C(n_55),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_751),
.B(n_56),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_786),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_818),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_768),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_900)
);

AO31x2_ASAP7_75t_L g901 ( 
.A1(n_791),
.A2(n_61),
.A3(n_59),
.B(n_60),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_773),
.A2(n_172),
.B1(n_176),
.B2(n_170),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_777),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_766),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_806),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_817),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_800),
.B(n_801),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_802),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_767),
.B(n_177),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_787),
.A2(n_180),
.B(n_178),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_778),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_794),
.A2(n_187),
.B(n_185),
.Y(n_912)
);

AND3x4_ASAP7_75t_L g913 ( 
.A(n_775),
.B(n_60),
.C(n_61),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_746),
.B(n_62),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_793),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_737),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_737),
.Y(n_917)
);

OA22x2_ASAP7_75t_L g918 ( 
.A1(n_779),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_L g919 ( 
.A(n_814),
.B(n_64),
.C(n_65),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_754),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_746),
.B(n_65),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_743),
.A2(n_189),
.B(n_188),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_822),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_788),
.A2(n_66),
.B(n_67),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_746),
.B(n_66),
.Y(n_925)
);

AND3x2_ASAP7_75t_L g926 ( 
.A(n_822),
.B(n_68),
.C(n_69),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_779),
.B(n_68),
.C(n_69),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_746),
.B(n_70),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_738),
.B(n_190),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_746),
.A2(n_193),
.B1(n_194),
.B2(n_191),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_746),
.B(n_70),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_822),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_746),
.B(n_71),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_796),
.A2(n_255),
.B1(n_373),
.B2(n_370),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_754),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_SL g936 ( 
.A(n_775),
.B(n_71),
.C(n_72),
.Y(n_936)
);

OAI21xp33_ASAP7_75t_L g937 ( 
.A1(n_746),
.A2(n_72),
.B(n_74),
.Y(n_937)
);

AO21x1_ASAP7_75t_L g938 ( 
.A1(n_788),
.A2(n_75),
.B(n_76),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_754),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_746),
.B(n_75),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_769),
.A2(n_199),
.B(n_198),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_796),
.A2(n_257),
.B1(n_369),
.B2(n_368),
.Y(n_942)
);

AO31x2_ASAP7_75t_L g943 ( 
.A1(n_746),
.A2(n_77),
.A3(n_78),
.B(n_79),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_746),
.B(n_77),
.Y(n_944)
);

AO31x2_ASAP7_75t_L g945 ( 
.A1(n_746),
.A2(n_79),
.A3(n_80),
.B(n_81),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_746),
.B(n_80),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_737),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_763),
.Y(n_948)
);

AO21x1_ASAP7_75t_L g949 ( 
.A1(n_788),
.A2(n_81),
.B(n_82),
.Y(n_949)
);

OA21x2_ASAP7_75t_L g950 ( 
.A1(n_743),
.A2(n_207),
.B(n_206),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_798),
.B(n_208),
.Y(n_951)
);

O2A1O1Ixp5_ASAP7_75t_L g952 ( 
.A1(n_788),
.A2(n_264),
.B(n_366),
.C(n_365),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_746),
.B(n_82),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_746),
.A2(n_262),
.B1(n_364),
.B2(n_362),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_745),
.B(n_209),
.Y(n_955)
);

AO31x2_ASAP7_75t_L g956 ( 
.A1(n_746),
.A2(n_83),
.A3(n_84),
.B(n_85),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_746),
.B(n_83),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_743),
.A2(n_214),
.B(n_212),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_746),
.B(n_85),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_754),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_824),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_825),
.A2(n_218),
.B(n_217),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_856),
.A2(n_274),
.B1(n_359),
.B2(n_358),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_932),
.B(n_87),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_868),
.Y(n_965)
);

OA21x2_ASAP7_75t_L g966 ( 
.A1(n_837),
.A2(n_225),
.B(n_221),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_864),
.Y(n_967)
);

AO21x2_ASAP7_75t_L g968 ( 
.A1(n_855),
.A2(n_228),
.B(n_227),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_883),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_SL g970 ( 
.A(n_888),
.B(n_89),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_851),
.A2(n_276),
.B(n_355),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_882),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_SL g973 ( 
.A1(n_859),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_846),
.B(n_94),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_SL g975 ( 
.A1(n_913),
.A2(n_95),
.B(n_96),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_835),
.B(n_97),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_922),
.A2(n_282),
.B(n_352),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_888),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_853),
.A2(n_270),
.B(n_349),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_828),
.A2(n_268),
.B1(n_348),
.B2(n_346),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_860),
.A2(n_267),
.B(n_345),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_888),
.B(n_916),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_857),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_923),
.B(n_97),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_845),
.B(n_98),
.C(n_100),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_865),
.A2(n_265),
.B(n_344),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_870),
.A2(n_261),
.B(n_342),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_854),
.A2(n_283),
.B1(n_341),
.B2(n_338),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_914),
.A2(n_98),
.B(n_100),
.C(n_101),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_921),
.A2(n_101),
.B(n_102),
.C(n_104),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_920),
.B(n_104),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_854),
.A2(n_285),
.B1(n_335),
.B2(n_334),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_948),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_849),
.B(n_105),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_841),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_873),
.A2(n_260),
.B1(n_332),
.B2(n_329),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_958),
.A2(n_256),
.B(n_324),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_935),
.B(n_105),
.Y(n_998)
);

CKINVDCx14_ASAP7_75t_R g999 ( 
.A(n_915),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_939),
.B(n_106),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_876),
.A2(n_284),
.B1(n_323),
.B2(n_320),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_916),
.B(n_253),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_890),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_904),
.Y(n_1004)
);

OAI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_925),
.A2(n_931),
.B1(n_959),
.B2(n_944),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_852),
.B(n_108),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_928),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_1007)
);

OA21x2_ASAP7_75t_L g1008 ( 
.A1(n_867),
.A2(n_252),
.B(n_313),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_898),
.B(n_110),
.Y(n_1009)
);

OA21x2_ASAP7_75t_L g1010 ( 
.A1(n_872),
.A2(n_286),
.B(n_311),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_L g1011 ( 
.A(n_933),
.B(n_111),
.C(n_112),
.Y(n_1011)
);

OA21x2_ASAP7_75t_L g1012 ( 
.A1(n_886),
.A2(n_287),
.B(n_310),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_SL g1013 ( 
.A1(n_838),
.A2(n_251),
.B(n_308),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_960),
.A2(n_249),
.B1(n_307),
.B2(n_306),
.Y(n_1014)
);

OA21x2_ASAP7_75t_L g1015 ( 
.A1(n_891),
.A2(n_245),
.B(n_304),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_875),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_862),
.A2(n_244),
.B(n_300),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_899),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_955),
.B(n_243),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_831),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_892),
.B(n_113),
.Y(n_1021)
);

BUFx2_ASAP7_75t_R g1022 ( 
.A(n_905),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_880),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_940),
.B(n_114),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_903),
.B(n_114),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_832),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_830),
.Y(n_1027)
);

INVx6_ASAP7_75t_L g1028 ( 
.A(n_917),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_955),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_946),
.A2(n_117),
.B(n_230),
.C(n_231),
.Y(n_1030)
);

INVx6_ASAP7_75t_L g1031 ( 
.A(n_917),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_953),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_917),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_947),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_918),
.B(n_947),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_877),
.A2(n_235),
.B(n_236),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_879),
.Y(n_1037)
);

BUFx8_ASAP7_75t_L g1038 ( 
.A(n_897),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_957),
.B(n_367),
.Y(n_1039)
);

CKINVDCx11_ASAP7_75t_R g1040 ( 
.A(n_871),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_908),
.A2(n_237),
.B(n_241),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_839),
.B(n_242),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_826),
.A2(n_289),
.B(n_290),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_863),
.B(n_291),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_947),
.B(n_296),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_840),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_844),
.B(n_298),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_937),
.A2(n_848),
.B(n_850),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_934),
.B(n_942),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_866),
.A2(n_927),
.B1(n_924),
.B2(n_949),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_911),
.A2(n_906),
.B1(n_878),
.B2(n_912),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_836),
.B(n_847),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_843),
.B(n_885),
.Y(n_1053)
);

BUFx2_ASAP7_75t_R g1054 ( 
.A(n_929),
.Y(n_1054)
);

AO21x1_ASAP7_75t_L g1055 ( 
.A1(n_941),
.A2(n_930),
.B(n_954),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_827),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_842),
.B(n_936),
.Y(n_1057)
);

NOR4xp25_ASAP7_75t_L g1058 ( 
.A(n_900),
.B(n_919),
.C(n_869),
.D(n_887),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_938),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_833),
.B(n_951),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_884),
.A2(n_952),
.B(n_858),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_911),
.B(n_829),
.Y(n_1062)
);

OAI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_881),
.A2(n_911),
.B1(n_871),
.B2(n_861),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_895),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_907),
.A2(n_950),
.B1(n_909),
.B2(n_896),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_943),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_874),
.A2(n_889),
.B(n_910),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_943),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_902),
.A2(n_894),
.B(n_926),
.C(n_945),
.Y(n_1069)
);

AOI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_894),
.A2(n_945),
.B(n_956),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_893),
.A2(n_856),
.B1(n_846),
.B2(n_796),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_901),
.A2(n_746),
.B(n_856),
.C(n_814),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_901),
.B(n_824),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_856),
.A2(n_779),
.B1(n_883),
.B2(n_882),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_859),
.B(n_678),
.Y(n_1075)
);

AO32x2_ASAP7_75t_L g1076 ( 
.A1(n_930),
.A2(n_779),
.A3(n_782),
.B1(n_621),
.B2(n_689),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_846),
.B(n_738),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_824),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_824),
.B(n_932),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_846),
.B(n_738),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_824),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_831),
.B(n_678),
.Y(n_1082)
);

OA21x2_ASAP7_75t_L g1083 ( 
.A1(n_825),
.A2(n_834),
.B(n_743),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_856),
.A2(n_779),
.B1(n_883),
.B2(n_882),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_967),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1082),
.B(n_1020),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_1075),
.B(n_1080),
.Y(n_1087)
);

OAI222xp33_ASAP7_75t_L g1088 ( 
.A1(n_1074),
.A2(n_1084),
.B1(n_969),
.B2(n_1003),
.C1(n_1057),
.C2(n_973),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1023),
.B(n_1005),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1016),
.B(n_1035),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_982),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_993),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_1078),
.B(n_1079),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1081),
.B(n_961),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1026),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_SL g1096 ( 
.A1(n_1024),
.A2(n_1056),
.B1(n_994),
.B2(n_1019),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1048),
.A2(n_1049),
.B1(n_985),
.B2(n_1011),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1021),
.Y(n_1098)
);

INVx6_ASAP7_75t_L g1099 ( 
.A(n_978),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_1072),
.A2(n_1071),
.B(n_1043),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1064),
.B(n_1053),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1059),
.B(n_1019),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1027),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1022),
.B(n_1006),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_SL g1105 ( 
.A(n_1038),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1027),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1077),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1046),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_978),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_974),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_976),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1018),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_995),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_991),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_989),
.A2(n_1007),
.B(n_972),
.C(n_990),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_965),
.Y(n_1116)
);

BUFx4_ASAP7_75t_R g1117 ( 
.A(n_1029),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_999),
.Y(n_1118)
);

BUFx2_ASAP7_75t_SL g1119 ( 
.A(n_1037),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1046),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_998),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1065),
.A2(n_1051),
.B(n_1066),
.Y(n_1122)
);

CKINVDCx6p67_ASAP7_75t_R g1123 ( 
.A(n_983),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1000),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1068),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1047),
.B(n_1044),
.Y(n_1126)
);

BUFx2_ASAP7_75t_SL g1127 ( 
.A(n_983),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1025),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1049),
.A2(n_1063),
.B1(n_1050),
.B2(n_963),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1033),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1034),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_975),
.B(n_1009),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_984),
.B(n_1039),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1058),
.B(n_1052),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1028),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1028),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_1004),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1062),
.B(n_1061),
.Y(n_1138)
);

AO21x1_ASAP7_75t_L g1139 ( 
.A1(n_1069),
.A2(n_1036),
.B(n_979),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1042),
.B(n_996),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1038),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1031),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1031),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1073),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1002),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1076),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1076),
.Y(n_1147)
);

BUFx4f_ASAP7_75t_L g1148 ( 
.A(n_964),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1076),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_964),
.B(n_1054),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1045),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1061),
.B(n_1060),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_970),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1083),
.B(n_971),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1030),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_981),
.B(n_987),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1040),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_986),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1013),
.Y(n_1159)
);

OR2x2_ASAP7_75t_SL g1160 ( 
.A(n_1012),
.B(n_1015),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_968),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_977),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1055),
.A2(n_1012),
.B1(n_1015),
.B2(n_980),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_977),
.B(n_997),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1032),
.B(n_1010),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1041),
.B(n_1067),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1017),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_997),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_SL g1169 ( 
.A1(n_962),
.A2(n_1014),
.B(n_1001),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_988),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_992),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_966),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1008),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1008),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1019),
.B(n_1079),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_1072),
.A2(n_1070),
.B(n_1071),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1137),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1086),
.B(n_1132),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1125),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1085),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1175),
.B(n_1103),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1087),
.B(n_1098),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1093),
.B(n_1116),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1108),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1175),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1096),
.B(n_1090),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1092),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1114),
.B(n_1121),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1096),
.B(n_1106),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1120),
.B(n_1104),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1099),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1118),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1124),
.B(n_1128),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1099),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1089),
.B(n_1101),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1116),
.B(n_1133),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1144),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1089),
.B(n_1102),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1134),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1129),
.A2(n_1126),
.B1(n_1158),
.B2(n_1097),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1102),
.B(n_1107),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1139),
.A2(n_1168),
.A3(n_1164),
.B(n_1173),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1095),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1099),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1138),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1152),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_1123),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1138),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1143),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1143),
.Y(n_1212)
);

OAI322xp33_ASAP7_75t_L g1213 ( 
.A1(n_1126),
.A2(n_1115),
.A3(n_1101),
.B1(n_1147),
.B2(n_1149),
.C1(n_1146),
.C2(n_1155),
.Y(n_1213)
);

OR2x6_ASAP7_75t_L g1214 ( 
.A(n_1145),
.B(n_1140),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1097),
.B(n_1094),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1112),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1130),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1119),
.B(n_1150),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1113),
.B(n_1129),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1153),
.B(n_1151),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1131),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1091),
.B(n_1135),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1112),
.B(n_1136),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1135),
.B(n_1156),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1100),
.A2(n_1140),
.B1(n_1171),
.B2(n_1170),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1159),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1122),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1162),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1148),
.B(n_1142),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1088),
.B(n_1100),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1115),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1143),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1172),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1109),
.B(n_1148),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1162),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1127),
.B(n_1109),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1165),
.B(n_1176),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1141),
.B(n_1157),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1157),
.B(n_1118),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1233),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1214),
.B(n_1166),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1201),
.B(n_1176),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1233),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1185),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1179),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1214),
.B(n_1166),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1228),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1187),
.B(n_1154),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1179),
.Y(n_1249)
);

NOR2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1219),
.B(n_1105),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1180),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1207),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1207),
.Y(n_1253)
);

NOR2xp67_ASAP7_75t_L g1254 ( 
.A(n_1177),
.B(n_1189),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1210),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1230),
.B(n_1208),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1237),
.B(n_1160),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1214),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1185),
.B(n_1167),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1195),
.B(n_1169),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1183),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1230),
.B(n_1174),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1193),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1202),
.A2(n_1163),
.B1(n_1161),
.B2(n_1088),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1228),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1191),
.B(n_1161),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1225),
.B(n_1163),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1182),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1188),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1235),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_R g1271 ( 
.A(n_1194),
.B(n_1105),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1204),
.B(n_1184),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1205),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1215),
.B(n_1117),
.Y(n_1274)
);

INVxp33_ASAP7_75t_L g1275 ( 
.A(n_1274),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1257),
.B(n_1198),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1247),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1240),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1257),
.B(n_1224),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1247),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1256),
.B(n_1262),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1262),
.B(n_1227),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1242),
.B(n_1227),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1265),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1242),
.B(n_1186),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1261),
.B(n_1199),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1260),
.B(n_1200),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1245),
.B(n_1199),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1265),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1240),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1270),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1270),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1243),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1249),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1252),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1252),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1253),
.Y(n_1297)
);

NOR2xp67_ASAP7_75t_SL g1298 ( 
.A(n_1244),
.B(n_1190),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1258),
.B(n_1226),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1266),
.B(n_1231),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1266),
.B(n_1192),
.Y(n_1301)
);

AND2x4_ASAP7_75t_SL g1302 ( 
.A(n_1259),
.B(n_1181),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1268),
.B(n_1197),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1253),
.B(n_1203),
.Y(n_1304)
);

AND2x4_ASAP7_75t_SL g1305 ( 
.A(n_1259),
.B(n_1181),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1279),
.B(n_1248),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1291),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1295),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1287),
.B(n_1255),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1275),
.B(n_1216),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1278),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1291),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1281),
.B(n_1285),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1275),
.B(n_1276),
.Y(n_1314)
);

OAI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1303),
.A2(n_1254),
.B1(n_1264),
.B2(n_1286),
.C(n_1234),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1296),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1290),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1297),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1290),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1301),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1281),
.B(n_1272),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1285),
.B(n_1272),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1293),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1300),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1277),
.B(n_1255),
.Y(n_1325)
);

OAI221xp5_ASAP7_75t_L g1326 ( 
.A1(n_1300),
.A2(n_1223),
.B1(n_1220),
.B2(n_1169),
.C(n_1218),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1312),
.B(n_1241),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1324),
.B(n_1282),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1320),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1310),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1322),
.B(n_1282),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1315),
.A2(n_1299),
.B(n_1294),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1326),
.A2(n_1241),
.B1(n_1246),
.B2(n_1250),
.Y(n_1333)
);

O2A1O1Ixp5_ASAP7_75t_L g1334 ( 
.A1(n_1309),
.A2(n_1298),
.B(n_1213),
.C(n_1299),
.Y(n_1334)
);

OAI322xp33_ASAP7_75t_L g1335 ( 
.A1(n_1306),
.A2(n_1288),
.A3(n_1304),
.B1(n_1280),
.B2(n_1284),
.C1(n_1292),
.C2(n_1289),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1307),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1312),
.B(n_1241),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1314),
.B(n_1283),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1313),
.B(n_1283),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1311),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1325),
.A2(n_1267),
.B(n_1246),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1311),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1340),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1342),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1327),
.Y(n_1345)
);

AOI31xp33_ASAP7_75t_L g1346 ( 
.A1(n_1332),
.A2(n_1271),
.A3(n_1194),
.B(n_1239),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1336),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_SL g1348 ( 
.A(n_1341),
.B(n_1190),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1333),
.A2(n_1318),
.B1(n_1308),
.B2(n_1316),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1331),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1347),
.B(n_1329),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1346),
.B(n_1330),
.Y(n_1352)
);

AOI331xp33_ASAP7_75t_L g1353 ( 
.A1(n_1344),
.A2(n_1334),
.A3(n_1319),
.B1(n_1323),
.B2(n_1317),
.B3(n_1269),
.C1(n_1251),
.Y(n_1353)
);

AOI221xp5_ASAP7_75t_L g1354 ( 
.A1(n_1349),
.A2(n_1335),
.B1(n_1338),
.B2(n_1328),
.C(n_1325),
.Y(n_1354)
);

OAI222xp33_ASAP7_75t_L g1355 ( 
.A1(n_1348),
.A2(n_1345),
.B1(n_1350),
.B2(n_1337),
.C1(n_1327),
.C2(n_1339),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_L g1356 ( 
.A(n_1352),
.B(n_1343),
.Y(n_1356)
);

NOR2x1_ASAP7_75t_L g1357 ( 
.A(n_1355),
.B(n_1343),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1351),
.Y(n_1358)
);

OAI211xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1354),
.A2(n_1345),
.B(n_1222),
.C(n_1273),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1353),
.A2(n_1305),
.B1(n_1302),
.B2(n_1337),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1352),
.A2(n_1325),
.B(n_1299),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1356),
.B(n_1313),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1358),
.B(n_1321),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1361),
.B(n_1360),
.C(n_1357),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1363),
.Y(n_1365)
);

NOR2xp67_ASAP7_75t_SL g1366 ( 
.A(n_1362),
.B(n_1209),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1365),
.B(n_1238),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1367),
.A2(n_1209),
.B1(n_1364),
.B2(n_1366),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1368),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1368),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1370),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1369),
.B(n_1178),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1371),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1372),
.Y(n_1374)
);

XNOR2xp5_ASAP7_75t_L g1375 ( 
.A(n_1374),
.B(n_1229),
.Y(n_1375)
);

AOI221x1_ASAP7_75t_L g1376 ( 
.A1(n_1373),
.A2(n_1359),
.B1(n_1232),
.B2(n_1212),
.C(n_1236),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1375),
.A2(n_1211),
.B(n_1221),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1376),
.A2(n_1117),
.B(n_1217),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1377),
.B(n_1193),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1378),
.A2(n_1212),
.B1(n_1232),
.B2(n_1206),
.C(n_1196),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1380),
.A2(n_1379),
.B1(n_1263),
.B2(n_1232),
.Y(n_1381)
);


endmodule