module fake_netlist_6_1593_n_254 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_32, n_66, n_78, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_27, n_38, n_61, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_41, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_254);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_32;
input n_66;
input n_78;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_27;
input n_38;
input n_61;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_41;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_254;

wire n_91;
wire n_146;
wire n_119;
wire n_163;
wire n_235;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_209;
wire n_98;
wire n_113;
wire n_223;
wire n_148;
wire n_199;
wire n_138;
wire n_161;
wire n_208;
wire n_226;
wire n_228;
wire n_252;
wire n_166;
wire n_184;
wire n_212;
wire n_158;
wire n_217;
wire n_210;
wire n_216;
wire n_83;
wire n_206;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_168;
wire n_153;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_227;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_189;
wire n_85;
wire n_99;
wire n_130;
wire n_84;
wire n_213;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_142;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_155;
wire n_219;
wire n_109;
wire n_150;
wire n_233;
wire n_122;
wire n_205;
wire n_140;
wire n_218;
wire n_234;
wire n_120;
wire n_251;
wire n_214;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_112;
wire n_172;
wire n_237;
wire n_81;
wire n_244;
wire n_181;
wire n_182;
wire n_124;
wire n_238;
wire n_239;
wire n_126;
wire n_243;
wire n_202;
wire n_94;
wire n_108;
wire n_97;
wire n_116;
wire n_211;
wire n_220;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_230;
wire n_93;
wire n_80;
wire n_141;
wire n_240;
wire n_135;
wire n_196;
wire n_200;
wire n_165;
wire n_139;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_248;
wire n_107;
wire n_229;
wire n_253;
wire n_190;
wire n_123;
wire n_136;
wire n_187;
wire n_89;
wire n_249;
wire n_173;
wire n_201;
wire n_250;
wire n_103;
wire n_111;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_232;
wire n_115;
wire n_128;
wire n_241;
wire n_79;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_221;

BUFx10_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_12),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_40),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_29),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_31),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_41),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_16),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_37),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_22),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_20),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_34),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_9),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_33),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_53),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_5),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_76),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_6),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_23),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_51),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_39),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_38),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_17),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_0),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_1),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_2),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_4),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_7),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_8),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_10),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_11),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_11),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_13),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_14),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_15),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_R g143 ( 
.A(n_112),
.B(n_17),
.Y(n_143)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_18),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_19),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_19),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

OR2x6_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_110),
.B1(n_91),
.B2(n_86),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_113),
.B1(n_116),
.B2(n_115),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_120),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_151),
.B1(n_129),
.B2(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_92),
.B1(n_93),
.B2(n_89),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_99),
.B1(n_101),
.B2(n_97),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_137),
.Y(n_162)
);

OR2x6_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_21),
.Y(n_163)
);

AO22x2_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_164)
);

AO22x2_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_109),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_119),
.B1(n_118),
.B2(n_117),
.Y(n_168)
);

BUFx6f_ASAP7_75t_SL g169 ( 
.A(n_132),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AO22x2_ASAP7_75t_L g171 ( 
.A1(n_125),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_144),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_167),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_131),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

NAND2x1p5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_133),
.Y(n_178)
);

NAND2x1p5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_128),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_161),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_181),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_147),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_147),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_148),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_191),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_142),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_134),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_136),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_184),
.Y(n_211)
);

OR2x6_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_175),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_185),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_163),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_180),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_209),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_200),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_216),
.B1(n_213),
.B2(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_214),
.B1(n_212),
.B2(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_222),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_218),
.B1(n_220),
.B2(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_228),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

BUFx2_ASAP7_75t_SL g238 ( 
.A(n_237),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NOR4xp25_ASAP7_75t_SL g245 ( 
.A(n_244),
.B(n_47),
.C(n_48),
.D(n_49),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_245),
.B1(n_55),
.B2(n_58),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_253)
);

AOI211xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_72),
.B(n_73),
.C(n_75),
.Y(n_254)
);


endmodule