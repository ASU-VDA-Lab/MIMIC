module fake_jpeg_30361_n_458 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_458);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_458;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_15),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_57),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_14),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_60),
.Y(n_100)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_68),
.Y(n_105)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_71),
.Y(n_106)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_13),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_13),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_42),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_32),
.B(n_0),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_18),
.C(n_34),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_89),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_31),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_33),
.B1(n_42),
.B2(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_95),
.B1(n_98),
.B2(n_104),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_43),
.B1(n_45),
.B2(n_42),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_94),
.A2(n_97),
.B1(n_113),
.B2(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_44),
.B1(n_35),
.B2(n_28),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_47),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_28),
.B1(n_35),
.B2(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_54),
.A2(n_29),
.B1(n_23),
.B2(n_37),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_108),
.A2(n_123),
.B1(n_139),
.B2(n_24),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_115),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_46),
.A2(n_41),
.B1(n_28),
.B2(n_35),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_41),
.B1(n_38),
.B2(n_27),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_131),
.B1(n_134),
.B2(n_41),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_12),
.B(n_10),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_34),
.B(n_18),
.C(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_135),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_77),
.B1(n_71),
.B2(n_64),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_41),
.B1(n_22),
.B2(n_27),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_63),
.A2(n_41),
.B1(n_26),
.B2(n_22),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_31),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_85),
.A2(n_78),
.B1(n_87),
.B2(n_81),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_26),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_142),
.B(n_143),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_58),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_155),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_162),
.Y(n_207)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g227 ( 
.A(n_146),
.Y(n_227)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_99),
.A2(n_52),
.B1(n_34),
.B2(n_18),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_170),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_156),
.B(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_65),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_160),
.A2(n_182),
.B1(n_138),
.B2(n_120),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_58),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_76),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_100),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_111),
.B(n_66),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_174),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_8),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_101),
.A2(n_17),
.B1(n_16),
.B2(n_78),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_179),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_141),
.A2(n_88),
.B1(n_17),
.B2(n_9),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_183),
.A2(n_98),
.B1(n_123),
.B2(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_119),
.B(n_9),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_185),
.C(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_95),
.B(n_9),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_109),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_17),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_92),
.B(n_1),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_16),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_121),
.C(n_92),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_191),
.C(n_215),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_92),
.C(n_101),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_92),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_196),
.A2(n_202),
.B(n_224),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_124),
.B1(n_96),
.B2(n_132),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_204),
.B1(n_228),
.B2(n_170),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_152),
.B1(n_165),
.B2(n_150),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_124),
.B1(n_102),
.B2(n_96),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_212),
.B1(n_217),
.B2(n_225),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_101),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_132),
.B1(n_102),
.B2(n_136),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_214),
.B(n_156),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_141),
.C(n_107),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_149),
.A2(n_129),
.B1(n_136),
.B2(n_110),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_162),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_171),
.A2(n_110),
.B1(n_122),
.B2(n_130),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_129),
.B1(n_122),
.B2(n_114),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_138),
.C(n_120),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_172),
.C(n_188),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_163),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_231),
.B(n_191),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_184),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_186),
.B1(n_175),
.B2(n_158),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_234),
.A2(n_247),
.B1(n_208),
.B2(n_221),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_235),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_237),
.B(n_242),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_164),
.B(n_185),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_214),
.B(n_208),
.Y(n_272)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_245),
.B1(n_248),
.B2(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_243),
.B(n_244),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

AO22x1_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_173),
.B1(n_166),
.B2(n_188),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_216),
.A2(n_144),
.B1(n_167),
.B2(n_173),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_155),
.B1(n_174),
.B2(n_173),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_197),
.A2(n_173),
.B1(n_168),
.B2(n_142),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_179),
.B1(n_159),
.B2(n_176),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_265),
.B1(n_225),
.B2(n_227),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_252),
.B(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_151),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_213),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_211),
.B(n_146),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_192),
.B(n_169),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_211),
.B(n_146),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_192),
.B(n_223),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_264),
.B(n_267),
.C(n_226),
.D(n_210),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_190),
.B(n_148),
.C(n_176),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_268),
.C(n_230),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_148),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_209),
.A2(n_159),
.B1(n_179),
.B2(n_130),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_189),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_125),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_190),
.B(n_126),
.C(n_125),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_275),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_210),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_260),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_276),
.A2(n_296),
.B1(n_247),
.B2(n_267),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_215),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_280),
.C(n_287),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_279),
.A2(n_286),
.B1(n_290),
.B2(n_301),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_191),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_202),
.A3(n_196),
.B1(n_213),
.B2(n_210),
.C1(n_205),
.C2(n_221),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_231),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_233),
.A2(n_234),
.B1(n_244),
.B2(n_252),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_230),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_294),
.C(n_237),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_199),
.B1(n_196),
.B2(n_216),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_220),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_202),
.C(n_220),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_242),
.A2(n_198),
.B(n_224),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_200),
.B1(n_217),
.B2(n_212),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_226),
.Y(n_298)
);

BUFx24_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_303),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_233),
.A2(n_201),
.B1(n_194),
.B2(n_229),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_232),
.A2(n_193),
.B(n_126),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_309),
.Y(n_339)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_307),
.A2(n_295),
.A3(n_272),
.B1(n_300),
.B2(n_294),
.C1(n_292),
.C2(n_273),
.Y(n_341)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_301),
.B1(n_283),
.B2(n_276),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_245),
.B1(n_265),
.B2(n_248),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_312),
.A2(n_330),
.B1(n_296),
.B2(n_273),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_261),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_322),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_321),
.C(n_328),
.Y(n_349)
);

XOR2x2_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_258),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_246),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_278),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_268),
.C(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_288),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_326),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_292),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_256),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_235),
.C(n_238),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_299),
.B(n_193),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_246),
.B1(n_241),
.B2(n_255),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_246),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_270),
.C(n_284),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_270),
.B(n_239),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_334),
.Y(n_346)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_323),
.B(n_325),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_336),
.A2(n_329),
.B(n_309),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_334),
.B(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_351),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_360),
.B1(n_331),
.B2(n_194),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_342),
.C(n_345),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_289),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_347),
.A2(n_358),
.B1(n_312),
.B2(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_274),
.Y(n_350)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_353),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_274),
.Y(n_355)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_355),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_274),
.C(n_269),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_357),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_120),
.C(n_138),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_311),
.A2(n_299),
.B1(n_194),
.B2(n_193),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_321),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_359),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_299),
.Y(n_360)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_361),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_353),
.B1(n_348),
.B2(n_342),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_336),
.A2(n_304),
.B(n_323),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_363),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_363),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_355),
.A2(n_319),
.B(n_330),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_350),
.A2(n_313),
.B(n_317),
.Y(n_368)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_337),
.B(n_316),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_374),
.B(n_380),
.Y(n_396)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_376),
.Y(n_387)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

AO221x1_ASAP7_75t_L g377 ( 
.A1(n_339),
.A2(n_333),
.B1(n_322),
.B2(n_313),
.C(n_195),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_381),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_379),
.A2(n_352),
.B1(n_361),
.B2(n_335),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_SL g380 ( 
.A(n_344),
.B(n_151),
.C(n_195),
.Y(n_380)
);

AO22x1_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_195),
.B1(n_2),
.B2(n_3),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_384),
.A2(n_375),
.B1(n_373),
.B2(n_376),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_338),
.A3(n_354),
.B1(n_340),
.B2(n_339),
.C1(n_348),
.C2(n_358),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_372),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_392),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_349),
.C(n_345),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_394),
.C(n_395),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_349),
.C(n_356),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_360),
.C(n_357),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_398),
.A2(n_371),
.B1(n_362),
.B2(n_384),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_335),
.C(n_16),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_402),
.C(n_365),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_400),
.B(n_366),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_379),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_381),
.B1(n_371),
.B2(n_364),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_16),
.C(n_17),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_390),
.B(n_383),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_405),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_409),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_408),
.A2(n_417),
.B1(n_377),
.B2(n_401),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_385),
.A2(n_364),
.B(n_369),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_1),
.Y(n_429)
);

NAND4xp25_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_389),
.C(n_380),
.D(n_396),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_412),
.Y(n_426)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_396),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_1),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_385),
.A2(n_369),
.B1(n_374),
.B2(n_367),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_414),
.A2(n_391),
.B1(n_397),
.B2(n_393),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_388),
.A2(n_383),
.B(n_380),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_1),
.B(n_2),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_367),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_416),
.B(n_370),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_370),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_419),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_394),
.C(n_395),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_422),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_407),
.B(n_402),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_406),
.A2(n_393),
.B1(n_397),
.B2(n_387),
.Y(n_424)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_405),
.A2(n_387),
.B1(n_400),
.B2(n_398),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_427),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_415),
.B(n_411),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_430),
.A2(n_409),
.B(n_412),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_431),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_437),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

BUFx24_ASAP7_75t_SL g438 ( 
.A(n_426),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_439),
.Y(n_447)
);

AO221x1_ASAP7_75t_L g439 ( 
.A1(n_420),
.A2(n_414),
.B1(n_404),
.B2(n_410),
.C(n_6),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_430),
.A2(n_404),
.B(n_4),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g445 ( 
.A1(n_441),
.A2(n_419),
.B(n_424),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_425),
.C(n_423),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_442),
.A2(n_449),
.B(n_445),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_423),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_443),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_446),
.Y(n_453)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_440),
.A2(n_429),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_2),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_436),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_437),
.B1(n_433),
.B2(n_7),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_450),
.A2(n_452),
.B(n_443),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_SL g451 ( 
.A(n_444),
.B(n_4),
.C(n_5),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_442),
.C(n_447),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_455),
.A2(n_456),
.B(n_454),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_457),
.B(n_453),
.Y(n_458)
);


endmodule