module fake_jpeg_12101_n_62 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_22),
.C(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_3),
.Y(n_34)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_34),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_25),
.B1(n_23),
.B2(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_13),
.C(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.C(n_47),
.Y(n_54)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_4),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_38),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_23),
.B1(n_8),
.B2(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NOR4xp25_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_55),
.C(n_57),
.D(n_49),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_54),
.B(n_56),
.C(n_21),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_17),
.C(n_20),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);


endmodule