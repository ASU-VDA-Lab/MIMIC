module real_jpeg_2379_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_288;
wire n_286;
wire n_83;
wire n_166;
wire n_176;
wire n_292;
wire n_249;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_283;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_39),
.B1(n_69),
.B2(n_71),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_3),
.A2(n_50),
.B1(n_69),
.B2(n_71),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_3),
.B(n_29),
.C(n_33),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_31),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_3),
.B(n_56),
.C(n_60),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_3),
.B(n_95),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_67),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_68),
.C(n_71),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_62),
.Y(n_234)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_6),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_6),
.A2(n_48),
.B1(n_69),
.B2(n_71),
.Y(n_159)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_9),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_11),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_11),
.A2(n_25),
.B1(n_59),
.B2(n_60),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_25),
.B1(n_69),
.B2(n_71),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_292),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_12),
.B(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_41),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_40),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_20),
.A2(n_27),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_26),
.B(n_49),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_31),
.B1(n_46),
.B2(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_49),
.Y(n_79)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_33),
.B(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_38),
.B(n_79),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_36),
.A2(n_47),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_37),
.B(n_43),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_80),
.B(n_291),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_76),
.C(n_78),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_44),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.C(n_64),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_45),
.A2(n_106),
.B1(n_143),
.B2(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_45),
.B(n_143),
.C(n_153),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_45),
.A2(n_106),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_51),
.A2(n_64),
.B1(n_265),
.B2(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_51),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_51)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_53),
.A2(n_62),
.B1(n_102),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_58),
.B(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

AOI22x1_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_58),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_72),
.Y(n_74)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_60),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_64),
.A2(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_64),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_64),
.B(n_128),
.C(n_266),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_73),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_66),
.A2(n_73),
.B1(n_90),
.B2(n_91),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_66),
.A2(n_73),
.B(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_67),
.A2(n_75),
.B1(n_116),
.B2(n_142),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_71),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_76),
.B(n_78),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_286),
.B(n_290),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_257),
.B(n_283),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_147),
.B(n_256),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_129),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_84),
.B(n_129),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_107),
.C(n_118),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_85),
.B(n_107),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_101),
.C(n_106),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_88),
.A2(n_89),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_88),
.A2(n_89),
.B1(n_207),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_89),
.B(n_202),
.C(n_207),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_89),
.B(n_158),
.C(n_234),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_94),
.A2(n_95),
.B1(n_123),
.B2(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_97),
.B(n_122),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_97),
.A2(n_122),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_127),
.C(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_101),
.A2(n_105),
.B1(n_169),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_101),
.A2(n_105),
.B1(n_124),
.B2(n_125),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_101),
.B(n_124),
.C(n_242),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_103),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_117),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_110),
.B(n_123),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_117),
.A2(n_133),
.B(n_138),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_118),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.C(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_119),
.A2(n_120),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_124),
.A2(n_125),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_124),
.B(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_128),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_127),
.A2(n_128),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_127),
.A2(n_128),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_128),
.B(n_277),
.C(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_146),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_139),
.B2(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_132),
.B(n_139),
.C(n_146),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B(n_145),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_143),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_177),
.C(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_143),
.A2(n_161),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_145),
.A2(n_261),
.B1(n_262),
.B2(n_270),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_145),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_251),
.B(n_255),
.Y(n_147)
);

OAI211xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_180),
.B(n_194),
.C(n_195),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_170),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_162),
.B2(n_163),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_165),
.C(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_157),
.A2(n_158),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_158),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_158),
.B(n_222),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_176),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_176),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_178),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_196),
.C(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_186),
.C(n_192),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_213),
.B(n_250),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_201),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_244),
.B(n_249),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_238),
.B(n_243),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_230),
.B(n_237),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_229),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B(n_223),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_236),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_273),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_272),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_272),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_270),
.C(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_282),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);


endmodule