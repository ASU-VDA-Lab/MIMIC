module fake_jpeg_29913_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_65),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_51),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_55),
.B1(n_47),
.B2(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_92),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_49),
.B(n_53),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_4),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_97),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_104),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_50),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_45),
.C(n_23),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_22),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_110),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_81),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_116),
.B1(n_6),
.B2(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_27),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_32),
.B(n_5),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_13),
.B(n_15),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_11),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_125),
.B(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_109),
.B1(n_106),
.B2(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_130),
.B(n_131),
.Y(n_136)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_18),
.B(n_20),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_99),
.C(n_29),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_137),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_126),
.C(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_129),
.B1(n_119),
.B2(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_134),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_143),
.C(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_24),
.Y(n_148)
);


endmodule