module real_aes_6569_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_310;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_0), .A2(n_32), .B1(n_356), .B2(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_1), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_2), .A2(n_217), .B1(n_380), .B2(n_487), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_3), .A2(n_674), .B1(n_698), .B2(n_699), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_3), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_4), .A2(n_24), .B1(n_360), .B2(n_362), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_5), .B(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_6), .A2(n_101), .B1(n_356), .B2(n_484), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_7), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_8), .A2(n_172), .B1(n_450), .B2(n_452), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_9), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_10), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_11), .A2(n_120), .B1(n_304), .B2(n_311), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_12), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_13), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_14), .A2(n_21), .B1(n_323), .B2(n_546), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_15), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_16), .A2(n_171), .B1(n_383), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_17), .A2(n_36), .B1(n_496), .B2(n_497), .Y(n_495) );
AO22x2_ASAP7_75t_L g257 ( .A1(n_18), .A2(n_65), .B1(n_249), .B2(n_254), .Y(n_257) );
INVx1_ASAP7_75t_L g670 ( .A(n_18), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_19), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_20), .A2(n_57), .B1(n_455), .B2(n_496), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_22), .B(n_549), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_23), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_25), .A2(n_211), .B1(n_362), .B2(n_458), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_26), .A2(n_156), .B1(n_375), .B2(n_377), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_27), .A2(n_126), .B1(n_448), .B2(n_594), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_28), .A2(n_185), .B1(n_448), .B2(n_653), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_29), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_30), .A2(n_158), .B1(n_352), .B2(n_353), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_31), .Y(n_639) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_33), .A2(n_70), .B1(n_249), .B2(n_250), .Y(n_259) );
INVx1_ASAP7_75t_L g671 ( .A(n_33), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_34), .A2(n_78), .B1(n_356), .B2(n_357), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_35), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_37), .A2(n_199), .B1(n_357), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_38), .A2(n_159), .B1(n_383), .B2(n_482), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_39), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_40), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_41), .A2(n_190), .B1(n_360), .B2(n_373), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_42), .A2(n_170), .B1(n_585), .B2(n_596), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_43), .A2(n_62), .B1(n_281), .B2(n_383), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_44), .A2(n_72), .B1(n_511), .B2(n_512), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_45), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_46), .A2(n_127), .B1(n_317), .B2(n_475), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_47), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_48), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_49), .A2(n_60), .B1(n_340), .B2(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_50), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_51), .A2(n_110), .B1(n_476), .B2(n_546), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_52), .Y(n_284) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_53), .A2(n_130), .B1(n_349), .B2(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_54), .B(n_405), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_55), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_56), .A2(n_74), .B1(n_380), .B2(n_381), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_58), .A2(n_64), .B1(n_383), .B2(n_455), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_59), .A2(n_153), .B1(n_482), .B2(n_484), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_61), .A2(n_122), .B1(n_504), .B2(n_507), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_63), .A2(n_124), .B1(n_319), .B2(n_323), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_66), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_67), .A2(n_69), .B1(n_103), .B2(n_300), .C1(n_323), .C2(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_68), .A2(n_128), .B1(n_287), .B2(n_501), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_71), .A2(n_207), .B1(n_306), .B2(n_349), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_73), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_75), .Y(n_720) );
AND2x2_ASAP7_75t_L g229 ( .A(n_76), .B(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_77), .A2(n_157), .B1(n_265), .B2(n_272), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_79), .A2(n_203), .B1(n_352), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_80), .A2(n_133), .B1(n_383), .B2(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_81), .A2(n_219), .B1(n_499), .B2(n_558), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_82), .Y(n_366) );
INVx1_ASAP7_75t_L g226 ( .A(n_83), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_84), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_85), .A2(n_108), .B1(n_313), .B2(n_349), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_86), .A2(n_95), .B1(n_357), .B2(n_638), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_87), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_88), .A2(n_154), .B1(n_243), .B2(n_260), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_89), .A2(n_191), .B1(n_327), .B2(n_330), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_90), .A2(n_214), .B1(n_313), .B2(n_341), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_91), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_92), .A2(n_186), .B1(n_561), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_93), .A2(n_96), .B1(n_341), .B2(n_553), .Y(n_552) );
OA22x2_ASAP7_75t_L g536 ( .A1(n_94), .A2(n_537), .B1(n_538), .B2(n_564), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_94), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_97), .B(n_312), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_98), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_99), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_100), .B(n_347), .Y(n_551) );
OA22x2_ASAP7_75t_L g565 ( .A1(n_102), .A2(n_566), .B1(n_567), .B2(n_588), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_102), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_104), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_105), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_106), .A2(n_111), .B1(n_327), .B2(n_330), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_107), .A2(n_134), .B1(n_360), .B2(n_509), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_109), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_112), .B(n_344), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_113), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_114), .Y(n_601) );
XNOR2x2_ASAP7_75t_L g238 ( .A(n_115), .B(n_239), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_116), .A2(n_137), .B1(n_645), .B2(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g230 ( .A(n_117), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_118), .A2(n_143), .B1(n_265), .B2(n_385), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_119), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_121), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_123), .B(n_549), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_125), .Y(n_529) );
INVx1_ASAP7_75t_L g707 ( .A(n_129), .Y(n_707) );
OA22x2_ASAP7_75t_L g710 ( .A1(n_129), .A2(n_707), .B1(n_711), .B2(n_731), .Y(n_710) );
AND2x6_ASAP7_75t_L g225 ( .A(n_131), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_131), .Y(n_664) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_132), .A2(n_180), .B1(n_249), .B2(n_250), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_135), .A2(n_152), .B1(n_455), .B2(n_456), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_136), .A2(n_166), .B1(n_695), .B2(n_696), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_138), .A2(n_223), .B(n_231), .C(n_672), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g316 ( .A1(n_139), .A2(n_187), .B1(n_317), .B2(n_321), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_140), .A2(n_201), .B1(n_482), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_141), .A2(n_169), .B1(n_402), .B2(n_458), .Y(n_582) );
INVx1_ASAP7_75t_L g459 ( .A(n_142), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_144), .A2(n_189), .B1(n_385), .B2(n_636), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_145), .A2(n_208), .B1(n_287), .B2(n_484), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_146), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_147), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_148), .B(n_321), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_149), .A2(n_196), .B1(n_561), .B2(n_562), .Y(n_560) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_150), .A2(n_193), .B1(n_249), .B2(n_254), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_151), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_155), .A2(n_173), .B1(n_484), .B2(n_653), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_160), .A2(n_182), .B1(n_266), .B2(n_558), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_161), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_162), .A2(n_168), .B1(n_265), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_163), .A2(n_188), .B1(n_260), .B2(n_365), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_164), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_165), .A2(n_195), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_167), .A2(n_369), .B1(n_416), .B2(n_417), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_167), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_174), .A2(n_200), .B1(n_365), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_175), .A2(n_205), .B1(n_340), .B2(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_176), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_177), .B(n_311), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_178), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_179), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_180), .B(n_669), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_181), .Y(n_527) );
INVx1_ASAP7_75t_L g590 ( .A(n_183), .Y(n_590) );
INVx1_ASAP7_75t_L g490 ( .A(n_184), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_192), .A2(n_212), .B1(n_383), .B2(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g667 ( .A(n_193), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_194), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_197), .A2(n_202), .B1(n_356), .B2(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_198), .Y(n_515) );
XNOR2x2_ASAP7_75t_L g641 ( .A(n_204), .B(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_206), .A2(n_492), .B1(n_531), .B2(n_532), .Y(n_491) );
INVx1_ASAP7_75t_L g531 ( .A(n_206), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_209), .Y(n_682) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_213), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_215), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_216), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_218), .A2(n_221), .B1(n_499), .B2(n_501), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_220), .Y(n_473) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_226), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_227), .A2(n_662), .B(n_706), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_419), .B1(n_657), .B2(n_658), .C(n_659), .Y(n_231) );
INVx1_ASAP7_75t_L g658 ( .A(n_232), .Y(n_658) );
AOI22xp5_ASAP7_75t_SL g232 ( .A1(n_233), .A2(n_234), .B1(n_367), .B2(n_418), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B1(n_332), .B2(n_333), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_240), .B(n_297), .Y(n_239) );
NOR3xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_276), .C(n_289), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_264), .Y(n_241) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx3_ASAP7_75t_L g373 ( .A(n_244), .Y(n_373) );
BUFx3_ASAP7_75t_L g496 ( .A(n_244), .Y(n_496) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx2_ASAP7_75t_SL g365 ( .A(n_245), .Y(n_365) );
INVx2_ASAP7_75t_L g483 ( .A(n_245), .Y(n_483) );
BUFx2_ASAP7_75t_SL g653 ( .A(n_245), .Y(n_653) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
AND2x6_ASAP7_75t_L g281 ( .A(n_246), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g292 ( .A(n_246), .B(n_271), .Y(n_292) );
AND2x6_ASAP7_75t_L g300 ( .A(n_246), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
AND2x2_ASAP7_75t_L g288 ( .A(n_247), .B(n_253), .Y(n_288) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_248), .B(n_253), .Y(n_263) );
AND2x2_ASAP7_75t_L g269 ( .A(n_248), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g310 ( .A(n_248), .B(n_257), .Y(n_310) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g254 ( .A(n_251), .Y(n_254) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g270 ( .A(n_253), .Y(n_270) );
INVx1_ASAP7_75t_L g309 ( .A(n_253), .Y(n_309) );
AND2x4_ASAP7_75t_L g261 ( .A(n_255), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g287 ( .A(n_255), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_255), .B(n_269), .Y(n_296) );
AND2x2_ASAP7_75t_L g363 ( .A(n_255), .B(n_269), .Y(n_363) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
AND2x2_ASAP7_75t_L g271 ( .A(n_256), .B(n_259), .Y(n_271) );
OR2x2_ASAP7_75t_L g283 ( .A(n_256), .B(n_259), .Y(n_283) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g301 ( .A(n_257), .B(n_259), .Y(n_301) );
AND2x2_ASAP7_75t_L g308 ( .A(n_258), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g392 ( .A(n_258), .Y(n_392) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
BUFx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g377 ( .A(n_261), .Y(n_377) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_261), .Y(n_448) );
BUFx2_ASAP7_75t_L g484 ( .A(n_261), .Y(n_484) );
BUFx3_ASAP7_75t_L g587 ( .A(n_261), .Y(n_587) );
AND2x2_ASAP7_75t_L g596 ( .A(n_262), .B(n_392), .Y(n_596) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x6_ASAP7_75t_L g274 ( .A(n_263), .B(n_275), .Y(n_274) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g451 ( .A(n_266), .Y(n_451) );
INVx4_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g354 ( .A(n_267), .Y(n_354) );
INVx3_ASAP7_75t_L g487 ( .A(n_267), .Y(n_487) );
INVx2_ASAP7_75t_L g511 ( .A(n_267), .Y(n_511) );
INVx5_ASAP7_75t_L g585 ( .A(n_267), .Y(n_585) );
INVx1_ASAP7_75t_L g729 ( .A(n_267), .Y(n_729) );
INVx8_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g325 ( .A(n_270), .Y(n_325) );
AND2x6_ASAP7_75t_L g331 ( .A(n_271), .B(n_288), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_271), .B(n_288), .Y(n_415) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g357 ( .A(n_273), .Y(n_357) );
BUFx4f_ASAP7_75t_SL g385 ( .A(n_273), .Y(n_385) );
BUFx2_ASAP7_75t_L g489 ( .A(n_273), .Y(n_489) );
BUFx2_ASAP7_75t_L g512 ( .A(n_273), .Y(n_512) );
INVx6_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g452 ( .A(n_274), .Y(n_452) );
INVx1_ASAP7_75t_SL g558 ( .A(n_274), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_274), .A2(n_396), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g320 ( .A(n_275), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B1(n_284), .B2(n_285), .Y(n_276) );
INVx2_ASAP7_75t_L g497 ( .A(n_278), .Y(n_497) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx5_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx4_ASAP7_75t_L g725 ( .A(n_280), .Y(n_725) );
INVx11_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx11_ASAP7_75t_L g361 ( .A(n_281), .Y(n_361) );
AND2x4_ASAP7_75t_L g329 ( .A(n_282), .B(n_288), .Y(n_329) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g410 ( .A(n_283), .B(n_411), .Y(n_410) );
INVx4_ASAP7_75t_L g456 ( .A(n_285), .Y(n_456) );
INVx4_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g356 ( .A(n_287), .Y(n_356) );
BUFx3_ASAP7_75t_L g376 ( .A(n_287), .Y(n_376) );
INVx2_ASAP7_75t_L g500 ( .A(n_287), .Y(n_500) );
BUFx3_ASAP7_75t_L g638 ( .A(n_287), .Y(n_638) );
INVx1_ASAP7_75t_L g411 ( .A(n_288), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_293), .B2(n_294), .Y(n_289) );
INVx2_ASAP7_75t_L g352 ( .A(n_291), .Y(n_352) );
INVx2_ASAP7_75t_L g380 ( .A(n_291), .Y(n_380) );
INVx3_ASAP7_75t_L g562 ( .A(n_291), .Y(n_562) );
INVx2_ASAP7_75t_L g645 ( .A(n_291), .Y(n_645) );
INVx6_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g458 ( .A(n_292), .Y(n_458) );
BUFx3_ASAP7_75t_L g506 ( .A(n_292), .Y(n_506) );
BUFx3_ASAP7_75t_L g695 ( .A(n_292), .Y(n_695) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_315), .Y(n_297) );
OAI21xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_302), .B(n_303), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
INVx4_ASAP7_75t_L g438 ( .A(n_300), .Y(n_438) );
BUFx3_ASAP7_75t_L g542 ( .A(n_300), .Y(n_542) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_300), .Y(n_581) );
AND2x4_ASAP7_75t_L g324 ( .A(n_301), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g397 ( .A(n_301), .Y(n_397) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g440 ( .A(n_306), .Y(n_440) );
INVx2_ASAP7_75t_L g523 ( .A(n_306), .Y(n_523) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g402 ( .A(n_307), .Y(n_402) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_307), .Y(n_476) );
BUFx4f_ASAP7_75t_SL g545 ( .A(n_307), .Y(n_545) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_307), .Y(n_718) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g314 ( .A(n_309), .Y(n_314) );
AND2x4_ASAP7_75t_L g313 ( .A(n_310), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g319 ( .A(n_310), .B(n_320), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_310), .B(n_392), .Y(n_391) );
BUFx4f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g618 ( .A(n_312), .Y(n_618) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
BUFx12f_ASAP7_75t_L g546 ( .A(n_313), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_326), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
BUFx3_ASAP7_75t_L g553 ( .A(n_319), .Y(n_553) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_SL g341 ( .A(n_324), .Y(n_341) );
INVx1_ASAP7_75t_L g398 ( .A(n_325), .Y(n_398) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx5_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
INVx2_ASAP7_75t_L g716 ( .A(n_328), .Y(n_716) );
INVx4_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g344 ( .A(n_331), .Y(n_344) );
INVx1_ASAP7_75t_SL g550 ( .A(n_331), .Y(n_550) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
XOR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_366), .Y(n_333) );
NAND3x1_ASAP7_75t_L g334 ( .A(n_335), .B(n_350), .C(n_358), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_342), .Y(n_335) );
OAI21xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_338), .B(n_339), .Y(n_336) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_337), .A2(n_400), .B1(n_401), .B2(n_403), .C(n_404), .Y(n_399) );
BUFx3_ASAP7_75t_L g405 ( .A(n_340), .Y(n_405) );
INVx2_ASAP7_75t_L g656 ( .A(n_340), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .C(n_348), .Y(n_342) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_364), .Y(n_358) );
INVx4_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g455 ( .A(n_361), .Y(n_455) );
INVx4_ASAP7_75t_L g561 ( .A(n_361), .Y(n_561) );
OAI21xp33_ASAP7_75t_SL g572 ( .A1(n_361), .A2(n_573), .B(n_574), .Y(n_572) );
BUFx3_ASAP7_75t_L g696 ( .A(n_362), .Y(n_696) );
BUFx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g383 ( .A(n_363), .Y(n_383) );
BUFx3_ASAP7_75t_L g509 ( .A(n_363), .Y(n_509) );
INVx1_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g417 ( .A(n_369), .Y(n_417) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_370), .B(n_386), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_378), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g501 ( .A(n_377), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR3xp33_ASAP7_75t_SL g386 ( .A(n_387), .B(n_399), .C(n_406), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_393), .B2(n_394), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_389), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_441) );
INVx3_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_391), .A2(n_473), .B1(n_474), .B2(n_477), .Y(n_472) );
BUFx3_ASAP7_75t_L g528 ( .A(n_391), .Y(n_528) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g444 ( .A(n_395), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g530 ( .A(n_396), .Y(n_530) );
OR2x6_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_412), .B2(n_413), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_408), .A2(n_431), .B1(n_432), .B2(n_433), .Y(n_430) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g678 ( .A(n_409), .Y(n_678) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g465 ( .A(n_410), .Y(n_465) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_410), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_410), .A2(n_414), .B1(n_601), .B2(n_602), .C(n_603), .Y(n_600) );
BUFx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
INVxp67_ASAP7_75t_L g657 ( .A(n_419), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_609), .B2(n_610), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
XNOR2xp5_ASAP7_75t_SL g421 ( .A(n_422), .B(n_534), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_491), .B2(n_533), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
XNOR2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_460), .Y(n_426) );
XOR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_459), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_445), .Y(n_428) );
NOR3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_435), .C(n_441), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_433), .A2(n_622), .B1(n_623), .B2(n_625), .Y(n_621) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_439), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g719 ( .A1(n_437), .A2(n_720), .B(n_721), .Y(n_719) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g469 ( .A1(n_438), .A2(n_470), .B(n_471), .Y(n_469) );
INVx4_ASAP7_75t_L g521 ( .A(n_438), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_453), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_457), .Y(n_453) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_490), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_478), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_469), .C(n_472), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_465), .A2(n_518), .B1(n_570), .B2(n_571), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_467), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g518 ( .A(n_468), .Y(n_518) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g628 ( .A(n_476), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_485), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g594 ( .A(n_483), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g533 ( .A(n_491), .Y(n_533) );
INVx2_ASAP7_75t_L g532 ( .A(n_492), .Y(n_532) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_493), .B(n_513), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .C(n_526), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_514) );
INVx1_ASAP7_75t_L g624 ( .A(n_516), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_523), .B2(n_524), .C(n_525), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_529), .B2(n_530), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_528), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_528), .A2(n_530), .B1(n_687), .B2(n_688), .Y(n_686) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_589), .B1(n_607), .B2(n_608), .Y(n_534) );
INVx1_ASAP7_75t_L g607 ( .A(n_535), .Y(n_607) );
XOR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_565), .Y(n_535) );
INVx1_ASAP7_75t_L g564 ( .A(n_538), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_554), .Y(n_538) );
NOR2xp67_ASAP7_75t_L g539 ( .A(n_540), .B(n_547), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_543), .B(n_544), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_541), .A2(n_605), .B(n_606), .Y(n_604) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g683 ( .A(n_545), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .C(n_552), .Y(n_547) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_578), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .C(n_575), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_583), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx2_ASAP7_75t_L g616 ( .A(n_581), .Y(n_616) );
INVx2_ASAP7_75t_SL g681 ( .A(n_581), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_585), .Y(n_636) );
INVx2_ASAP7_75t_SL g608 ( .A(n_589), .Y(n_608) );
XNOR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NOR4xp75_ASAP7_75t_L g591 ( .A(n_592), .B(n_597), .C(n_600), .D(n_604), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_593), .B(n_595), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_599), .Y(n_597) );
CKINVDCx16_ASAP7_75t_R g609 ( .A(n_610), .Y(n_609) );
OAI22xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_612), .B1(n_640), .B2(n_641), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
XOR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_639), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_630), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_621), .C(n_626), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_619), .C(n_620), .Y(n_615) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND4xp75_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .C(n_650), .D(n_654), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
AND2x2_ASAP7_75t_SL g647 ( .A(n_648), .B(n_649), .Y(n_647) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_665), .Y(n_660) );
OR2x2_ASAP7_75t_SL g734 ( .A(n_661), .B(n_666), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_662), .Y(n_701) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_663), .B(n_703), .Y(n_706) );
CKINVDCx16_ASAP7_75t_R g703 ( .A(n_664), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OAI322xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_700), .A3(n_702), .B1(n_704), .B2(n_707), .C1(n_708), .C2(n_732), .Y(n_672) );
INVx2_ASAP7_75t_SL g699 ( .A(n_674), .Y(n_699) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_689), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_680), .C(n_686), .Y(n_675) );
OAI221xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B1(n_683), .B2(n_684), .C(n_685), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
CKINVDCx16_ASAP7_75t_R g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g731 ( .A(n_711), .Y(n_731) );
NAND2x1p5_ASAP7_75t_L g711 ( .A(n_712), .B(n_722), .Y(n_711) );
NOR2xp67_ASAP7_75t_SL g712 ( .A(n_713), .B(n_719), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .C(n_717), .Y(n_713) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
endmodule