module fake_jpeg_19726_n_142 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_17),
.B1(n_18),
.B2(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_17),
.B(n_18),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_34),
.B1(n_25),
.B2(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_31),
.B1(n_34),
.B2(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_46),
.B1(n_23),
.B2(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_12),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_23),
.B1(n_27),
.B2(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_57),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_61),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_45),
.B(n_42),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_35),
.B(n_43),
.C(n_42),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_22),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_42),
.C(n_35),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_22),
.C(n_32),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_57),
.B(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_47),
.B1(n_58),
.B2(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_77),
.B1(n_40),
.B2(n_26),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_51),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_82),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_16),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_67),
.C(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_26),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_92),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_60),
.B1(n_61),
.B2(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_62),
.B1(n_24),
.B2(n_14),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_59),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_55),
.C(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_18),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_21),
.B1(n_32),
.B2(n_15),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_77),
.C(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_99),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_21),
.B1(n_16),
.B2(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_102),
.B1(n_90),
.B2(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_83),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_94),
.C(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_112),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_103),
.B1(n_19),
.B2(n_13),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_83),
.C(n_13),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_116),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_103),
.B(n_4),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_13),
.C(n_10),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_10),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_117),
.Y(n_125)
);

OAI31xp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_5),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_3),
.B(n_4),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_111),
.B1(n_110),
.B2(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_128),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_5),
.B(n_6),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_133),
.C(n_6),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_19),
.B1(n_7),
.B2(n_9),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_126),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_7),
.B(n_9),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_135),
.B1(n_19),
.B2(n_9),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_10),
.Y(n_142)
);


endmodule