module fake_aes_9448_n_29 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
OA21x2_ASAP7_75t_L g14 ( .A1(n_4), .A2(n_3), .B(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
OR2x6_ASAP7_75t_L g19 ( .A(n_1), .B(n_10), .Y(n_19) );
AOI221xp5_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_0), .B1(n_2), .B2(n_5), .C(n_6), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
NOR2xp33_ASAP7_75t_SL g23 ( .A(n_22), .B(n_16), .Y(n_23) );
AOI211xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_20), .B(n_15), .C(n_19), .Y(n_24) );
XNOR2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_19), .Y(n_25) );
OAI31xp33_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_14), .A3(n_12), .B(n_13), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_27), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_25), .B1(n_14), .B2(n_11), .Y(n_29) );
endmodule