module fake_jpeg_24848_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_1),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_16),
.Y(n_23)
);

INVx5_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_18),
.B1(n_10),
.B2(n_8),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_7),
.B(n_6),
.C(n_12),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_3),
.B1(n_10),
.B2(n_6),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_10),
.B1(n_8),
.B2(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.C(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_19),
.C(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_17),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_18),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_30),
.B(n_33),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_32),
.C(n_22),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_34),
.Y(n_40)
);

NAND2x1p5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_15),
.Y(n_41)
);


endmodule