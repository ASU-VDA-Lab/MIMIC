module fake_jpeg_18064_n_33 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

OAI22x1_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_16),
.B1(n_2),
.B2(n_11),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_16),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

AOI31xp67_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_23),
.A3(n_13),
.B(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_26),
.B1(n_23),
.B2(n_9),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_33)
);


endmodule