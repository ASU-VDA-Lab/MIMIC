module fake_jpeg_9284_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_47),
.B1(n_18),
.B2(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_53),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_38),
.B1(n_43),
.B2(n_30),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_75),
.B1(n_89),
.B2(n_16),
.Y(n_106)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_41),
.B1(n_38),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_72),
.B1(n_85),
.B2(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_38),
.B1(n_39),
.B2(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_84),
.B1(n_26),
.B2(n_31),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_83),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_33),
.B1(n_18),
.B2(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_80),
.B1(n_82),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_39),
.B1(n_16),
.B2(n_24),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_18),
.B1(n_26),
.B2(n_31),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_42),
.B(n_80),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_63),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_68),
.A3(n_105),
.B1(n_113),
.B2(n_116),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_94),
.Y(n_123)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_29),
.B1(n_22),
.B2(n_19),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_99),
.B(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_116),
.B(n_22),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_88),
.B1(n_83),
.B2(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_35),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_77),
.B(n_67),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_45),
.B(n_62),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_127),
.B(n_97),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_143),
.B1(n_86),
.B2(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_67),
.B1(n_39),
.B2(n_49),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_118),
.B1(n_60),
.B2(n_86),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_76),
.B1(n_62),
.B2(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_140),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_21),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_65),
.B1(n_81),
.B2(n_49),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_65),
.B1(n_81),
.B2(n_49),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_35),
.CI(n_36),
.CON(n_136),
.SN(n_136)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_145),
.Y(n_149)
);

XOR2x2_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_106),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_36),
.CI(n_40),
.CON(n_165),
.SN(n_165)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_24),
.B1(n_57),
.B2(n_21),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_29),
.B(n_91),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_20),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_20),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_57),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_40),
.B(n_36),
.C(n_35),
.D(n_27),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_136),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_148),
.B(n_165),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_166),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_93),
.B1(n_117),
.B2(n_94),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_164),
.B1(n_171),
.B2(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_142),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_161),
.B(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_14),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_160),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_63),
.C(n_95),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.C(n_167),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_63),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2x1_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_35),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_112),
.B1(n_118),
.B2(n_57),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_63),
.C(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_11),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_126),
.A2(n_86),
.B1(n_27),
.B2(n_28),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_133),
.B(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_124),
.B(n_28),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_40),
.C(n_36),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_137),
.C(n_40),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_122),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_122),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_134),
.B1(n_135),
.B2(n_125),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_120),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_194),
.C(n_195),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_182),
.B1(n_191),
.B2(n_171),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_132),
.B1(n_129),
.B2(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_191),
.B1(n_193),
.B2(n_180),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_196),
.B(n_208),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_178),
.B1(n_162),
.B2(n_159),
.Y(n_191)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_147),
.B1(n_136),
.B2(n_140),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_137),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_27),
.B1(n_17),
.B2(n_36),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_40),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_203),
.C(n_177),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_40),
.A3(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_202),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_79),
.C(n_73),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_166),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_204),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_154),
.A2(n_149),
.B(n_170),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_152),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_212),
.B(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_209),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_179),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_214),
.B(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_165),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_217),
.B(n_227),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_151),
.B1(n_167),
.B2(n_162),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_220),
.B1(n_13),
.B2(n_12),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_151),
.B1(n_173),
.B2(n_176),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_165),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_225),
.C(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_196),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_172),
.B(n_155),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_79),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_199),
.Y(n_232)
);

CKINVDCx11_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_186),
.A2(n_193),
.B1(n_181),
.B2(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_0),
.C(n_1),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_203),
.C(n_200),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_193),
.B1(n_183),
.B2(n_189),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_246),
.B1(n_229),
.B2(n_212),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_210),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_224),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_217),
.Y(n_258)
);

FAx1_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_183),
.CI(n_195),
.CON(n_242),
.SN(n_242)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_240),
.C(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_216),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_0),
.C(n_2),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_250),
.C(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_224),
.C(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_235),
.B(n_245),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_226),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_243),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_253),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_264),
.C(n_268),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_213),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_223),
.C(n_219),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_247),
.B(n_222),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_2),
.C(n_3),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_3),
.C(n_4),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_3),
.C(n_4),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_4),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_237),
.B1(n_254),
.B2(n_236),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_275),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_237),
.B1(n_236),
.B2(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_281),
.C(n_271),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_281),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_248),
.B1(n_242),
.B2(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_242),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_283),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_268),
.B1(n_259),
.B2(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_296),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_292),
.B1(n_6),
.B2(n_7),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_9),
.B(n_12),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_295),
.B(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_300),
.Y(n_306)
);

AOI21x1_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_276),
.B(n_280),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_302),
.B1(n_287),
.B2(n_292),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_280),
.B1(n_7),
.B2(n_8),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_8),
.C(n_6),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_308),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_286),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_294),
.B(n_305),
.Y(n_314)
);

OR2x6_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_301),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_306),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_311),
.B(n_6),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_7),
.Y(n_320)
);


endmodule