module fake_jpeg_20879_n_257 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_6),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_24),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_48),
.B1(n_54),
.B2(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_33),
.Y(n_79)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_42),
.B1(n_30),
.B2(n_25),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_27),
.B1(n_31),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_42),
.B1(n_45),
.B2(n_63),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_31),
.B1(n_27),
.B2(n_40),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_42),
.B1(n_45),
.B2(n_31),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_27),
.C(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_32),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_54),
.B1(n_62),
.B2(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_91),
.B1(n_50),
.B2(n_70),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_55),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_89),
.Y(n_119)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_90),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_53),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_73),
.B(n_65),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_99),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_96),
.Y(n_102)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_60),
.B1(n_56),
.B2(n_52),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_66),
.B(n_68),
.C(n_52),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_80),
.B1(n_65),
.B2(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_82),
.B(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_59),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_75),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_114),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_117),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_50),
.B1(n_64),
.B2(n_56),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_18),
.B(n_15),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_90),
.B1(n_99),
.B2(n_88),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_125),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_133),
.B1(n_102),
.B2(n_105),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_96),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_28),
.B1(n_20),
.B2(n_13),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_59),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_140),
.Y(n_147)
);

CKINVDCx12_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

AO221x1_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_109),
.B1(n_116),
.B2(n_21),
.C(n_23),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_32),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_20),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_59),
.C(n_21),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_109),
.C(n_14),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_23),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_20),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_16),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_17),
.B1(n_13),
.B2(n_23),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_116),
.B(n_117),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_146),
.B(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_16),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_19),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_109),
.C(n_14),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_164),
.C(n_12),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_18),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_109),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_127),
.B1(n_123),
.B2(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_16),
.B1(n_18),
.B2(n_15),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_15),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_136),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_14),
.C(n_12),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_176),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_12),
.C(n_28),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_153),
.C(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_12),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_181),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_1),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_161),
.B1(n_163),
.B2(n_143),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_SL g187 ( 
.A(n_184),
.B(n_162),
.C(n_145),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_200),
.B(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_185),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_148),
.C(n_164),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_152),
.C(n_148),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_163),
.C(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_17),
.C(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_17),
.C(n_23),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_7),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_203),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_194),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_168),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_190),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_176),
.B(n_170),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_213),
.B(n_174),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_178),
.B(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_179),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_221),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_188),
.B1(n_193),
.B2(n_210),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_177),
.B1(n_183),
.B2(n_180),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_222),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_210),
.C(n_208),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_212),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_169),
.B(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_211),
.B(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_209),
.C(n_207),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_19),
.C(n_2),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_6),
.C(n_2),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_240),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_222),
.Y(n_239)
);

FAx1_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_8),
.CI(n_3),
.CON(n_246),
.SN(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_7),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_230),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_242),
.B(n_7),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_245),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_5),
.B(n_2),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_8),
.B(n_3),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_238),
.C(n_236),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_239),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_8),
.C2(n_9),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.C(n_249),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_1),
.A3(n_4),
.B1(n_10),
.B2(n_11),
.C1(n_237),
.C2(n_236),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_4),
.B(n_10),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_10),
.C(n_11),
.Y(n_255)
);

NAND2x1p5_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_11),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_1),
.Y(n_257)
);


endmodule