module fake_netlist_5_1251_n_1616 (n_29, n_16, n_43, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_1616);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_1616;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_82;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_111;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_105;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_87;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_51;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_101;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_94;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_59;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_72;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_48;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_114;
wire n_96;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_129;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_49;
wire n_310;
wire n_54;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_70;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_91;
wire n_1565;
wire n_182;
wire n_143;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_117;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_53;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_71;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_121;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_64;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_103;
wire n_97;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_52;
wire n_784;
wire n_110;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_61;
wire n_678;
wire n_697;
wire n_127;
wire n_1222;
wire n_75;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_116;
wire n_284;
wire n_1128;
wire n_139;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_47;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_100;
wire n_1443;
wire n_1008;
wire n_1539;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_133;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_106;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_93;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_122;
wire n_331;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_90;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_123;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_131;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_109;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_88;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_65;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_69;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_73;
wire n_309;
wire n_512;
wire n_1591;
wire n_84;
wire n_130;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_112;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_55;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_102;
wire n_77;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_83;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_58;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_128;
wire n_120;
wire n_327;
wire n_135;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_62;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_136;
wire n_86;
wire n_146;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_74;
wire n_1139;
wire n_515;
wire n_57;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_132;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_50;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_107;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_85;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1516;
wire n_876;
wire n_1190;
wire n_118;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_108;
wire n_487;
wire n_1584;
wire n_665;
wire n_66;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_126;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_89;
wire n_1524;
wire n_1485;
wire n_115;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_137;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_124;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_119;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1281;
wire n_67;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_68;
wire n_867;
wire n_186;
wire n_134;
wire n_587;
wire n_63;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_138;
wire n_961;
wire n_771;
wire n_276;
wire n_95;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_104;
wire n_682;
wire n_1567;
wire n_56;
wire n_141;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_145;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_140;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_78;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_98;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_80;
wire n_1315;
wire n_277;
wire n_1061;
wire n_92;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_79;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_76;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_81;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_60;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_113;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_99;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_1),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_6),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_10),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_78),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_48),
.B1(n_83),
.B2(n_88),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_57),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_83),
.B1(n_88),
.B2(n_52),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_57),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_66),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_110),
.Y(n_142)
);

OR2x6_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_64),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_111),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_118),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_71),
.B1(n_100),
.B2(n_97),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_103),
.B1(n_90),
.B2(n_59),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_111),
.Y(n_151)
);

OR2x6_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_66),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_112),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_112),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_87),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_87),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_77),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

BUFx4f_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_124),
.A2(n_77),
.B1(n_56),
.B2(n_73),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_59),
.B1(n_84),
.B2(n_86),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_119),
.B(n_97),
.Y(n_184)
);

AOI21x1_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_90),
.B(n_84),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_127),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_99),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_105),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_139),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_137),
.B(n_62),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_140),
.B(n_93),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_137),
.B(n_75),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_194),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_167),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_135),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_135),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_132),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_132),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_132),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_144),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_132),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_141),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_189),
.B(n_120),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_137),
.C(n_120),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_117),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

BUFx6f_ASAP7_75t_SL g226 ( 
.A(n_157),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_189),
.B(n_137),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_143),
.B(n_137),
.Y(n_229)
);

BUFx6f_ASAP7_75t_SL g230 ( 
.A(n_157),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_172),
.B(n_137),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_143),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_107),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_127),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_143),
.A2(n_71),
.B1(n_55),
.B2(n_65),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_74),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_143),
.A2(n_117),
.B1(n_81),
.B2(n_65),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_148),
.B(n_126),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_58),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_161),
.A2(n_60),
.B1(n_117),
.B2(n_126),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_171),
.B(n_127),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_186),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_127),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_127),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_149),
.B(n_76),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_198),
.B(n_79),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_157),
.B(n_127),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_168),
.B(n_177),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_149),
.B(n_68),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_150),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_143),
.B(n_139),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_150),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_142),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_150),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_157),
.B(n_117),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_181),
.B(n_70),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_181),
.B(n_80),
.Y(n_265)
);

OR2x2_ASAP7_75t_SL g266 ( 
.A(n_148),
.B(n_177),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_157),
.B(n_117),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_168),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_157),
.B(n_117),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_161),
.A2(n_117),
.B1(n_126),
.B2(n_55),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_143),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_166),
.A2(n_117),
.B(n_134),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_152),
.B(n_117),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_174),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_196),
.B(n_63),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_196),
.B(n_89),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_152),
.B(n_117),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_152),
.A2(n_65),
.B1(n_81),
.B2(n_86),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_92),
.B1(n_69),
.B2(n_72),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_145),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_152),
.B(n_139),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_152),
.B(n_122),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_145),
.Y(n_284)
);

BUFx12f_ASAP7_75t_SL g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_151),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_151),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_179),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_179),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_152),
.A2(n_91),
.B1(n_67),
.B2(n_61),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_166),
.B(n_82),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_202),
.B(n_82),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_158),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_147),
.B(n_122),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_154),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_158),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_153),
.A2(n_69),
.B1(n_72),
.B2(n_92),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_204),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_268),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_212),
.B(n_155),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_192),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_243),
.B(n_82),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_217),
.B(n_182),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_204),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_217),
.B(n_293),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_205),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_214),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_182),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_212),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_208),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_237),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_244),
.A2(n_153),
.B(n_155),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_208),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_214),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_268),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_207),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_215),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_254),
.A2(n_180),
.B(n_193),
.C(n_199),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_215),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_261),
.B(n_162),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_204),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_266),
.A2(n_81),
.B1(n_82),
.B2(n_3),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_209),
.B(n_182),
.Y(n_330)
);

NAND2x2_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_0),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_182),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_182),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_162),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_220),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_247),
.A2(n_162),
.B1(n_147),
.B2(n_156),
.Y(n_337)
);

NOR3xp33_ASAP7_75t_L g338 ( 
.A(n_218),
.B(n_147),
.C(n_156),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_225),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_225),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_235),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_38),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_266),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_156),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_245),
.B(n_2),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_156),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_241),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_236),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_236),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_220),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_250),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_276),
.A2(n_147),
.B1(n_180),
.B2(n_199),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_259),
.B(n_37),
.Y(n_355)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_206),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_259),
.B(n_42),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_238),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_238),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g360 ( 
.A(n_232),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_287),
.B(n_180),
.Y(n_361)
);

NOR2x2_ASAP7_75t_L g362 ( 
.A(n_245),
.B(n_176),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_250),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_233),
.A2(n_4),
.B1(n_9),
.B2(n_11),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_221),
.B(n_203),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_227),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_219),
.A2(n_193),
.B1(n_197),
.B2(n_201),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_287),
.A2(n_197),
.B1(n_193),
.B2(n_178),
.Y(n_370)
);

O2A1O1Ixp33_ASAP7_75t_SL g371 ( 
.A1(n_263),
.A2(n_197),
.B(n_200),
.C(n_187),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_229),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_251),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_277),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_289),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_232),
.A2(n_201),
.B1(n_200),
.B2(n_195),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

AND2x6_ASAP7_75t_SL g380 ( 
.A(n_282),
.B(n_9),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_258),
.Y(n_381)
);

BUFx12f_ASAP7_75t_L g382 ( 
.A(n_271),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_316),
.B(n_366),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_SL g384 ( 
.A(n_364),
.B(n_240),
.C(n_222),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_316),
.B(n_221),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_301),
.B(n_285),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_316),
.A2(n_234),
.B(n_227),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_316),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_322),
.B(n_271),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

BUFx8_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_349),
.B(n_221),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_342),
.A2(n_222),
.B(n_290),
.C(n_270),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_316),
.A2(n_234),
.B(n_227),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_SL g402 ( 
.A(n_307),
.B(n_290),
.C(n_291),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_234),
.B(n_223),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_327),
.B(n_257),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_321),
.B(n_270),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_378),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_303),
.Y(n_410)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_330),
.A2(n_291),
.B(n_228),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_303),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_366),
.A2(n_302),
.B(n_365),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_322),
.B(n_206),
.Y(n_414)
);

A2O1A1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_374),
.A2(n_229),
.B(n_231),
.C(n_283),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_314),
.B(n_210),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_310),
.B(n_211),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_356),
.A2(n_216),
.B1(n_213),
.B2(n_274),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_356),
.A2(n_305),
.B1(n_334),
.B2(n_300),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_356),
.B(n_274),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

O2A1O1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_304),
.A2(n_264),
.B(n_265),
.C(n_297),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_302),
.A2(n_223),
.B(n_252),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_318),
.B(n_221),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_320),
.B(n_226),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_375),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_304),
.B(n_221),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_323),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_356),
.A2(n_334),
.B1(n_300),
.B2(n_302),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_317),
.A2(n_224),
.B(n_239),
.C(n_248),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_303),
.Y(n_433)
);

OR2x6_ASAP7_75t_L g434 ( 
.A(n_355),
.B(n_278),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_315),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_355),
.B(n_280),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_324),
.A2(n_255),
.B(n_249),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_361),
.B(n_221),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_361),
.B(n_221),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_303),
.A2(n_253),
.B(n_246),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_313),
.A2(n_206),
.B(n_267),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

NOR2x1_ASAP7_75t_SL g443 ( 
.A(n_356),
.B(n_253),
.Y(n_443)
);

O2A1O1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_336),
.A2(n_352),
.B(n_353),
.C(n_372),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_300),
.B(n_280),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_SL g446 ( 
.A1(n_338),
.A2(n_272),
.B(n_258),
.C(n_260),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_306),
.A2(n_224),
.B(n_273),
.C(n_269),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_303),
.B(n_295),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_370),
.A2(n_294),
.B(n_295),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_309),
.B(n_206),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_372),
.A2(n_279),
.B(n_275),
.C(n_262),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_326),
.A2(n_260),
.B(n_190),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_SL g453 ( 
.A(n_344),
.B(n_280),
.C(n_230),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_355),
.B(n_280),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_346),
.B(n_226),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_331),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_SL g458 ( 
.A1(n_363),
.A2(n_242),
.B(n_201),
.C(n_176),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_328),
.B(n_206),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_363),
.B(n_206),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_376),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_346),
.A2(n_230),
.B1(n_226),
.B2(n_138),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_357),
.Y(n_463)
);

NAND2x1p5_ASAP7_75t_L g464 ( 
.A(n_357),
.B(n_230),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_348),
.Y(n_465)
);

NOR3xp33_ASAP7_75t_SL g466 ( 
.A(n_329),
.B(n_12),
.C(n_13),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_360),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_340),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_379),
.A2(n_178),
.B1(n_174),
.B2(n_190),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_340),
.A2(n_341),
.B1(n_358),
.B2(n_359),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_299),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_331),
.A2(n_325),
.B1(n_299),
.B2(n_339),
.Y(n_472)
);

AOI21x1_ASAP7_75t_L g473 ( 
.A1(n_319),
.A2(n_201),
.B(n_200),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_341),
.B(n_16),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_332),
.A2(n_347),
.B(n_333),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_319),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_350),
.B(n_17),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_335),
.A2(n_174),
.B(n_178),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_325),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_350),
.B(n_21),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_339),
.B(n_200),
.Y(n_482)
);

INVx6_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_371),
.A2(n_195),
.B(n_191),
.C(n_187),
.Y(n_484)
);

A2O1A1Ixp33_ASAP7_75t_L g485 ( 
.A1(n_358),
.A2(n_195),
.B(n_191),
.C(n_154),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_343),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_348),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_359),
.A2(n_195),
.B(n_191),
.C(n_154),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_351),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_345),
.A2(n_174),
.B(n_190),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_384),
.B(n_466),
.C(n_398),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_414),
.B(n_351),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_405),
.A2(n_308),
.B(n_337),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_407),
.A2(n_384),
.B1(n_463),
.B2(n_453),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_380),
.Y(n_495)
);

INVx8_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_387),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_407),
.A2(n_367),
.B1(n_377),
.B2(n_362),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_406),
.B(n_381),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_415),
.A2(n_354),
.B(n_381),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_411),
.A2(n_175),
.B(n_154),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_390),
.A2(n_401),
.B(n_389),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_406),
.B(n_362),
.Y(n_504)
);

CKINVDCx11_ASAP7_75t_R g505 ( 
.A(n_397),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_449),
.A2(n_191),
.B(n_160),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_453),
.A2(n_175),
.B1(n_187),
.B2(n_183),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_438),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_399),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_437),
.A2(n_173),
.B(n_183),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_427),
.B(n_138),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_429),
.B(n_160),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_417),
.B(n_160),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_441),
.A2(n_432),
.B(n_424),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

AOI21xp33_ASAP7_75t_L g517 ( 
.A1(n_445),
.A2(n_22),
.B(n_23),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_417),
.B(n_176),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_394),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_462),
.B(n_190),
.Y(n_521)
);

AO31x2_ASAP7_75t_L g522 ( 
.A1(n_421),
.A2(n_175),
.A3(n_173),
.B(n_170),
.Y(n_522)
);

A2O1A1Ixp33_ASAP7_75t_L g523 ( 
.A1(n_402),
.A2(n_173),
.B(n_170),
.C(n_138),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_478),
.A2(n_170),
.B(n_190),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_403),
.B(n_170),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_404),
.B(n_190),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_435),
.B(n_22),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_455),
.A2(n_122),
.B1(n_116),
.B2(n_115),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_44),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_408),
.B(n_122),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_394),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_447),
.A2(n_116),
.B(n_115),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_386),
.A2(n_122),
.B1(n_116),
.B2(n_115),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_392),
.B(n_24),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_484),
.A2(n_27),
.B(n_28),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_409),
.B(n_122),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_439),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_R g540 ( 
.A(n_479),
.B(n_30),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_490),
.A2(n_452),
.B(n_413),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_392),
.B(n_436),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_468),
.B(n_30),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_456),
.Y(n_544)
);

AO21x1_ASAP7_75t_L g545 ( 
.A1(n_444),
.A2(n_31),
.B(n_32),
.Y(n_545)
);

OA21x2_ASAP7_75t_L g546 ( 
.A1(n_475),
.A2(n_113),
.B(n_115),
.Y(n_546)
);

OAI21x1_ASAP7_75t_SL g547 ( 
.A1(n_443),
.A2(n_33),
.B(n_34),
.Y(n_547)
);

OAI22x1_ASAP7_75t_L g548 ( 
.A1(n_457),
.A2(n_454),
.B1(n_464),
.B2(n_477),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_391),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_433),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_SL g551 ( 
.A(n_472),
.B(n_33),
.C(n_34),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

OAI22x1_ASAP7_75t_L g553 ( 
.A1(n_464),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_483),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_440),
.A2(n_113),
.B(n_115),
.Y(n_555)
);

AOI211x1_ASAP7_75t_L g556 ( 
.A1(n_460),
.A2(n_113),
.B(n_115),
.C(n_116),
.Y(n_556)
);

AO31x2_ASAP7_75t_L g557 ( 
.A1(n_485),
.A2(n_113),
.A3(n_115),
.B(n_116),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_SL g558 ( 
.A(n_474),
.B(n_113),
.C(n_115),
.Y(n_558)
);

AOI221x1_ASAP7_75t_L g559 ( 
.A1(n_419),
.A2(n_116),
.B1(n_431),
.B2(n_481),
.C(n_477),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_420),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_468),
.B(n_116),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_385),
.A2(n_116),
.B(n_425),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_385),
.A2(n_116),
.B(n_383),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_462),
.B(n_472),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_433),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_450),
.B(n_467),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_383),
.A2(n_446),
.B(n_396),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_461),
.Y(n_568)
);

OA22x2_ASAP7_75t_L g569 ( 
.A1(n_466),
.A2(n_434),
.B1(n_480),
.B2(n_476),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_448),
.A2(n_469),
.B(n_482),
.Y(n_570)
);

AO31x2_ASAP7_75t_L g571 ( 
.A1(n_488),
.A2(n_470),
.A3(n_481),
.B(n_474),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_446),
.A2(n_434),
.B(n_426),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_471),
.B(n_489),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_R g574 ( 
.A(n_434),
.B(n_459),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_487),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

AO31x2_ASAP7_75t_L g577 ( 
.A1(n_486),
.A2(n_393),
.A3(n_400),
.B(n_430),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_448),
.A2(n_465),
.B(n_423),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_483),
.A2(n_456),
.B1(n_467),
.B2(n_486),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_410),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_458),
.A2(n_451),
.B(n_422),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_467),
.B(n_412),
.Y(n_582)
);

AO22x2_ASAP7_75t_L g583 ( 
.A1(n_412),
.A2(n_458),
.B1(n_483),
.B2(n_467),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_422),
.A2(n_316),
.B(n_366),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_405),
.A2(n_316),
.B(n_366),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_398),
.A2(n_415),
.B(n_254),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_429),
.B(n_418),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_473),
.A2(n_449),
.B(n_401),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_387),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_414),
.B(n_392),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_398),
.A2(n_254),
.B(n_244),
.C(n_349),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_407),
.A2(n_398),
.B1(n_384),
.B2(n_266),
.Y(n_592)
);

NOR2xp67_ASAP7_75t_SL g593 ( 
.A(n_397),
.B(n_301),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_456),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_405),
.A2(n_316),
.B(n_366),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_429),
.B(n_418),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_429),
.B(n_418),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_428),
.B(n_321),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_429),
.B(n_418),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_428),
.B(n_349),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_428),
.B(n_321),
.Y(n_601)
);

AOI21xp33_ASAP7_75t_L g602 ( 
.A1(n_407),
.A2(n_254),
.B(n_244),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_524),
.A2(n_506),
.B(n_493),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_559),
.A2(n_515),
.B(n_586),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_SL g605 ( 
.A(n_591),
.B(n_491),
.C(n_545),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_602),
.A2(n_592),
.B1(n_564),
.B2(n_551),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_557),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_581),
.A2(n_562),
.B(n_570),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_577),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_505),
.Y(n_611)
);

AO31x2_ASAP7_75t_L g612 ( 
.A1(n_592),
.A2(n_572),
.A3(n_567),
.B(n_498),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_585),
.A2(n_595),
.B(n_555),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_602),
.B(n_494),
.C(n_539),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_563),
.A2(n_546),
.B(n_578),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_557),
.Y(n_616)
);

AOI21x1_ASAP7_75t_L g617 ( 
.A1(n_501),
.A2(n_546),
.B(n_511),
.Y(n_617)
);

AO21x2_ASAP7_75t_L g618 ( 
.A1(n_500),
.A2(n_536),
.B(n_558),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_496),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_533),
.A2(n_511),
.B(n_584),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_513),
.A2(n_507),
.B(n_531),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_577),
.Y(n_623)
);

AO21x2_ASAP7_75t_L g624 ( 
.A1(n_536),
.A2(n_523),
.B(n_547),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_587),
.A2(n_597),
.B(n_596),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_531),
.A2(n_537),
.B(n_526),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_494),
.A2(n_504),
.B1(n_569),
.B2(n_498),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_529),
.B(n_590),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_537),
.A2(n_526),
.B(n_525),
.Y(n_629)
);

INVx6_ASAP7_75t_SL g630 ( 
.A(n_492),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_587),
.A2(n_599),
.B(n_596),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_522),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_508),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_497),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_503),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_542),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_569),
.A2(n_514),
.B(n_518),
.Y(n_637)
);

AO21x2_ASAP7_75t_L g638 ( 
.A1(n_521),
.A2(n_599),
.B(n_597),
.Y(n_638)
);

AOI221x1_ASAP7_75t_L g639 ( 
.A1(n_517),
.A2(n_548),
.B1(n_539),
.B2(n_583),
.C(n_553),
.Y(n_639)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_514),
.A2(n_518),
.B(n_517),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_509),
.A2(n_565),
.B(n_550),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_589),
.Y(n_642)
);

OA21x2_ASAP7_75t_L g643 ( 
.A1(n_568),
.A2(n_573),
.B(n_561),
.Y(n_643)
);

AO21x2_ASAP7_75t_L g644 ( 
.A1(n_528),
.A2(n_568),
.B(n_573),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_552),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_535),
.B(n_540),
.C(n_543),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_561),
.A2(n_575),
.B(n_560),
.Y(n_647)
);

AO21x2_ASAP7_75t_L g648 ( 
.A1(n_534),
.A2(n_530),
.B(n_499),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_529),
.B(n_590),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_516),
.A2(n_549),
.B(n_580),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_492),
.B(n_566),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g652 ( 
.A1(n_556),
.A2(n_571),
.B(n_574),
.Y(n_652)
);

AO31x2_ASAP7_75t_L g653 ( 
.A1(n_571),
.A2(n_583),
.A3(n_598),
.B(n_601),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_571),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_579),
.A2(n_583),
.B(n_527),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_600),
.A2(n_532),
.B(n_508),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_508),
.A2(n_512),
.B(n_582),
.Y(n_657)
);

NAND2x1p5_ASAP7_75t_L g658 ( 
.A(n_508),
.B(n_593),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_496),
.A2(n_538),
.B(n_594),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_496),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_520),
.B(n_594),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_554),
.A2(n_495),
.B(n_576),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_520),
.B(n_510),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_594),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_544),
.B(n_519),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_491),
.A2(n_346),
.B1(n_266),
.B2(n_407),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_550),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_602),
.A2(n_402),
.B1(n_491),
.B2(n_592),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_541),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_598),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_550),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_508),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_587),
.B(n_596),
.Y(n_674)
);

CKINVDCx11_ASAP7_75t_R g675 ( 
.A(n_505),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_587),
.B(n_596),
.Y(n_676)
);

AO21x2_ASAP7_75t_L g677 ( 
.A1(n_586),
.A2(n_515),
.B(n_602),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_529),
.B(n_590),
.Y(n_678)
);

AOI21x1_ASAP7_75t_L g679 ( 
.A1(n_581),
.A2(n_502),
.B(n_493),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_592),
.B(n_587),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_602),
.A2(n_586),
.B(n_591),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_592),
.B(n_587),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_602),
.A2(n_402),
.B1(n_491),
.B2(n_592),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_550),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_577),
.Y(n_685)
);

OA21x2_ASAP7_75t_L g686 ( 
.A1(n_559),
.A2(n_515),
.B(n_586),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_588),
.A2(n_502),
.B(n_541),
.Y(n_687)
);

AO21x2_ASAP7_75t_L g688 ( 
.A1(n_586),
.A2(n_515),
.B(n_602),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_577),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_588),
.A2(n_502),
.B(n_541),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_577),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_559),
.A2(n_411),
.A3(n_398),
.B(n_581),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_577),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_602),
.A2(n_591),
.B(n_592),
.C(n_586),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_588),
.A2(n_502),
.B(n_541),
.Y(n_695)
);

OAI21x1_ASAP7_75t_SL g696 ( 
.A1(n_500),
.A2(n_567),
.B(n_572),
.Y(n_696)
);

AO21x2_ASAP7_75t_L g697 ( 
.A1(n_586),
.A2(n_515),
.B(n_602),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_505),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_588),
.A2(n_502),
.B(n_541),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_496),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_588),
.A2(n_502),
.B(n_541),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_602),
.A2(n_402),
.B1(n_491),
.B2(n_592),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_677),
.B(n_688),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_677),
.B(n_688),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_631),
.A2(n_681),
.B(n_694),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_694),
.A2(n_614),
.B(n_681),
.C(n_606),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_667),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_674),
.B(n_676),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_677),
.B(n_688),
.Y(n_709)
);

AOI21x1_ASAP7_75t_SL g710 ( 
.A1(n_661),
.A2(n_676),
.B(n_674),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_631),
.A2(n_625),
.B(n_641),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_625),
.B(n_666),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_667),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_677),
.B(n_688),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_636),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_666),
.B(n_668),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_683),
.A2(n_702),
.B1(n_670),
.B2(n_627),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_673),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_697),
.B(n_612),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_635),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_673),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_614),
.A2(n_646),
.B1(n_682),
.B2(n_680),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_660),
.B(n_635),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_680),
.B(n_682),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_697),
.B(n_612),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_612),
.B(n_654),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_697),
.B(n_612),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_697),
.B(n_612),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_673),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_605),
.A2(n_646),
.B(n_696),
.C(n_662),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_675),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_634),
.Y(n_732)
);

OA21x2_ASAP7_75t_L g733 ( 
.A1(n_608),
.A2(n_639),
.B(n_615),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_612),
.B(n_653),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_671),
.B(n_684),
.Y(n_735)
);

O2A1O1Ixp5_ASAP7_75t_L g736 ( 
.A1(n_654),
.A2(n_662),
.B(n_679),
.C(n_632),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_635),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_673),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_SL g739 ( 
.A1(n_604),
.A2(n_686),
.B(n_658),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_605),
.A2(n_696),
.B(n_661),
.C(n_658),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_660),
.B(n_651),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_609),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_673),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_653),
.B(n_654),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_628),
.A2(n_678),
.B1(n_649),
.B2(n_651),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_655),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_608),
.A2(n_639),
.B(n_615),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_663),
.A2(n_651),
.B1(n_658),
.B2(n_665),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_SL g750 ( 
.A1(n_604),
.A2(n_686),
.B(n_648),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_SL g751 ( 
.A1(n_604),
.A2(n_686),
.B(n_648),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_SL g752 ( 
.A1(n_611),
.A2(n_698),
.B1(n_665),
.B2(n_660),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_L g753 ( 
.A1(n_618),
.A2(n_642),
.B1(n_634),
.B2(n_645),
.C(n_651),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_653),
.B(n_638),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_653),
.B(n_638),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_628),
.B(n_678),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_647),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_628),
.B(n_678),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_628),
.B(n_678),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_618),
.A2(n_642),
.B(n_648),
.C(n_645),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_657),
.A2(n_656),
.B(n_655),
.C(n_613),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_690),
.A2(n_620),
.B(n_699),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_653),
.B(n_638),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_647),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_621),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_653),
.B(n_638),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_643),
.B(n_652),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_618),
.A2(n_648),
.B(n_624),
.C(n_664),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_SL g769 ( 
.A1(n_644),
.A2(n_618),
.B(n_700),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_623),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_652),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_649),
.B(n_619),
.Y(n_772)
);

AOI21x1_ASAP7_75t_SL g773 ( 
.A1(n_649),
.A2(n_656),
.B(n_624),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_621),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_690),
.A2(n_620),
.B(n_699),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_649),
.B(n_643),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_619),
.B(n_700),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_613),
.A2(n_673),
.B(n_644),
.Y(n_778)
);

O2A1O1Ixp5_ASAP7_75t_L g779 ( 
.A1(n_669),
.A2(n_616),
.B(n_607),
.C(n_610),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_673),
.B(n_664),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_619),
.A2(n_700),
.B1(n_630),
.B2(n_633),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_692),
.B(n_691),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_685),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_643),
.B(n_644),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_643),
.B(n_652),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_685),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_652),
.B(n_637),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_657),
.A2(n_637),
.B(n_622),
.C(n_659),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_624),
.A2(n_640),
.B(n_644),
.C(n_669),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_624),
.A2(n_640),
.B(n_633),
.C(n_691),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_637),
.B(n_692),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_742),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_706),
.B(n_633),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_787),
.B(n_791),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_742),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_757),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_787),
.B(n_607),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_713),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_737),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_746),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_769),
.B(n_701),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_748),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_778),
.A2(n_695),
.B(n_687),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_748),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_764),
.B(n_607),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_724),
.B(n_705),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_791),
.B(n_610),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_765),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_770),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_755),
.B(n_692),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_774),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_774),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_737),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_786),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_750),
.A2(n_617),
.B(n_689),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_755),
.B(n_692),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_786),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_761),
.B(n_616),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_783),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_770),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_719),
.B(n_616),
.Y(n_822)
);

AO21x1_ASAP7_75t_SL g823 ( 
.A1(n_782),
.A2(n_693),
.B(n_689),
.Y(n_823)
);

AOI222xp33_ASAP7_75t_L g824 ( 
.A1(n_716),
.A2(n_693),
.B1(n_633),
.B2(n_629),
.C1(n_622),
.C2(n_626),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_718),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_719),
.B(n_616),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_732),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_720),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_725),
.B(n_610),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_713),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_720),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_722),
.B(n_640),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_767),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_777),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_782),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_767),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_725),
.B(n_727),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_776),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_788),
.B(n_723),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_746),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_744),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_711),
.A2(n_617),
.B(n_672),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_784),
.B(n_726),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_707),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_726),
.B(n_692),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_727),
.B(n_610),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_728),
.B(n_692),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_785),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_703),
.B(n_672),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_723),
.B(n_623),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_771),
.Y(n_852)
);

BUFx4f_ASAP7_75t_SL g853 ( 
.A(n_715),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_771),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_785),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_723),
.B(n_623),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_762),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_750),
.A2(n_672),
.B(n_603),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_754),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_760),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_734),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_734),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_754),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_712),
.B(n_640),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_728),
.B(n_626),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_763),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_833),
.B(n_704),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_792),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_807),
.B(n_763),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_792),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_796),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_833),
.B(n_709),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_795),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_839),
.B(n_833),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_795),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_839),
.B(n_709),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_803),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_794),
.B(n_766),
.Y(n_879)
);

OAI221xp5_ASAP7_75t_SL g880 ( 
.A1(n_832),
.A2(n_730),
.B1(n_753),
.B2(n_751),
.C(n_740),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_794),
.B(n_766),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_803),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_800),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_793),
.A2(n_717),
.B1(n_749),
.B2(n_708),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_805),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_836),
.B(n_714),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_800),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_805),
.Y(n_888)
);

OA21x2_ASAP7_75t_L g889 ( 
.A1(n_804),
.A2(n_779),
.B(n_736),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_794),
.B(n_714),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_800),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_840),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_836),
.B(n_704),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_853),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_807),
.B(n_703),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_852),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_836),
.B(n_747),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_848),
.B(n_747),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_848),
.B(n_747),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_848),
.B(n_733),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_837),
.B(n_733),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_839),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_857),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_837),
.B(n_733),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_838),
.B(n_735),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_809),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_852),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_853),
.A2(n_832),
.B1(n_860),
.B2(n_745),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_838),
.B(n_751),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_855),
.B(n_769),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_857),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_809),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_839),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_837),
.B(n_865),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_812),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_865),
.B(n_739),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_857),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_857),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_857),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_813),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_867),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_855),
.B(n_739),
.Y(n_922)
);

OAI221xp5_ASAP7_75t_L g923 ( 
.A1(n_793),
.A2(n_768),
.B1(n_731),
.B2(n_752),
.C(n_781),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_840),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_865),
.B(n_789),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_839),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_813),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_864),
.B(n_790),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_815),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_815),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_855),
.B(n_775),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_854),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_867),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_798),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_867),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_867),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_840),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_863),
.B(n_775),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_830),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_854),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_818),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_830),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_835),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_863),
.B(n_775),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_822),
.B(n_762),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_818),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_820),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_820),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_883),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_894),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_914),
.B(n_866),
.Y(n_952)
);

OA21x2_ASAP7_75t_L g953 ( 
.A1(n_928),
.A2(n_860),
.B(n_804),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_894),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_914),
.B(n_866),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_891),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_934),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_896),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_872),
.Y(n_959)
);

AOI221xp5_ASAP7_75t_L g960 ( 
.A1(n_880),
.A2(n_864),
.B1(n_844),
.B2(n_861),
.C(n_862),
.Y(n_960)
);

AND4x1_ASAP7_75t_L g961 ( 
.A(n_884),
.B(n_824),
.C(n_861),
.D(n_862),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_947),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_883),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_L g964 ( 
.A1(n_880),
.A2(n_844),
.B1(n_866),
.B2(n_847),
.C(n_859),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_883),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_947),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_875),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_884),
.A2(n_756),
.B1(n_847),
.B2(n_741),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_923),
.A2(n_741),
.B1(n_772),
.B2(n_756),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_923),
.A2(n_758),
.B1(n_759),
.B2(n_834),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_875),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_895),
.B(n_859),
.Y(n_972)
);

OAI31xp33_ASAP7_75t_L g973 ( 
.A1(n_908),
.A2(n_819),
.A3(n_756),
.B(n_847),
.Y(n_973)
);

AOI31xp33_ASAP7_75t_L g974 ( 
.A1(n_908),
.A2(n_731),
.A3(n_824),
.B(n_777),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_870),
.A2(n_741),
.B1(n_772),
.B2(n_630),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_896),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_891),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_928),
.A2(n_819),
.B(n_827),
.Y(n_978)
);

NAND4xp25_ASAP7_75t_L g979 ( 
.A(n_895),
.B(n_870),
.C(n_909),
.D(n_905),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_875),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_905),
.B(n_909),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_R g982 ( 
.A(n_934),
.B(n_718),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_875),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_947),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_910),
.B(n_835),
.C(n_843),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_939),
.A2(n_819),
.B(n_827),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_948),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_875),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_910),
.B(n_843),
.C(n_819),
.Y(n_989)
);

AO21x2_ASAP7_75t_L g990 ( 
.A1(n_911),
.A2(n_842),
.B(n_804),
.Y(n_990)
);

OAI332xp33_ASAP7_75t_L g991 ( 
.A1(n_910),
.A2(n_811),
.A3(n_817),
.B1(n_843),
.B2(n_845),
.B3(n_851),
.C1(n_841),
.C2(n_814),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_R g992 ( 
.A(n_891),
.B(n_819),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_890),
.B(n_798),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_948),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_L g995 ( 
.A(n_925),
.B(n_798),
.C(n_811),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_890),
.B(n_841),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_914),
.B(n_834),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_L g998 ( 
.A(n_925),
.B(n_817),
.C(n_811),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_875),
.Y(n_999)
);

OAI221xp5_ASAP7_75t_SL g1000 ( 
.A1(n_922),
.A2(n_817),
.B1(n_845),
.B2(n_849),
.C(n_801),
.Y(n_1000)
);

AOI31xp33_ASAP7_75t_L g1001 ( 
.A1(n_902),
.A2(n_777),
.A3(n_845),
.B(n_772),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_922),
.A2(n_834),
.B1(n_825),
.B2(n_802),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_925),
.A2(n_822),
.B(n_826),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_890),
.B(n_851),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_939),
.A2(n_799),
.B1(n_814),
.B2(n_828),
.C(n_831),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_879),
.B(n_808),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_916),
.A2(n_799),
.B1(n_814),
.B2(n_828),
.C(n_831),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_L g1008 ( 
.A(n_922),
.B(n_849),
.C(n_799),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_948),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_879),
.B(n_808),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_879),
.B(n_808),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_883),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_887),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_869),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_916),
.A2(n_630),
.B1(n_829),
.B2(n_846),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_902),
.B(n_913),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_916),
.A2(n_630),
.B1(n_829),
.B2(n_846),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_942),
.A2(n_846),
.B1(n_829),
.B2(n_826),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_868),
.B(n_849),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_872),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_869),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_902),
.A2(n_913),
.B1(n_926),
.B2(n_877),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_942),
.A2(n_822),
.B1(n_826),
.B2(n_816),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_887),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_881),
.B(n_797),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_887),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_871),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_881),
.B(n_797),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_868),
.B(n_797),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_907),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_877),
.A2(n_816),
.B1(n_802),
.B2(n_825),
.Y(n_1032)
);

AOI331xp33_ASAP7_75t_L g1033 ( 
.A1(n_871),
.A2(n_710),
.A3(n_823),
.B1(n_842),
.B2(n_773),
.B3(n_816),
.C1(n_801),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_902),
.A2(n_802),
.B1(n_825),
.B2(n_743),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_907),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_881),
.B(n_856),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_871),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_R g1038 ( 
.A(n_913),
.B(n_729),
.Y(n_1038)
);

AOI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_901),
.A2(n_856),
.B1(n_850),
.B2(n_806),
.C(n_821),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_868),
.B(n_856),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_887),
.B(n_721),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_886),
.B(n_856),
.Y(n_1042)
);

AO21x2_ASAP7_75t_L g1043 ( 
.A1(n_911),
.A2(n_842),
.B(n_816),
.Y(n_1043)
);

INVx5_ASAP7_75t_L g1044 ( 
.A(n_903),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_924),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_913),
.A2(n_802),
.B1(n_825),
.B2(n_743),
.Y(n_1046)
);

OAI33xp33_ASAP7_75t_L g1047 ( 
.A1(n_874),
.A2(n_821),
.A3(n_810),
.B1(n_823),
.B2(n_816),
.B3(n_858),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_926),
.B(n_801),
.Y(n_1048)
);

OAI211xp5_ASAP7_75t_SL g1049 ( 
.A1(n_911),
.A2(n_867),
.B(n_821),
.C(n_823),
.Y(n_1049)
);

OAI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_926),
.A2(n_802),
.B1(n_825),
.B2(n_801),
.C(n_780),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_874),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_926),
.A2(n_825),
.B1(n_802),
.B2(n_743),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_874),
.Y(n_1053)
);

AOI22x1_ASAP7_75t_L g1054 ( 
.A1(n_892),
.A2(n_825),
.B1(n_802),
.B2(n_738),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_901),
.A2(n_850),
.B(n_856),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_924),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1012),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_1017),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_1038),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1017),
.B(n_877),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1015),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_959),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_981),
.B(n_943),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1022),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1028),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_951),
.B(n_877),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1037),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_1017),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_959),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_988),
.B(n_901),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1021),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1021),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1051),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_988),
.B(n_904),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1043),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1053),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_962),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_958),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1043),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_966),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_950),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_1044),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_984),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1038),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_987),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_994),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_961),
.B(n_974),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_963),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1009),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_998),
.B(n_886),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_973),
.B(n_892),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_1032),
.A2(n_917),
.B(n_919),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_SL g1093 ( 
.A(n_964),
.B(n_892),
.C(n_937),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_951),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_990),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_958),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_982),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_990),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_976),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_976),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1031),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1044),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1031),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_982),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1035),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1044),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1035),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1020),
.Y(n_1108)
);

INVx4_ASAP7_75t_SL g1109 ( 
.A(n_1041),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1033),
.A2(n_801),
.B(n_932),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1044),
.Y(n_1111)
);

INVx4_ASAP7_75t_SL g1112 ( 
.A(n_1041),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_956),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1048),
.B(n_877),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1041),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_960),
.A2(n_932),
.B(n_940),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_956),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_977),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_1041),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_996),
.Y(n_1120)
);

CKINVDCx6p67_ASAP7_75t_R g1121 ( 
.A(n_954),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_1041),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_977),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_1025),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_999),
.B(n_904),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_953),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_999),
.B(n_904),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1004),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_965),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_972),
.B(n_886),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_967),
.B(n_945),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_970),
.B(n_940),
.C(n_943),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_953),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1030),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1048),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_953),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_971),
.B(n_945),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1040),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1042),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_980),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1056),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_985),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1048),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1056),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1026),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1029),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1008),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1057),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1142),
.B(n_979),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1059),
.B(n_952),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1057),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1061),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1121),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1061),
.Y(n_1154)
);

AOI31xp33_ASAP7_75t_L g1155 ( 
.A1(n_1087),
.A2(n_969),
.A3(n_992),
.B(n_1052),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1064),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1142),
.B(n_1003),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1059),
.B(n_955),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_1132),
.B(n_968),
.C(n_1024),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1147),
.B(n_1007),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1064),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1107),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1065),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1084),
.B(n_1006),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1147),
.B(n_1090),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_SL g1166 ( 
.A1(n_1091),
.A2(n_995),
.B1(n_978),
.B2(n_989),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1065),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1084),
.B(n_1097),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1097),
.B(n_1010),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1067),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1094),
.B(n_1121),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1063),
.B(n_1005),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1063),
.B(n_991),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1126),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1107),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1126),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1104),
.B(n_1011),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1109),
.B(n_986),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1104),
.B(n_1036),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1109),
.B(n_1032),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1113),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1102),
.A2(n_1068),
.B(n_1058),
.Y(n_1182)
);

OAI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1091),
.A2(n_1093),
.B1(n_1132),
.B2(n_1116),
.C(n_1094),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1115),
.B(n_997),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1067),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1115),
.B(n_983),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1073),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1119),
.B(n_1023),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1073),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_R g1190 ( 
.A(n_1094),
.B(n_937),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1093),
.A2(n_1033),
.B(n_1000),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1126),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1113),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1076),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1145),
.B(n_993),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1119),
.B(n_1122),
.Y(n_1196)
);

NOR3xp33_ASAP7_75t_L g1197 ( 
.A(n_1094),
.B(n_1050),
.C(n_1047),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1122),
.B(n_1013),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1121),
.B(n_1066),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1109),
.B(n_1025),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1141),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1141),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1145),
.B(n_957),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1109),
.B(n_1027),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1078),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1146),
.B(n_1019),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1146),
.B(n_1139),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1090),
.B(n_1000),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1133),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1105),
.B(n_1019),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1076),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1143),
.A2(n_968),
.B1(n_975),
.B2(n_1016),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1109),
.B(n_1027),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1105),
.B(n_1024),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1112),
.B(n_1014),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1130),
.B(n_873),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1130),
.B(n_873),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1134),
.B(n_873),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1133),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1078),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1112),
.B(n_877),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1077),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1077),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1134),
.B(n_873),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1112),
.B(n_1052),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1110),
.B(n_1054),
.C(n_975),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1112),
.B(n_1045),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1080),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1081),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1229),
.B(n_1120),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1220),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1162),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1168),
.B(n_1060),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1168),
.B(n_1060),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1175),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1202),
.B(n_1196),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1193),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1148),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1225),
.B(n_1221),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1165),
.B(n_1096),
.Y(n_1240)
);

NOR5xp2_ASAP7_75t_L g1241 ( 
.A(n_1183),
.B(n_1116),
.C(n_1049),
.D(n_1103),
.E(n_1101),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1202),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1148),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1174),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1151),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1151),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1152),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1152),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1161),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1165),
.B(n_1096),
.Y(n_1250)
);

NAND2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1153),
.B(n_1082),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1174),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1181),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1214),
.B(n_1099),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1225),
.B(n_1060),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1176),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1214),
.B(n_1099),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1176),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1161),
.Y(n_1259)
);

NAND4xp25_ASAP7_75t_L g1260 ( 
.A(n_1191),
.B(n_1110),
.C(n_1016),
.D(n_1018),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1221),
.B(n_1060),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1196),
.B(n_1112),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1210),
.B(n_1100),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1227),
.B(n_1102),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1167),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1171),
.B(n_1139),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1180),
.B(n_1114),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1180),
.B(n_1114),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1149),
.B(n_1120),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1192),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1173),
.B(n_1128),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1227),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1167),
.Y(n_1273)
);

OAI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1166),
.A2(n_1018),
.B(n_1055),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1199),
.B(n_1160),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1180),
.B(n_1114),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1190),
.Y(n_1277)
);

NAND2xp33_ASAP7_75t_L g1278 ( 
.A(n_1197),
.B(n_1082),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1170),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1200),
.B(n_1114),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1200),
.B(n_1114),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1150),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1208),
.A2(n_1068),
.B1(n_1058),
.B2(n_1135),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1204),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1210),
.B(n_1206),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1205),
.B(n_1100),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1170),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1204),
.B(n_1144),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1192),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1185),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1185),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1236),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1242),
.B(n_1201),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1247),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1282),
.B(n_1157),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1247),
.Y(n_1296)
);

NOR2x1_ASAP7_75t_L g1297 ( 
.A(n_1242),
.B(n_1155),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1253),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1239),
.B(n_1150),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1248),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1236),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1236),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1278),
.A2(n_1159),
.B(n_1172),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1275),
.B(n_1208),
.Y(n_1304)
);

AOI21xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1285),
.A2(n_1277),
.B(n_1251),
.Y(n_1305)
);

BUFx2_ASAP7_75t_SL g1306 ( 
.A(n_1262),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1230),
.B(n_1207),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1251),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1251),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1262),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1239),
.B(n_1158),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1240),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1285),
.B(n_1269),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1248),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_SL g1315 ( 
.A(n_1264),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1288),
.A2(n_1182),
.B(n_1102),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1272),
.B(n_1158),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1274),
.A2(n_1226),
.B1(n_1212),
.B2(n_1178),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1233),
.B(n_1184),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1232),
.B(n_1164),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1235),
.B(n_1164),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1249),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1278),
.B(n_1179),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1284),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1240),
.Y(n_1326)
);

AND2x2_ASAP7_75t_SL g1327 ( 
.A(n_1241),
.B(n_1178),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1271),
.B(n_1169),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1263),
.B(n_1254),
.Y(n_1329)
);

AOI222xp33_ASAP7_75t_L g1330 ( 
.A1(n_1231),
.A2(n_1178),
.B1(n_1047),
.B2(n_1188),
.C1(n_1177),
.C2(n_1203),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1263),
.B(n_1195),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1264),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1249),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1259),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1284),
.B(n_1213),
.Y(n_1335)
);

NOR2x1_ASAP7_75t_L g1336 ( 
.A(n_1231),
.B(n_1264),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1266),
.B(n_1179),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1288),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1259),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_1233),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1265),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_R g1342 ( 
.A(n_1254),
.B(n_1213),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1234),
.A2(n_1255),
.B1(n_1267),
.B2(n_1276),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1260),
.A2(n_1177),
.B1(n_1188),
.B2(n_1143),
.Y(n_1344)
);

AOI222xp33_ASAP7_75t_L g1345 ( 
.A1(n_1255),
.A2(n_1143),
.B1(n_1198),
.B2(n_1088),
.C1(n_1081),
.C2(n_1129),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1234),
.B(n_1184),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1250),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1250),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1280),
.B(n_1215),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1257),
.B(n_1216),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1336),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1299),
.B(n_1280),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1327),
.A2(n_1267),
.B1(n_1268),
.B2(n_1276),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1312),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_R g1355 ( 
.A(n_1342),
.B(n_1286),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1312),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1308),
.B(n_1332),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1327),
.A2(n_1268),
.B1(n_1257),
.B2(n_1281),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1326),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1298),
.B(n_1286),
.Y(n_1361)
);

AOI211xp5_ASAP7_75t_L g1362 ( 
.A1(n_1303),
.A2(n_1281),
.B(n_1246),
.C(n_1243),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1310),
.B(n_1238),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1297),
.A2(n_1182),
.B(n_1245),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1326),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1304),
.A2(n_1287),
.B1(n_1279),
.B2(n_1273),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1304),
.B(n_1265),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1329),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1292),
.B(n_1290),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1342),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1315),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1340),
.A2(n_1261),
.B1(n_1001),
.B2(n_1143),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1294),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1317),
.B(n_1216),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1292),
.B(n_1290),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1296),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1344),
.A2(n_1261),
.B1(n_1143),
.B2(n_1129),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1344),
.A2(n_1143),
.B1(n_1088),
.B2(n_1068),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1318),
.A2(n_1291),
.B(n_1215),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1300),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1314),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1301),
.B(n_1291),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1311),
.B(n_1198),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1301),
.B(n_1154),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1308),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1322),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1330),
.A2(n_1143),
.B1(n_1135),
.B2(n_1058),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1324),
.A2(n_1068),
.B1(n_1058),
.B2(n_1135),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1302),
.B(n_1156),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1302),
.B(n_1163),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1345),
.B(n_1082),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1306),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1305),
.B(n_1252),
.C(n_1244),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1333),
.Y(n_1394)
);

AOI31xp33_ASAP7_75t_L g1395 ( 
.A1(n_1324),
.A2(n_1313),
.A3(n_1293),
.B(n_1337),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_1187),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1349),
.B(n_1186),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1319),
.B(n_1186),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1295),
.A2(n_992),
.B1(n_1082),
.B2(n_1144),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1334),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1332),
.B(n_1144),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1308),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1339),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1341),
.Y(n_1404)
);

AOI222xp33_ASAP7_75t_L g1405 ( 
.A1(n_1337),
.A2(n_1289),
.B1(n_1270),
.B2(n_1258),
.C1(n_1256),
.C2(n_1252),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1332),
.B(n_1244),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1347),
.A2(n_1082),
.B1(n_1144),
.B2(n_1118),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1325),
.B(n_1194),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1371),
.B(n_1328),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1358),
.B(n_1320),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1351),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1392),
.B(n_1325),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1370),
.B(n_1348),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1354),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1387),
.A2(n_1343),
.B1(n_1335),
.B2(n_1346),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1355),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1356),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1360),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1355),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1365),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1370),
.B(n_1321),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_SL g1422 ( 
.A(n_1359),
.B(n_1309),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1357),
.B(n_1335),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1352),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1361),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1395),
.B(n_1323),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1368),
.B(n_1335),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_L g1428 ( 
.A(n_1367),
.B(n_1364),
.C(n_1351),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1369),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1362),
.B(n_1353),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1391),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1379),
.B(n_1307),
.Y(n_1432)
);

AND2x4_ASAP7_75t_SL g1433 ( 
.A(n_1383),
.B(n_1309),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1366),
.B(n_1406),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1363),
.B(n_1391),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1366),
.B(n_1331),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1401),
.Y(n_1437)
);

OAI31xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1377),
.A2(n_1316),
.A3(n_1258),
.B(n_1289),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1398),
.B(n_1397),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1375),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1406),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1382),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1384),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1397),
.B(n_1385),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1407),
.B(n_1316),
.Y(n_1445)
);

AND2x2_ASAP7_75t_SL g1446 ( 
.A(n_1373),
.B(n_1350),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1385),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_1256),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1389),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1402),
.B(n_1270),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1405),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1423),
.B(n_1399),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_1428),
.B(n_1393),
.C(n_1378),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1434),
.A2(n_1407),
.B(n_1399),
.C(n_1404),
.Y(n_1454)
);

AOI221x1_ASAP7_75t_L g1455 ( 
.A1(n_1428),
.A2(n_1376),
.B1(n_1403),
.B2(n_1400),
.C(n_1380),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1445),
.A2(n_1396),
.B(n_1408),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1419),
.A2(n_1372),
.B1(n_1386),
.B2(n_1381),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1409),
.B(n_1374),
.Y(n_1458)
);

OAI211xp5_ASAP7_75t_L g1459 ( 
.A1(n_1430),
.A2(n_1390),
.B(n_1394),
.C(n_1388),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1445),
.A2(n_1219),
.B(n_1209),
.Y(n_1460)
);

OAI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1422),
.A2(n_1082),
.B1(n_1102),
.B2(n_1106),
.C(n_1111),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1435),
.B(n_1082),
.C(n_1209),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1446),
.Y(n_1463)
);

NAND4xp25_ASAP7_75t_L g1464 ( 
.A(n_1409),
.B(n_1219),
.C(n_1135),
.D(n_1106),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1423),
.B(n_1117),
.Y(n_1465)
);

AOI322xp5_ASAP7_75t_L g1466 ( 
.A1(n_1426),
.A2(n_1133),
.A3(n_1136),
.B1(n_1079),
.B2(n_1075),
.C1(n_1101),
.C2(n_1103),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1447),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1431),
.A2(n_1117),
.B1(n_1118),
.B2(n_1123),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1435),
.A2(n_1106),
.B(n_1111),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1436),
.A2(n_1111),
.B(n_1136),
.C(n_1223),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1432),
.A2(n_1136),
.B1(n_1117),
.B2(n_1123),
.C(n_1118),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1438),
.A2(n_1123),
.B1(n_1228),
.B2(n_1223),
.C(n_1222),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1446),
.Y(n_1473)
);

NOR4xp25_ASAP7_75t_SL g1474 ( 
.A(n_1414),
.B(n_1228),
.C(n_1189),
.D(n_1222),
.Y(n_1474)
);

NOR4xp25_ASAP7_75t_L g1475 ( 
.A(n_1441),
.B(n_1189),
.C(n_1211),
.D(n_1075),
.Y(n_1475)
);

NAND4xp25_ASAP7_75t_L g1476 ( 
.A(n_1415),
.B(n_1211),
.C(n_1039),
.D(n_1002),
.Y(n_1476)
);

OAI211xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1410),
.A2(n_1075),
.B(n_1079),
.C(n_1095),
.Y(n_1477)
);

OAI211xp5_ASAP7_75t_L g1478 ( 
.A1(n_1412),
.A2(n_1092),
.B(n_1079),
.C(n_1095),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1413),
.A2(n_1092),
.B(n_1124),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1421),
.A2(n_1092),
.B1(n_1124),
.B2(n_1034),
.C(n_1046),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1439),
.A2(n_1049),
.B(n_1124),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1427),
.B(n_1424),
.C(n_1437),
.D(n_1444),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1425),
.A2(n_1095),
.B1(n_1098),
.B2(n_1080),
.C(n_1086),
.Y(n_1483)
);

OAI33xp33_ASAP7_75t_L g1484 ( 
.A1(n_1417),
.A2(n_1098),
.A3(n_1224),
.B1(n_1218),
.B2(n_1083),
.B3(n_1086),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1443),
.A2(n_1092),
.B1(n_1224),
.B2(n_1218),
.C(n_1098),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1411),
.A2(n_1083),
.B1(n_1108),
.B2(n_1128),
.C(n_1062),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1473),
.Y(n_1487)
);

OA211x2_ASAP7_75t_L g1488 ( 
.A1(n_1452),
.A2(n_1447),
.B(n_1411),
.C(n_1448),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1453),
.A2(n_1433),
.B1(n_1420),
.B2(n_1418),
.Y(n_1489)
);

XOR2x2_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1449),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1463),
.B(n_1429),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1467),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1482),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1458),
.B(n_1440),
.Y(n_1494)
);

AOI21xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1454),
.A2(n_1442),
.B(n_1450),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1451),
.A2(n_1092),
.B1(n_1108),
.B2(n_1138),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1457),
.A2(n_1217),
.B1(n_1138),
.B2(n_1085),
.Y(n_1497)
);

OAI32xp33_ASAP7_75t_L g1498 ( 
.A1(n_1461),
.A2(n_1217),
.A3(n_924),
.B1(n_1070),
.B2(n_1074),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1456),
.A2(n_659),
.B(n_1138),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1465),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1457),
.A2(n_1468),
.B1(n_1472),
.B2(n_1462),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1459),
.A2(n_1085),
.B(n_1089),
.C(n_1069),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1455),
.Y(n_1503)
);

AOI221xp5_ASAP7_75t_L g1504 ( 
.A1(n_1469),
.A2(n_1062),
.B1(n_1069),
.B2(n_1071),
.C(n_1072),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1476),
.A2(n_801),
.B1(n_889),
.B2(n_1069),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1480),
.A2(n_1089),
.B1(n_1085),
.B2(n_1140),
.Y(n_1506)
);

OAI211xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1470),
.A2(n_1062),
.B(n_1072),
.C(n_1071),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1460),
.A2(n_1089),
.B(n_1071),
.C(n_1072),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1464),
.B(n_1140),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1484),
.A2(n_889),
.B1(n_1140),
.B2(n_924),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1486),
.Y(n_1511)
);

AOI211x1_ASAP7_75t_SL g1512 ( 
.A1(n_1471),
.A2(n_911),
.B(n_917),
.C(n_918),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1475),
.A2(n_1127),
.B1(n_1125),
.B2(n_1074),
.C(n_1070),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1466),
.A2(n_1479),
.B(n_1481),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_SL g1515 ( 
.A(n_1474),
.B(n_1074),
.C(n_1070),
.Y(n_1515)
);

INVxp67_ASAP7_75t_SL g1516 ( 
.A(n_1483),
.Y(n_1516)
);

INVxp33_ASAP7_75t_SL g1517 ( 
.A(n_1477),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1487),
.B(n_1478),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1492),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1500),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1503),
.B(n_1493),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1495),
.B(n_1517),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1489),
.B(n_1490),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1491),
.B(n_1501),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1494),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1511),
.B(n_1125),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1488),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1515),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1515),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1514),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1498),
.A2(n_1127),
.B1(n_1125),
.B2(n_937),
.C(n_1131),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1497),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1506),
.B(n_1505),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1127),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1512),
.B(n_1131),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1496),
.B(n_1131),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_L g1539 ( 
.A(n_1507),
.B(n_1137),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1510),
.B(n_1137),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_L g1541 ( 
.A(n_1504),
.B(n_718),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1502),
.Y(n_1542)
);

NAND4xp75_ASAP7_75t_L g1543 ( 
.A(n_1532),
.B(n_1513),
.C(n_1507),
.D(n_1508),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_R g1544 ( 
.A(n_1542),
.B(n_718),
.Y(n_1544)
);

INVx3_ASAP7_75t_SL g1545 ( 
.A(n_1519),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1523),
.B(n_1137),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1522),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1530),
.B(n_903),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1527),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1524),
.A2(n_1540),
.B1(n_1528),
.B2(n_1521),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1531),
.Y(n_1551)
);

XNOR2xp5_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_889),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_SL g1553 ( 
.A(n_1518),
.B(n_721),
.Y(n_1553)
);

NAND4xp75_ASAP7_75t_L g1554 ( 
.A(n_1524),
.B(n_931),
.C(n_889),
.D(n_938),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1529),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1526),
.B(n_721),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_903),
.Y(n_1557)
);

AO22x2_ASAP7_75t_L g1558 ( 
.A1(n_1535),
.A2(n_917),
.B1(n_918),
.B2(n_919),
.Y(n_1558)
);

OAI322xp33_ASAP7_75t_L g1559 ( 
.A1(n_1538),
.A2(n_917),
.A3(n_918),
.B1(n_919),
.B2(n_921),
.C1(n_936),
.C2(n_933),
.Y(n_1559)
);

NAND3x1_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_903),
.C(n_931),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_R g1561 ( 
.A(n_1545),
.B(n_1541),
.Y(n_1561)
);

AND4x2_ASAP7_75t_L g1562 ( 
.A(n_1543),
.B(n_1533),
.C(n_1541),
.D(n_1538),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1547),
.B(n_1537),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1550),
.A2(n_1536),
.B(n_743),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1551),
.A2(n_738),
.B1(n_743),
.B2(n_729),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1544),
.Y(n_1566)
);

NAND4xp75_ASAP7_75t_L g1567 ( 
.A(n_1555),
.B(n_931),
.C(n_938),
.D(n_889),
.Y(n_1567)
);

NOR3xp33_ASAP7_75t_L g1568 ( 
.A(n_1549),
.B(n_738),
.C(n_903),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1546),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1557),
.B(n_903),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1553),
.B(n_918),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1548),
.B(n_919),
.C(n_921),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1552),
.B(n_1556),
.C(n_1558),
.Y(n_1573)
);

NAND4xp75_ASAP7_75t_L g1574 ( 
.A(n_1558),
.B(n_938),
.C(n_889),
.D(n_944),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1554),
.B(n_921),
.Y(n_1575)
);

NAND4xp25_ASAP7_75t_L g1576 ( 
.A(n_1560),
.B(n_893),
.C(n_921),
.D(n_933),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1569),
.B(n_1559),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1566),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1563),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1573),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1564),
.A2(n_933),
.B1(n_935),
.B2(n_936),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1561),
.B(n_933),
.Y(n_1582)
);

NAND3x1_ASAP7_75t_L g1583 ( 
.A(n_1562),
.B(n_945),
.C(n_938),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1574),
.B(n_935),
.Y(n_1584)
);

XOR2x2_ASAP7_75t_L g1585 ( 
.A(n_1565),
.B(n_893),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_L g1586 ( 
.A(n_1568),
.B(n_936),
.C(n_935),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1571),
.B(n_935),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1575),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1579),
.A2(n_1570),
.B1(n_1572),
.B2(n_1567),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1580),
.B(n_1576),
.C(n_936),
.Y(n_1590)
);

AOI322xp5_ASAP7_75t_L g1591 ( 
.A1(n_1578),
.A2(n_893),
.A3(n_897),
.B1(n_898),
.B2(n_899),
.C1(n_900),
.C2(n_944),
.Y(n_1591)
);

XOR2x2_ASAP7_75t_L g1592 ( 
.A(n_1583),
.B(n_893),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1577),
.A2(n_912),
.B1(n_885),
.B2(n_946),
.C(n_888),
.Y(n_1593)
);

AOI322xp5_ASAP7_75t_L g1594 ( 
.A1(n_1588),
.A2(n_897),
.A3(n_898),
.B1(n_899),
.B2(n_900),
.C1(n_944),
.C2(n_930),
.Y(n_1594)
);

OAI322xp33_ASAP7_75t_L g1595 ( 
.A1(n_1582),
.A2(n_885),
.A3(n_946),
.B1(n_941),
.B2(n_930),
.C1(n_929),
.C2(n_927),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1592),
.Y(n_1596)
);

INVx3_ASAP7_75t_SL g1597 ( 
.A(n_1589),
.Y(n_1597)
);

OAI22x1_ASAP7_75t_L g1598 ( 
.A1(n_1590),
.A2(n_1584),
.B1(n_1587),
.B2(n_1585),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1593),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1595),
.B(n_1586),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_SL g1601 ( 
.A1(n_1596),
.A2(n_1581),
.B(n_1594),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1598),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1600),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1599),
.B(n_1597),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1602),
.A2(n_1591),
.B1(n_729),
.B2(n_721),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1604),
.Y(n_1606)
);

AOI22x1_ASAP7_75t_L g1607 ( 
.A1(n_1603),
.A2(n_729),
.B1(n_721),
.B2(n_941),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_R g1608 ( 
.A1(n_1601),
.A2(n_915),
.B1(n_878),
.B2(n_946),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1606),
.A2(n_1607),
.B(n_1608),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1605),
.A2(n_729),
.B1(n_915),
.B2(n_941),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_885),
.B1(n_876),
.B2(n_930),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1610),
.A2(n_882),
.B1(n_878),
.B2(n_929),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1611),
.A2(n_650),
.B(n_949),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_1612),
.B(n_906),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_882),
.B1(n_929),
.B2(n_927),
.C(n_920),
.Y(n_1615)
);

AOI211xp5_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_882),
.B(n_927),
.C(n_920),
.Y(n_1616)
);


endmodule