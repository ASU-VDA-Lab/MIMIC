module fake_aes_2047_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
BUFx3_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_8), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_6), .B(n_1), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_13), .B(n_0), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_15), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_11), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_19), .B(n_14), .Y(n_23) );
AO31x2_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_21), .A3(n_22), .B(n_14), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_20), .B(n_12), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
NAND2x1_ASAP7_75t_L g27 ( .A(n_26), .B(n_22), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_17), .B1(n_2), .B2(n_5), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_29), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_28), .B(n_25), .Y(n_31) );
XNOR2x1_ASAP7_75t_L g32 ( .A(n_30), .B(n_2), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
INVxp67_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
AOI211x1_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_24), .B(n_10), .C(n_3), .Y(n_36) );
INVxp67_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
NOR2x1_ASAP7_75t_L g39 ( .A(n_36), .B(n_33), .Y(n_39) );
BUFx2_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
INVx2_ASAP7_75t_SL g41 ( .A(n_39), .Y(n_41) );
AOI22xp5_ASAP7_75t_SL g42 ( .A1(n_40), .A2(n_27), .B1(n_35), .B2(n_41), .Y(n_42) );
endmodule