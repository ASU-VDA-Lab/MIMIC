module fake_jpeg_30772_n_499 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_499);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_499;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_9),
.B(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_53),
.B(n_58),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_54),
.B(n_88),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_17),
.B(n_14),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_27),
.B(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_83),
.Y(n_113)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_25),
.B(n_1),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_92),
.Y(n_139)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_23),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_39),
.B(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_99),
.B(n_23),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_45),
.C(n_41),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_54),
.B(n_45),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_37),
.B(n_46),
.C(n_43),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_109),
.B(n_153),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_39),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_118),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_57),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_48),
.B1(n_44),
.B2(n_37),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_143),
.B1(n_66),
.B2(n_78),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_28),
.B(n_50),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_48),
.B1(n_44),
.B2(n_50),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_142),
.B1(n_22),
.B2(n_38),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_70),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_151),
.Y(n_188)
);

AND2x4_ASAP7_75t_SL g135 ( 
.A(n_60),
.B(n_36),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_140),
.Y(n_189)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_30),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_73),
.A2(n_48),
.B1(n_44),
.B2(n_50),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_55),
.A2(n_97),
.B1(n_59),
.B2(n_94),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_64),
.A2(n_41),
.B1(n_48),
.B2(n_44),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_18),
.B1(n_35),
.B2(n_31),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_92),
.B1(n_65),
.B2(n_89),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_154),
.A2(n_159),
.B1(n_163),
.B2(n_167),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_155),
.B(n_162),
.Y(n_229)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_88),
.B1(n_86),
.B2(n_82),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_157),
.B(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_99),
.A2(n_75),
.B1(n_74),
.B2(n_52),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g243 ( 
.A1(n_165),
.A2(n_111),
.B(n_30),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_61),
.B1(n_28),
.B2(n_46),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_100),
.B(n_31),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_168),
.B(n_174),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_90),
.B1(n_46),
.B2(n_43),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_169),
.A2(n_180),
.B1(n_204),
.B2(n_124),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_170),
.A2(n_199),
.B1(n_144),
.B2(n_149),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_22),
.B1(n_38),
.B2(n_35),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_191),
.B1(n_192),
.B2(n_139),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_131),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_173),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_113),
.B(n_43),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_22),
.B1(n_38),
.B2(n_35),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_106),
.B1(n_107),
.B2(n_148),
.Y(n_217)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_185),
.B(n_196),
.Y(n_248)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_119),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_139),
.A2(n_29),
.B1(n_18),
.B2(n_40),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_29),
.B1(n_18),
.B2(n_40),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_202),
.B1(n_130),
.B2(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_138),
.B(n_2),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_127),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_197),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_201),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_127),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_30),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_200),
.B(n_23),
.CI(n_3),
.CON(n_249),
.SN(n_249)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_139),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_124),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_110),
.A2(n_120),
.B1(n_152),
.B2(n_126),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_207),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_140),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_225),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_210),
.A2(n_213),
.B(n_228),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_109),
.B(n_140),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_110),
.B1(n_152),
.B2(n_120),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_196),
.A2(n_107),
.B1(n_145),
.B2(n_106),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_128),
.B(n_148),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_221),
.B(n_226),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_104),
.Y(n_225)
);

NAND2x1_ASAP7_75t_SL g226 ( 
.A(n_169),
.B(n_111),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_104),
.C(n_149),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_247),
.C(n_163),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_144),
.B(n_103),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_134),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_237),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_199),
.A2(n_147),
.B1(n_130),
.B2(n_134),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_232),
.A2(n_235),
.B1(n_243),
.B2(n_167),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_112),
.B1(n_101),
.B2(n_147),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_40),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_40),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_40),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_112),
.C(n_101),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_192),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_267),
.Y(n_297)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_207),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_252),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_168),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_253),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_174),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_254),
.Y(n_312)
);

AO21x2_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_157),
.B(n_237),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_275),
.B(n_216),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_180),
.B1(n_159),
.B2(n_157),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_258),
.A2(n_263),
.B1(n_286),
.B2(n_242),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_155),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_279),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_226),
.A2(n_187),
.B1(n_161),
.B2(n_158),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_266),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_200),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_270),
.Y(n_298)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_164),
.C(n_188),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_197),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_171),
.B1(n_154),
.B2(n_182),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_274),
.A2(n_285),
.B1(n_236),
.B2(n_244),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_205),
.B(n_157),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_203),
.B1(n_183),
.B2(n_185),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_281),
.B1(n_282),
.B2(n_215),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_241),
.B(n_172),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_162),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_173),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_287),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_181),
.B1(n_186),
.B2(n_177),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_178),
.B1(n_175),
.B2(n_179),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_235),
.A2(n_190),
.B1(n_202),
.B2(n_23),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_221),
.B1(n_245),
.B2(n_206),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_231),
.B(n_156),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_213),
.A2(n_156),
.B(n_193),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_249),
.C(n_232),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_206),
.B(n_23),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_259),
.B1(n_275),
.B2(n_286),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_227),
.C(n_247),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_293),
.B(n_259),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_228),
.B(n_248),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_294),
.A2(n_320),
.B(n_288),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_248),
.C(n_222),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

NAND2x1p5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_220),
.Y(n_296)
);

AO22x2_ASAP7_75t_SL g361 ( 
.A1(n_296),
.A2(n_304),
.B1(n_294),
.B2(n_303),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_307),
.A2(n_322),
.B1(n_261),
.B2(n_272),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_309),
.A2(n_268),
.B(n_292),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_249),
.C(n_224),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_315),
.C(n_270),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_236),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_253),
.B(n_233),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_313),
.B(n_314),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_233),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_224),
.C(n_230),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_230),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_317),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_208),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_208),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_324),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_273),
.A2(n_214),
.B(n_244),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_242),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_277),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_2),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_283),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_325),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_3),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_251),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_330),
.A2(n_352),
.B1(n_353),
.B2(n_291),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_345),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_360),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_301),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_333),
.B(n_358),
.Y(n_388)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_334),
.Y(n_371)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_343),
.B(n_360),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_342),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_255),
.B(n_259),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_275),
.B1(n_258),
.B2(n_256),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_348),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_267),
.C(n_255),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_355),
.C(n_356),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_319),
.A2(n_256),
.B1(n_261),
.B2(n_281),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_351),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_299),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_350),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_306),
.B(n_289),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_322),
.A2(n_282),
.B1(n_256),
.B2(n_250),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_256),
.B1(n_284),
.B2(n_269),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_336),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_293),
.C(n_297),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_266),
.C(n_251),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_300),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_292),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_359),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_309),
.A2(n_264),
.B(n_23),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_362),
.A2(n_364),
.B1(n_368),
.B2(n_387),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_330),
.A2(n_304),
.B1(n_296),
.B2(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_353),
.A2(n_304),
.B1(n_296),
.B2(n_302),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_315),
.C(n_310),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_382),
.C(n_386),
.Y(n_397)
);

NOR3xp33_ASAP7_75t_SL g372 ( 
.A(n_338),
.B(n_302),
.C(n_308),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_385),
.C(n_336),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_325),
.Y(n_376)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_305),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_337),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_361),
.A2(n_305),
.B(n_321),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_341),
.C(n_332),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_361),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_351),
.Y(n_410)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_326),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_321),
.B1(n_326),
.B2(n_328),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_338),
.B(n_4),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_389),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_4),
.Y(n_390)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_391),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_404),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_374),
.B(n_344),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_406),
.Y(n_417)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_343),
.B1(n_346),
.B2(n_335),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_401),
.A2(n_407),
.B1(n_357),
.B2(n_378),
.Y(n_430)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_339),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_372),
.B(n_340),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_331),
.B1(n_349),
.B2(n_345),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_413),
.B1(n_415),
.B2(n_375),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_356),
.C(n_337),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_409),
.B(n_382),
.C(n_369),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_410),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_348),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_411),
.Y(n_422)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_386),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_427),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_416),
.A2(n_383),
.B(n_370),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_364),
.B(n_368),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_414),
.A2(n_373),
.B1(n_362),
.B2(n_379),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_426),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_432),
.C(n_397),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_414),
.A2(n_379),
.B1(n_377),
.B2(n_367),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_367),
.B1(n_387),
.B2(n_385),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_413),
.A2(n_388),
.B1(n_334),
.B2(n_375),
.Y(n_428)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_430),
.A2(n_392),
.B1(n_398),
.B2(n_394),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_365),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_401),
.A2(n_365),
.B(n_354),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_407),
.B(n_410),
.C(n_411),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_441),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_397),
.C(n_396),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_448),
.Y(n_453)
);

AO221x1_ASAP7_75t_L g444 ( 
.A1(n_417),
.A2(n_399),
.B1(n_412),
.B2(n_402),
.C(n_400),
.Y(n_444)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_420),
.B(n_403),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_447),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_423),
.A2(n_394),
.B(n_415),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_4),
.C(n_5),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_436),
.Y(n_457)
);

XNOR2x1_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_11),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_433),
.C(n_418),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_452),
.A2(n_427),
.B1(n_424),
.B2(n_426),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_455),
.A2(n_459),
.B1(n_449),
.B2(n_438),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_435),
.B(n_421),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_438),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_461),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_419),
.B1(n_422),
.B2(n_428),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_451),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_432),
.C(n_430),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_466),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_5),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_467),
.B(n_470),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_465),
.B(n_446),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_469),
.Y(n_483)
);

NOR3xp33_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_438),
.C(n_449),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_471),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_464),
.A2(n_5),
.B(n_6),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_460),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_478),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_6),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_477),
.Y(n_487)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

NAND3xp33_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_476),
.C(n_472),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_479),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_463),
.C(n_453),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_485),
.A2(n_6),
.B(n_7),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_480),
.B(n_453),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_489),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_455),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_456),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_492),
.C(n_487),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_493),
.A2(n_484),
.B(n_482),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_486),
.C(n_481),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_495),
.A2(n_7),
.B(n_10),
.Y(n_497)
);

OAI321xp33_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_497),
.A3(n_7),
.B1(n_11),
.B2(n_494),
.C(n_476),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_498),
.B(n_7),
.Y(n_499)
);


endmodule