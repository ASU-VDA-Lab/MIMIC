module fake_jpeg_12008_n_640 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_640);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_640;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_5),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_67),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_76),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_77),
.Y(n_159)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_84),
.Y(n_150)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_87),
.B(n_111),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_88),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_93),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_92),
.Y(n_206)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_96),
.Y(n_207)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_101),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_18),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_9),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_10),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_109),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_112),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_7),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_18),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

INVx5_ASAP7_75t_SL g173 ( 
.A(n_116),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_19),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_40),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_121),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_25),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_25),
.Y(n_124)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_125),
.Y(n_180)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_81),
.B(n_46),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_128),
.B(n_44),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_130),
.B(n_131),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_35),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_134),
.B(n_141),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_137),
.A2(n_208),
.B1(n_47),
.B2(n_57),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_95),
.B(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_21),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_142),
.B(n_154),
.Y(n_245)
);

INVx6_ASAP7_75t_SL g148 ( 
.A(n_67),
.Y(n_148)
);

CKINVDCx12_ASAP7_75t_R g231 ( 
.A(n_148),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_86),
.B(n_46),
.Y(n_154)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_77),
.A2(n_56),
.B1(n_36),
.B2(n_33),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_171),
.A2(n_47),
.B(n_22),
.Y(n_254)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_62),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_182),
.Y(n_269)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_103),
.B(n_42),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_188),
.B(n_203),
.Y(n_271)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_99),
.B(n_42),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_125),
.A2(n_56),
.B1(n_41),
.B2(n_36),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_68),
.Y(n_209)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_214),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_138),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_217),
.B(n_218),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_133),
.B(n_48),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_219),
.A2(n_226),
.B1(n_273),
.B2(n_53),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_220),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_139),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_223),
.B(n_230),
.Y(n_303)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_171),
.B1(n_147),
.B2(n_206),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_227),
.Y(n_309)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_48),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_132),
.B(n_56),
.C(n_60),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_261),
.C(n_159),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_98),
.B1(n_83),
.B2(n_70),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_237),
.A2(n_169),
.B1(n_162),
.B2(n_191),
.Y(n_334)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_43),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_240),
.B(n_243),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_242),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_164),
.B(n_60),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_186),
.A2(n_71),
.B1(n_90),
.B2(n_58),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_249),
.Y(n_295)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_149),
.Y(n_250)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_250),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_167),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_251),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_150),
.B(n_122),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_252),
.B(n_253),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_150),
.B(n_113),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_254),
.A2(n_200),
.B(n_151),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_182),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_258),
.Y(n_294)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_257),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_190),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_165),
.B(n_59),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_268),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_135),
.B(n_166),
.C(n_156),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_264),
.Y(n_335)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_157),
.Y(n_265)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

INVx11_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_152),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_152),
.A2(n_24),
.B(n_44),
.C(n_30),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g342 ( 
.A1(n_270),
.A2(n_155),
.B(n_58),
.Y(n_342)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_146),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_204),
.A2(n_79),
.B1(n_102),
.B2(n_96),
.Y(n_273)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_285),
.Y(n_293)
);

OR2x4_ASAP7_75t_L g277 ( 
.A(n_174),
.B(n_24),
.Y(n_277)
);

AOI22x1_ASAP7_75t_L g328 ( 
.A1(n_277),
.A2(n_45),
.B1(n_53),
.B2(n_162),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_55),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_280),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_175),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_210),
.B(n_30),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_282),
.Y(n_336)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_184),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_184),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_284),
.Y(n_343)
);

OAI32xp33_ASAP7_75t_L g284 ( 
.A1(n_201),
.A2(n_53),
.A3(n_41),
.B1(n_45),
.B2(n_123),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_22),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_298),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_297),
.C(n_300),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_172),
.C(n_159),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_211),
.B(n_57),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_180),
.C(n_196),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_270),
.A2(n_180),
.B1(n_196),
.B2(n_207),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_334),
.B1(n_286),
.B2(n_330),
.Y(n_346)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_229),
.B(n_202),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_304),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_158),
.B1(n_197),
.B2(n_204),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_306),
.A2(n_333),
.B1(n_267),
.B2(n_239),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_235),
.B(n_202),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_312),
.B(n_329),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_319),
.B(n_339),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_216),
.B(n_153),
.C(n_151),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_338),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_158),
.B1(n_197),
.B2(n_153),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_342),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_224),
.B(n_169),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g330 ( 
.A(n_225),
.B(n_275),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_330),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_244),
.B(n_129),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_55),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_345),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_231),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_246),
.B(n_191),
.C(n_178),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_236),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_276),
.B(n_200),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_346),
.A2(n_353),
.B1(n_360),
.B2(n_361),
.Y(n_428)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_343),
.A2(n_319),
.B1(n_333),
.B2(n_336),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_355),
.A2(n_380),
.B(n_332),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_357),
.Y(n_394)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_288),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_322),
.A2(n_251),
.B1(n_213),
.B2(n_214),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_304),
.A2(n_228),
.B1(n_266),
.B2(n_248),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_262),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_362),
.B(n_374),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_257),
.B1(n_259),
.B2(n_237),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_285),
.Y(n_367)
);

A2O1A1O1Ixp25_ASAP7_75t_L g400 ( 
.A1(n_367),
.A2(n_381),
.B(n_316),
.C(n_287),
.D(n_313),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_304),
.A2(n_178),
.B1(n_207),
.B2(n_144),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_286),
.B1(n_317),
.B2(n_292),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_312),
.A2(n_291),
.B1(n_328),
.B2(n_300),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_369),
.A2(n_388),
.B1(n_293),
.B2(n_311),
.Y(n_411)
);

INVx13_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_377),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_264),
.Y(n_374)
);

BUFx12_ASAP7_75t_L g377 ( 
.A(n_309),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_385),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_289),
.B(n_263),
.Y(n_380)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_308),
.B(n_255),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_298),
.B(n_212),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_383),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_212),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_317),
.A2(n_269),
.B1(n_221),
.B2(n_249),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_384),
.A2(n_330),
.B1(n_332),
.B2(n_331),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_327),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_269),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_387),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_297),
.B(n_255),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_293),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_390),
.Y(n_397)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_290),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_307),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_410),
.B1(n_359),
.B2(n_375),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_400),
.B(n_309),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_303),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_402),
.B(n_421),
.C(n_372),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_357),
.A2(n_322),
.B(n_331),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_406),
.A2(n_417),
.B(n_425),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_349),
.B(n_296),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_408),
.B(n_426),
.Y(n_460)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_320),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_412),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_376),
.A2(n_328),
.B1(n_290),
.B2(n_311),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_411),
.A2(n_413),
.B1(n_423),
.B2(n_427),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_363),
.B(n_369),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_350),
.A2(n_344),
.B1(n_301),
.B2(n_292),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_376),
.A2(n_325),
.B(n_335),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_430),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_307),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_350),
.A2(n_344),
.B1(n_301),
.B2(n_299),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_375),
.A2(n_299),
.B(n_295),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_349),
.B(n_295),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_350),
.A2(n_222),
.B1(n_215),
.B2(n_220),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_363),
.B(n_321),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_377),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_347),
.B(n_340),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_434),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_399),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_386),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g492 ( 
.A1(n_435),
.A2(n_451),
.B(n_457),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_423),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_410),
.A2(n_352),
.B1(n_367),
.B2(n_379),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_437),
.A2(n_438),
.B1(n_436),
.B2(n_442),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_428),
.A2(n_406),
.B1(n_394),
.B2(n_418),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_346),
.B(n_354),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_439),
.A2(n_442),
.B(n_446),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_383),
.Y(n_440)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_351),
.B(n_356),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_380),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_450),
.Y(n_473)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_444),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_425),
.A2(n_356),
.B(n_385),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_411),
.A2(n_368),
.B1(n_382),
.B2(n_361),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_449),
.A2(n_393),
.B1(n_407),
.B2(n_413),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_365),
.Y(n_450)
);

NOR2x1_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_389),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_420),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_466),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_455),
.C(n_465),
.Y(n_482)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_454),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_402),
.C(n_412),
.Y(n_455)
);

FAx1_ASAP7_75t_SL g456 ( 
.A(n_395),
.B(n_381),
.CI(n_371),
.CON(n_456),
.SN(n_456)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_462),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_397),
.A2(n_390),
.B(n_366),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_459),
.B(n_396),
.Y(n_484)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_405),
.Y(n_461)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_461),
.Y(n_498)
);

INVx8_ASAP7_75t_L g464 ( 
.A(n_416),
.Y(n_464)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_464),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_340),
.C(n_321),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_391),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_405),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_467),
.Y(n_483)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_468),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_455),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_470),
.B(n_472),
.C(n_474),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_395),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_429),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_401),
.Y(n_475)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_441),
.A2(n_418),
.B1(n_396),
.B2(n_426),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_476),
.A2(n_490),
.B1(n_492),
.B2(n_483),
.Y(n_511)
);

OAI21xp33_ASAP7_75t_L g479 ( 
.A1(n_433),
.A2(n_398),
.B(n_415),
.Y(n_479)
);

HAxp5_ASAP7_75t_SL g520 ( 
.A(n_479),
.B(n_456),
.CON(n_520),
.SN(n_520)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_435),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_430),
.Y(n_485)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_439),
.B(n_407),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_496),
.C(n_497),
.Y(n_514)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_400),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_463),
.C(n_438),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_447),
.A2(n_437),
.B(n_463),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_499),
.A2(n_414),
.B(n_416),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_501),
.A2(n_525),
.B(n_488),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_473),
.B(n_469),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_502),
.B(n_526),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_431),
.Y(n_503)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_503),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_432),
.Y(n_504)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_504),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_505),
.B(n_520),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_471),
.B(n_432),
.Y(n_507)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_478),
.B(n_460),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_508),
.B(n_521),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_435),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_518),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_511),
.A2(n_524),
.B1(n_324),
.B2(n_373),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_466),
.Y(n_515)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_515),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_467),
.C(n_461),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_519),
.C(n_523),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_451),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_470),
.B(n_454),
.C(n_444),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_494),
.B(n_460),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_472),
.B(n_419),
.C(n_449),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_499),
.A2(n_456),
.B1(n_427),
.B2(n_445),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_496),
.B(n_416),
.Y(n_526)
);

XNOR2x2_ASAP7_75t_L g527 ( 
.A(n_484),
.B(n_445),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_489),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_477),
.B(n_464),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_528),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_483),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_529),
.B(n_498),
.Y(n_531)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_531),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_525),
.Y(n_532)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_493),
.Y(n_533)
);

MAJx2_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_552),
.C(n_528),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_535),
.A2(n_501),
.B(n_515),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_524),
.A2(n_497),
.B1(n_487),
.B2(n_481),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_538),
.A2(n_543),
.B1(n_544),
.B2(n_227),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_490),
.B1(n_492),
.B2(n_476),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_539),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g575 ( 
.A(n_540),
.B(n_542),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_513),
.B(n_489),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_530),
.A2(n_487),
.B1(n_495),
.B2(n_491),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_522),
.A2(n_486),
.B1(n_500),
.B2(n_468),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_513),
.B(n_377),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_518),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_519),
.B(n_514),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_554),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_506),
.A2(n_500),
.B1(n_464),
.B2(n_378),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_544),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_358),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_553),
.A2(n_520),
.B1(n_370),
.B2(n_233),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_377),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_516),
.C(n_512),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_557),
.B(n_564),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_548),
.C(n_512),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_559),
.B(n_574),
.Y(n_595)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_560),
.Y(n_585)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_562),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_523),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_535),
.A2(n_522),
.B(n_517),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_568),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_546),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_549),
.B(n_509),
.C(n_527),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_567),
.B(n_573),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_505),
.Y(n_568)
);

OAI321xp33_ASAP7_75t_L g569 ( 
.A1(n_547),
.A2(n_507),
.A3(n_504),
.B1(n_503),
.B2(n_506),
.C(n_517),
.Y(n_569)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_571),
.A2(n_572),
.B1(n_577),
.B2(n_556),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_221),
.C(n_280),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_538),
.B(n_280),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_576),
.A2(n_533),
.B1(n_532),
.B2(n_537),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_555),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_578),
.B(n_594),
.Y(n_604)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_536),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_582),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_536),
.Y(n_582)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_583),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_558),
.A2(n_543),
.B1(n_551),
.B2(n_534),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_586),
.B(n_591),
.Y(n_607)
);

BUFx24_ASAP7_75t_SL g588 ( 
.A(n_563),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_588),
.B(n_568),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_557),
.B(n_540),
.C(n_534),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_SL g608 ( 
.A(n_590),
.B(n_589),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_558),
.A2(n_552),
.B1(n_45),
.B2(n_236),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_570),
.A2(n_577),
.B1(n_565),
.B2(n_562),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_236),
.C(n_175),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_567),
.B(n_560),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_596),
.B(n_598),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_593),
.A2(n_595),
.B(n_584),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_597),
.A2(n_608),
.B(n_3),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_581),
.B(n_566),
.C(n_575),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_579),
.B(n_575),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_599),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_573),
.C(n_571),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_58),
.C(n_6),
.Y(n_616)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_601),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_163),
.C(n_123),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_603),
.B(n_11),
.Y(n_619)
);

AOI221xp5_ASAP7_75t_L g606 ( 
.A1(n_587),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.C(n_3),
.Y(n_606)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_606),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_605),
.B(n_585),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_611),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_609),
.A2(n_590),
.B1(n_580),
.B2(n_578),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_602),
.A2(n_579),
.B1(n_58),
.B2(n_7),
.Y(n_612)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_612),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_0),
.C(n_1),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_4),
.B(n_14),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_617),
.A2(n_619),
.B1(n_620),
.B2(n_13),
.Y(n_627)
);

AOI322xp5_ASAP7_75t_L g623 ( 
.A1(n_615),
.A2(n_607),
.A3(n_599),
.B1(n_604),
.B2(n_600),
.C1(n_598),
.C2(n_606),
.Y(n_623)
);

AO21x1_ASAP7_75t_L g631 ( 
.A1(n_623),
.A2(n_627),
.B(n_614),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_624),
.B(n_625),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_618),
.B(n_15),
.C(n_3),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_15),
.C(n_3),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_626),
.B(n_617),
.C(n_616),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_621),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_628),
.A2(n_631),
.B(n_623),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_629),
.B(n_630),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_622),
.A2(n_613),
.B(n_612),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_SL g635 ( 
.A1(n_634),
.A2(n_632),
.B(n_13),
.C(n_14),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_635),
.A2(n_636),
.B(n_0),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_633),
.A2(n_13),
.B(n_1),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_637),
.A2(n_0),
.B(n_2),
.C(n_615),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_0),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_2),
.C(n_242),
.Y(n_640)
);


endmodule