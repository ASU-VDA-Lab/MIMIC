module fake_jpeg_1924_n_528 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_6),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_57),
.Y(n_108)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_6),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_59),
.Y(n_158)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_13),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_66),
.B(n_72),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_13),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_74),
.B(n_80),
.Y(n_155)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_19),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_83),
.Y(n_109)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_17),
.B(n_5),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_5),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_94),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_35),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_97),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_36),
.B(n_0),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_31),
.B1(n_39),
.B2(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_114),
.A2(n_121),
.B1(n_138),
.B2(n_150),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_27),
.B1(n_40),
.B2(n_37),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_27),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_125),
.B(n_127),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_37),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_56),
.B(n_40),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_129),
.B(n_132),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_45),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g183 ( 
.A(n_130),
.B(n_59),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_56),
.B(n_39),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_48),
.B(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_139),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_34),
.B1(n_45),
.B2(n_41),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_55),
.B(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_76),
.B(n_43),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_143),
.B(n_145),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_96),
.B(n_43),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_82),
.A2(n_41),
.B1(n_16),
.B2(n_33),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_84),
.B(n_36),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_36),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_97),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_58),
.B(n_36),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_162),
.Y(n_222)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_79),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_172),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_60),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_202),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_95),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_177),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_91),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_108),
.B(n_92),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_190),
.Y(n_228)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_183),
.B(n_196),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_63),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_186),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_SL g186 ( 
.A(n_114),
.B(n_54),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_111),
.B(n_68),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_189),
.B(n_192),
.Y(n_242)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_193),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

CKINVDCx12_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_134),
.A2(n_16),
.B1(n_41),
.B2(n_86),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_101),
.B(n_64),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_142),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_152),
.B1(n_124),
.B2(n_144),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_218),
.A2(n_223),
.B1(n_233),
.B2(n_102),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_144),
.B1(n_158),
.B2(n_116),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_172),
.A2(n_156),
.B1(n_124),
.B2(n_152),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_230),
.B1(n_151),
.B2(n_115),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_134),
.B(n_116),
.C(n_117),
.Y(n_229)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_172),
.A2(n_174),
.B1(n_197),
.B2(n_186),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_178),
.A2(n_142),
.B1(n_117),
.B2(n_49),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_195),
.B(n_104),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_173),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_206),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_246),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_242),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_171),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_170),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_170),
.C(n_205),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_258),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_251),
.B(n_253),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_210),
.A2(n_65),
.B1(n_61),
.B2(n_53),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_254),
.A2(n_164),
.B1(n_184),
.B2(n_234),
.Y(n_291)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_161),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_227),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_163),
.C(n_169),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_260),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_221),
.B(n_230),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_275),
.Y(n_301)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_264),
.A2(n_148),
.B1(n_180),
.B2(n_241),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_201),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_268),
.Y(n_303)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_266),
.A2(n_236),
.B1(n_166),
.B2(n_244),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_188),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_221),
.B(n_199),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_213),
.Y(n_307)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

OA22x2_ASAP7_75t_SL g274 ( 
.A1(n_229),
.A2(n_207),
.B1(n_198),
.B2(n_181),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_190),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_103),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_243),
.B(n_226),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_243),
.B(n_219),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_299),
.B(n_304),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_243),
.B1(n_211),
.B2(n_219),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_286),
.A2(n_288),
.B1(n_291),
.B2(n_294),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_243),
.B1(n_211),
.B2(n_167),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_261),
.B(n_237),
.CI(n_235),
.CON(n_289),
.SN(n_289)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_249),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_267),
.A2(n_241),
.B1(n_236),
.B2(n_217),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_248),
.A2(n_165),
.B1(n_234),
.B2(n_237),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_253),
.A2(n_216),
.B1(n_238),
.B2(n_151),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_302),
.B1(n_306),
.B2(n_308),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_235),
.B(n_212),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_267),
.A2(n_276),
.B(n_256),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_216),
.B1(n_212),
.B2(n_217),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_307),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_252),
.A2(n_216),
.B1(n_238),
.B2(n_215),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_248),
.C(n_250),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_316),
.C(n_339),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_310),
.B(n_254),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_279),
.B(n_268),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_311),
.B(n_314),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_312),
.B(n_322),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_296),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_313),
.B(n_331),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_250),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_281),
.B(n_246),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_318),
.B(n_319),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_281),
.B(n_259),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_249),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_337),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_247),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_260),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_270),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_262),
.B1(n_276),
.B2(n_253),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_307),
.B1(n_295),
.B2(n_291),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_335),
.Y(n_350)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_258),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_297),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_308),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_258),
.C(n_265),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_265),
.Y(n_340)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_341),
.Y(n_384)
);

OAI22x1_ASAP7_75t_SL g343 ( 
.A1(n_328),
.A2(n_304),
.B1(n_289),
.B2(n_277),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_343),
.A2(n_364),
.B1(n_365),
.B2(n_371),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_282),
.C(n_278),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_352),
.C(n_370),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_323),
.A2(n_298),
.B1(n_280),
.B2(n_278),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_346),
.A2(n_274),
.B1(n_329),
.B2(n_326),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_307),
.B(n_280),
.Y(n_347)
);

AOI21xp33_ASAP7_75t_L g379 ( 
.A1(n_347),
.A2(n_336),
.B(n_330),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_287),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_348),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_303),
.C(n_300),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_300),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_353),
.Y(n_402)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_287),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_357),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_303),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_366),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_286),
.Y(n_363)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_317),
.A2(n_289),
.B1(n_254),
.B2(n_275),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_317),
.B(n_271),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_271),
.C(n_306),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_213),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_373),
.B(n_331),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_365),
.A2(n_334),
.B1(n_325),
.B2(n_327),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_377),
.A2(n_378),
.B1(n_381),
.B2(n_399),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_334),
.B1(n_325),
.B2(n_327),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_347),
.B(n_353),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_343),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_346),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_360),
.A2(n_330),
.B1(n_329),
.B2(n_320),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_329),
.Y(n_385)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_387),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_389),
.A2(n_363),
.B1(n_355),
.B2(n_367),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_369),
.B(n_273),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_356),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_255),
.C(n_266),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_394),
.C(n_395),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_255),
.C(n_266),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_215),
.C(n_245),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_344),
.C(n_352),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_390),
.C(n_395),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_371),
.A2(n_326),
.B1(n_264),
.B2(n_274),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_354),
.A2(n_274),
.B1(n_238),
.B2(n_236),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_401),
.B1(n_157),
.B2(n_136),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_361),
.A2(n_274),
.B1(n_245),
.B2(n_225),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_416),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_366),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_413),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_391),
.B(n_359),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_409),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_411),
.B(n_414),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_370),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_402),
.A2(n_350),
.B(n_358),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_350),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_362),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_426),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_358),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_429),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_419),
.B(n_168),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_349),
.Y(n_420)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_402),
.A2(n_380),
.B(n_378),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_375),
.B(n_401),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_396),
.Y(n_424)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_424),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_382),
.B1(n_374),
.B2(n_376),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_367),
.C(n_225),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_427),
.A2(n_389),
.B1(n_386),
.B2(n_385),
.Y(n_440)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_383),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_168),
.Y(n_429)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_418),
.C(n_412),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_433),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_403),
.C(n_374),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_377),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_434),
.B(n_439),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_398),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_440),
.A2(n_443),
.B1(n_445),
.B2(n_427),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_382),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_435),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_408),
.A2(n_399),
.B1(n_400),
.B2(n_381),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_425),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_448),
.B(n_449),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_422),
.B(n_104),
.Y(n_449)
);

AOI322xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_50),
.A3(n_52),
.B1(n_105),
.B2(n_119),
.C1(n_35),
.C2(n_148),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_119),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_187),
.Y(n_451)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_451),
.Y(n_463)
);

AOI321xp33_ASAP7_75t_L g452 ( 
.A1(n_407),
.A2(n_141),
.A3(n_90),
.B1(n_126),
.B2(n_115),
.C(n_119),
.Y(n_452)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_406),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_468),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_454),
.A2(n_467),
.B1(n_133),
.B2(n_32),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_437),
.A2(n_423),
.B(n_404),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_456),
.A2(n_465),
.B(n_436),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_416),
.Y(n_458)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g459 ( 
.A(n_446),
.B(n_433),
.CI(n_437),
.CON(n_459),
.SN(n_459)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_460),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_408),
.B1(n_410),
.B2(n_415),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_466),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_445),
.A2(n_429),
.B1(n_157),
.B2(n_136),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_141),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_126),
.Y(n_469)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_71),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_8),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_432),
.C(n_441),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_475),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_458),
.A2(n_444),
.B1(n_447),
.B2(n_451),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_478),
.B1(n_479),
.B2(n_488),
.Y(n_494)
);

AO21x1_ASAP7_75t_L g489 ( 
.A1(n_474),
.A2(n_459),
.B(n_463),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_436),
.C(n_16),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_465),
.A2(n_26),
.B1(n_32),
.B2(n_5),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_32),
.C(n_26),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_480),
.A2(n_468),
.B(n_470),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_457),
.B(n_8),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_481),
.B(n_483),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_8),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_461),
.B(n_7),
.Y(n_485)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_485),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_489),
.A2(n_499),
.B(n_475),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_474),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_498),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_471),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_484),
.A2(n_459),
.B(n_469),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_487),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_501),
.Y(n_509)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_478),
.Y(n_507)
);

AOI21xp33_ASAP7_75t_L g503 ( 
.A1(n_489),
.A2(n_472),
.B(n_476),
.Y(n_503)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_504),
.B(n_506),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_491),
.A2(n_480),
.B(n_479),
.Y(n_506)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_496),
.A2(n_477),
.B(n_7),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_11),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_133),
.C(n_35),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_498),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_514),
.C(n_515),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_493),
.C(n_494),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_508),
.Y(n_516)
);

AOI322xp5_ASAP7_75t_L g521 ( 
.A1(n_516),
.A2(n_510),
.A3(n_518),
.B1(n_493),
.B2(n_517),
.C1(n_497),
.C2(n_35),
.Y(n_521)
);

AOI211x1_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_512),
.B(n_505),
.C(n_492),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_519),
.A2(n_521),
.B(n_4),
.Y(n_523)
);

AOI322xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_11),
.A3(n_4),
.B1(n_9),
.B2(n_3),
.C1(n_1),
.C2(n_2),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_9),
.C(n_11),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_523),
.A2(n_524),
.B(n_520),
.Y(n_525)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_525),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_0),
.C(n_1),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_0),
.B(n_1),
.Y(n_528)
);


endmodule