module fake_aes_10966_n_638 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_638);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_638;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_SL g78 ( .A(n_9), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_31), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_12), .Y(n_80) );
INVx3_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_12), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_75), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_77), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_68), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_15), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_64), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_55), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_71), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_67), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_35), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_48), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_23), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_53), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_33), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_26), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_46), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_32), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_0), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_63), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_19), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_61), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_20), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_44), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_22), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_42), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_51), .Y(n_121) );
BUFx8_ASAP7_75t_L g122 ( .A(n_104), .Y(n_122) );
BUFx8_ASAP7_75t_L g123 ( .A(n_104), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_78), .B(n_1), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_78), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_81), .B(n_2), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_111), .B(n_97), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_111), .B(n_3), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_111), .B(n_30), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_97), .B(n_3), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_108), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_83), .B(n_4), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_82), .B(n_4), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_80), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_90), .B(n_5), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_110), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_110), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_94), .B(n_5), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
NOR2xp33_ASAP7_75t_SL g154 ( .A(n_89), .B(n_36), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_86), .Y(n_155) );
INVx4_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_96), .B(n_6), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_114), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_131), .B(n_80), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_129), .B(n_121), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_130), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_131), .B(n_94), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_156), .B(n_112), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_134), .B(n_121), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_156), .B(n_95), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_130), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_156), .B(n_95), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_131), .B(n_112), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_131), .B(n_117), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_155), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_122), .B(n_116), .Y(n_178) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_143), .B(n_120), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVxp67_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_147), .B(n_116), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_137), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_122), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_144), .Y(n_193) );
INVx4_ASAP7_75t_SL g194 ( .A(n_133), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_124), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_137), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_122), .B(n_88), .Y(n_200) );
INVx5_ASAP7_75t_L g201 ( .A(n_133), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_124), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_149), .B(n_127), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_204), .B(n_134), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_204), .B(n_122), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_192), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_184), .Y(n_211) );
AO22x1_ASAP7_75t_L g212 ( .A1(n_203), .A2(n_133), .B1(n_134), .B2(n_143), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
NOR2x1p5_ASAP7_75t_L g215 ( .A(n_184), .B(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_166), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_177), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_166), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_172), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_192), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_159), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_181), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_202), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_169), .B(n_134), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_163), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_162), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_174), .B(n_168), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_202), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_170), .B(n_123), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
AO22x1_ASAP7_75t_L g235 ( .A1(n_203), .A2(n_133), .B1(n_152), .B2(n_92), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_182), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_158), .B(n_127), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_197), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_173), .B(n_123), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_160), .B(n_123), .Y(n_240) );
BUFx4f_ASAP7_75t_L g241 ( .A(n_169), .Y(n_241) );
INVxp67_ASAP7_75t_L g242 ( .A(n_199), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_160), .B(n_123), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_205), .Y(n_244) );
INVxp67_ASAP7_75t_SL g245 ( .A(n_162), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_162), .Y(n_246) );
INVxp67_ASAP7_75t_SL g247 ( .A(n_179), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_176), .A2(n_152), .B1(n_140), .B2(n_139), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_179), .B(n_152), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_198), .B(n_152), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_189), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_160), .B(n_128), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_205), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_205), .Y(n_255) );
INVx5_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_189), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_179), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_183), .Y(n_261) );
BUFx5_ASAP7_75t_L g262 ( .A(n_188), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_185), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_227), .A2(n_176), .B1(n_136), .B2(n_158), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_236), .B(n_176), .Y(n_265) );
AO32x2_ASAP7_75t_L g266 ( .A1(n_246), .A2(n_198), .A3(n_167), .B1(n_151), .B2(n_153), .Y(n_266) );
NAND2x2_ASAP7_75t_L g267 ( .A(n_215), .B(n_125), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_258), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_206), .Y(n_269) );
INVx8_ASAP7_75t_L g270 ( .A(n_250), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
AND2x6_ASAP7_75t_L g273 ( .A(n_258), .B(n_191), .Y(n_273) );
OR2x6_ASAP7_75t_L g274 ( .A(n_236), .B(n_126), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_224), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_218), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_222), .Y(n_277) );
NAND2xp33_ASAP7_75t_L g278 ( .A(n_262), .B(n_201), .Y(n_278) );
INVx5_ASAP7_75t_L g279 ( .A(n_258), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_206), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_226), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_241), .A2(n_191), .B1(n_103), .B2(n_200), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_210), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_250), .B(n_178), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_232), .Y(n_287) );
INVx5_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g289 ( .A1(n_241), .A2(n_109), .B1(n_138), .B2(n_146), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_228), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_247), .B(n_194), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_241), .B(n_201), .Y(n_292) );
OR2x6_ASAP7_75t_L g293 ( .A(n_250), .B(n_132), .Y(n_293) );
CKINVDCx8_ASAP7_75t_R g294 ( .A(n_218), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_207), .B(n_128), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_230), .A2(n_201), .B1(n_138), .B2(n_136), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_232), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_245), .A2(n_157), .B1(n_154), .B2(n_146), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_213), .Y(n_301) );
AOI221x1_ASAP7_75t_L g302 ( .A1(n_237), .A2(n_150), .B1(n_145), .B2(n_140), .C(n_139), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_213), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_209), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_207), .B(n_194), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_207), .B(n_194), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_214), .Y(n_307) );
INVx5_ASAP7_75t_L g308 ( .A(n_259), .Y(n_308) );
NOR2xp33_ASAP7_75t_SL g309 ( .A(n_211), .B(n_201), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_227), .A2(n_150), .B1(n_145), .B2(n_151), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_216), .A2(n_153), .B1(n_201), .B2(n_84), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_208), .B(n_201), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_252), .B(n_93), .C(n_107), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_209), .Y(n_314) );
OAI22x1_ASAP7_75t_L g315 ( .A1(n_242), .A2(n_93), .B1(n_120), .B2(n_115), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_SL g316 ( .A1(n_312), .A2(n_239), .B(n_233), .C(n_234), .Y(n_316) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_270), .A2(n_257), .B1(n_240), .B2(n_243), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_274), .B(n_253), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_289), .A2(n_216), .B1(n_229), .B2(n_223), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g320 ( .A1(n_270), .A2(n_231), .B1(n_223), .B2(n_229), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
AOI22xp5_ASAP7_75t_SL g322 ( .A1(n_276), .A2(n_235), .B1(n_212), .B2(n_98), .Y(n_322) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_300), .A2(n_225), .B(n_251), .Y(n_323) );
BUFx2_ASAP7_75t_SL g324 ( .A(n_288), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_271), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_288), .B(n_225), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_289), .A2(n_214), .B1(n_244), .B2(n_254), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_310), .B(n_249), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_271), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_301), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g331 ( .A1(n_265), .A2(n_148), .B1(n_235), .B2(n_212), .C1(n_234), .C2(n_238), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_270), .A2(n_238), .B1(n_260), .B2(n_255), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_310), .A2(n_244), .B1(n_254), .B2(n_255), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_264), .A2(n_148), .B1(n_113), .B2(n_115), .C(n_99), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_271), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_267), .A2(n_148), .B1(n_260), .B2(n_102), .C(n_101), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_267), .A2(n_100), .B1(n_105), .B2(n_106), .C(n_118), .Y(n_338) );
AOI21x1_ASAP7_75t_L g339 ( .A1(n_302), .A2(n_193), .B(n_187), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_264), .A2(n_164), .B1(n_165), .B2(n_171), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_282), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_298), .A2(n_164), .B(n_165), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_283), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g344 ( .A1(n_274), .A2(n_259), .B1(n_194), .B2(n_256), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_283), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_307), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_288), .A2(n_262), .B1(n_259), .B2(n_256), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_278), .A2(n_259), .B(n_248), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_339), .A2(n_298), .B(n_314), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_338), .A2(n_274), .B1(n_294), .B2(n_275), .C(n_276), .Y(n_352) );
AOI21xp33_ASAP7_75t_L g353 ( .A1(n_320), .A2(n_315), .B(n_286), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_319), .A2(n_293), .B1(n_286), .B2(n_288), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_339), .A2(n_314), .B(n_304), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_286), .B(n_293), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_328), .A2(n_295), .B1(n_284), .B2(n_271), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
OAI221xp5_ASAP7_75t_SL g359 ( .A1(n_327), .A2(n_293), .B1(n_311), .B2(n_285), .C(n_290), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_328), .A2(n_313), .B1(n_268), .B2(n_303), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g361 ( .A1(n_331), .A2(n_311), .B(n_296), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g362 ( .A1(n_322), .A2(n_309), .B1(n_277), .B2(n_268), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_336), .A2(n_307), .B1(n_272), .B2(n_269), .C(n_280), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_334), .A2(n_287), .B1(n_297), .B2(n_279), .C(n_305), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_318), .B(n_279), .Y(n_366) );
INVxp33_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_330), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_337), .B(n_297), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_337), .B(n_273), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_317), .A2(n_279), .B(n_292), .C(n_171), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_331), .A2(n_279), .B(n_292), .C(n_187), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_346), .A2(n_277), .B1(n_281), .B2(n_308), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_346), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_332), .A2(n_281), .B1(n_277), .B2(n_304), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_341), .B(n_266), .Y(n_377) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_352), .B(n_340), .C(n_333), .D(n_326), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_368), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_351), .B(n_324), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_361), .A2(n_333), .B(n_340), .Y(n_381) );
OA21x2_ASAP7_75t_L g382 ( .A1(n_350), .A2(n_349), .B(n_342), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_361), .A2(n_326), .B1(n_324), .B2(n_323), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g384 ( .A1(n_359), .A2(n_348), .B(n_345), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_353), .A2(n_326), .B1(n_316), .B2(n_323), .C(n_344), .Y(n_385) );
INVx8_ASAP7_75t_L g386 ( .A(n_370), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_368), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_370), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_358), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_364), .A2(n_372), .B(n_357), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_369), .B(n_341), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_369), .B(n_348), .Y(n_393) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_354), .A2(n_343), .B1(n_345), .B2(n_273), .C1(n_305), .C2(n_306), .Y(n_394) );
AOI322xp5_ASAP7_75t_L g395 ( .A1(n_356), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_375), .B(n_329), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_356), .B(n_323), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_353), .B(n_175), .C(n_193), .D(n_180), .Y(n_398) );
AND2x4_ASAP7_75t_SL g399 ( .A(n_375), .B(n_343), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_357), .A2(n_335), .B1(n_329), .B2(n_325), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_363), .B(n_266), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_364), .A2(n_347), .B1(n_335), .B2(n_329), .C(n_325), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_363), .B(n_266), .Y(n_405) );
OAI222xp33_ASAP7_75t_L g406 ( .A1(n_362), .A2(n_325), .B1(n_335), .B2(n_308), .C1(n_266), .C2(n_14), .Y(n_406) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_366), .B(n_175), .C(n_180), .D(n_185), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_377), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_360), .A2(n_306), .B1(n_190), .B2(n_195), .C(n_196), .Y(n_409) );
AOI31xp67_ASAP7_75t_L g410 ( .A1(n_383), .A2(n_371), .A3(n_190), .B(n_350), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_389), .B(n_367), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_408), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_408), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_386), .B(n_377), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_381), .A2(n_376), .B1(n_371), .B2(n_365), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_388), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_408), .B(n_355), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_392), .B(n_355), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_403), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_395), .B(n_373), .C(n_374), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_401), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_386), .B(n_374), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_403), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_392), .B(n_7), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_378), .A2(n_277), .B1(n_273), .B2(n_278), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_390), .B(n_8), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_399), .Y(n_433) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_400), .B(n_291), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_397), .B(n_342), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_393), .B(n_10), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_386), .B(n_13), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_402), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_400), .A2(n_308), .B1(n_299), .B2(n_291), .Y(n_440) );
AND2x4_ASAP7_75t_SL g441 ( .A(n_396), .B(n_308), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_397), .B(n_13), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_380), .B(n_15), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_396), .B(n_16), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_405), .B(n_16), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_391), .B(n_299), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_384), .B(n_385), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_382), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_17), .B1(n_273), .B2(n_196), .C1(n_195), .C2(n_186), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_382), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_404), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_429), .B(n_398), .Y(n_457) );
NOR2xp67_ASAP7_75t_SL g458 ( .A(n_421), .B(n_407), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_430), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_452), .A2(n_394), .B1(n_409), .B2(n_273), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_451), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_426), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_429), .B(n_17), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_414), .B(n_21), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_447), .B(n_24), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_446), .B(n_25), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_447), .B(n_196), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_412), .B(n_196), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_446), .B(n_27), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_435), .B(n_196), .Y(n_471) );
NOR3xp33_ASAP7_75t_SL g472 ( .A(n_425), .B(n_28), .C(n_34), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_413), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_437), .B(n_38), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_430), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_432), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_39), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_437), .B(n_43), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_428), .B(n_45), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_433), .Y(n_480) );
NOR3xp33_ASAP7_75t_SL g481 ( .A(n_425), .B(n_50), .C(n_52), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_432), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_416), .B(n_54), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_442), .B(n_56), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_426), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_415), .Y(n_486) );
NOR3xp33_ASAP7_75t_SL g487 ( .A(n_438), .B(n_57), .C(n_58), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_442), .B(n_59), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_421), .B(n_62), .Y(n_490) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_443), .B(n_186), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_435), .B(n_186), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_436), .B(n_66), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_452), .B(n_186), .C(n_195), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_417), .Y(n_495) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_434), .B(n_69), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_417), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_454), .A2(n_195), .B1(n_256), .B2(n_221), .C(n_220), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_419), .Y(n_499) );
NAND3xp33_ASAP7_75t_SL g500 ( .A(n_431), .B(n_72), .C(n_74), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_423), .B(n_76), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_419), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_426), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_426), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_441), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_439), .B(n_217), .Y(n_506) );
NOR2x1p5_ASAP7_75t_L g507 ( .A(n_427), .B(n_219), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_476), .B(n_450), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_482), .B(n_450), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_456), .B(n_434), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g512 ( .A1(n_494), .A2(n_454), .B(n_445), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_480), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_456), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_459), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_475), .B(n_424), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_473), .B(n_444), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_500), .B(n_449), .C(n_418), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_505), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_459), .B(n_422), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_486), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_488), .B(n_422), .Y(n_523) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_461), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_495), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_497), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_504), .B(n_436), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_499), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_457), .A2(n_431), .B1(n_463), .B2(n_500), .Y(n_529) );
AOI31xp33_ASAP7_75t_L g530 ( .A1(n_460), .A2(n_418), .A3(n_436), .B(n_420), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_472), .A2(n_420), .B(n_448), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_493), .B(n_434), .Y(n_532) );
AOI21xp5_ASAP7_75t_SL g533 ( .A1(n_493), .A2(n_440), .B(n_424), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_502), .B(n_424), .Y(n_534) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_493), .B(n_453), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_496), .A2(n_441), .B(n_448), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_468), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_492), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_491), .B(n_411), .C(n_453), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_462), .B(n_441), .Y(n_540) );
INVx5_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_485), .B(n_410), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_485), .B(n_410), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_472), .A2(n_219), .B(n_220), .C(n_221), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_484), .B(n_248), .C(n_261), .Y(n_545) );
INVxp33_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_503), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g548 ( .A(n_460), .B(n_263), .C(n_256), .D(n_262), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_507), .B(n_263), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_489), .B(n_262), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_471), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_465), .B(n_262), .Y(n_552) );
XOR2x2_ASAP7_75t_L g553 ( .A(n_513), .B(n_496), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_514), .Y(n_554) );
AOI221x1_ASAP7_75t_L g555 ( .A1(n_519), .A2(n_533), .B1(n_512), .B2(n_539), .C(n_545), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_509), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_515), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_514), .B(n_481), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_535), .A2(n_481), .B(n_478), .C(n_474), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_546), .B(n_501), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_520), .B(n_483), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g562 ( .A1(n_530), .A2(n_487), .B1(n_467), .B2(n_466), .C(n_470), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_548), .B(n_477), .Y(n_563) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_530), .A2(n_487), .B1(n_498), .B2(n_479), .C(n_506), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_541), .B(n_464), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_529), .B(n_262), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_522), .B(n_517), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_518), .B(n_537), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_512), .B(n_543), .C(n_542), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_525), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_538), .B(n_551), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_526), .B(n_528), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_541), .B(n_531), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_541), .B(n_536), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_548), .B(n_540), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_524), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_534), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_511), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_549), .Y(n_580) );
OAI221xp5_ASAP7_75t_SL g581 ( .A1(n_532), .A2(n_547), .B1(n_552), .B2(n_550), .C(n_549), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_544), .B(n_508), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_524), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_529), .B(n_512), .C(n_530), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_509), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_514), .B(n_541), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_508), .B(n_510), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_513), .B(n_523), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_509), .Y(n_591) );
XOR2x2_ASAP7_75t_L g592 ( .A(n_513), .B(n_496), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_521), .B(n_513), .Y(n_593) );
XNOR2x1_ASAP7_75t_L g594 ( .A(n_511), .B(n_218), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
NAND2x1_ASAP7_75t_L g596 ( .A(n_533), .B(n_513), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_509), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_509), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_521), .B(n_527), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_554), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_554), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_585), .A2(n_592), .B1(n_553), .B2(n_594), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_553), .A2(n_592), .B1(n_594), .B2(n_576), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g604 ( .A1(n_596), .A2(n_562), .B1(n_560), .B2(n_584), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_593), .B(n_599), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_559), .B(n_558), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_589), .B(n_578), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_555), .A2(n_559), .B(n_558), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_563), .A2(n_574), .B(n_583), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_573), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_590), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_575), .A2(n_574), .B(n_588), .C(n_581), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_575), .B(n_588), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_567), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_602), .A2(n_582), .B1(n_579), .B2(n_564), .C(n_570), .Y(n_615) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_608), .A2(n_580), .B(n_569), .C(n_566), .Y(n_616) );
XNOR2x2_ASAP7_75t_L g617 ( .A(n_603), .B(n_565), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_606), .A2(n_589), .B1(n_568), .B2(n_586), .C(n_556), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_611), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_610), .Y(n_620) );
AO22x1_ASAP7_75t_L g621 ( .A1(n_613), .A2(n_557), .B1(n_561), .B2(n_577), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_606), .A2(n_572), .B1(n_598), .B2(n_597), .C1(n_591), .C2(n_587), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_612), .B(n_571), .C(n_595), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_615), .A2(n_612), .B(n_609), .C(n_601), .Y(n_624) );
OR3x1_ASAP7_75t_L g625 ( .A(n_616), .B(n_604), .C(n_614), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_619), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_618), .B(n_565), .C(n_607), .D(n_605), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_617), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_626), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_628), .B(n_622), .Y(n_630) );
XOR2xp5_ASAP7_75t_L g631 ( .A(n_625), .B(n_623), .Y(n_631) );
INVx4_ASAP7_75t_L g632 ( .A(n_629), .Y(n_632) );
AO22x2_ASAP7_75t_L g633 ( .A1(n_631), .A2(n_620), .B1(n_624), .B2(n_621), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_632), .Y(n_634) );
BUFx2_ASAP7_75t_L g635 ( .A(n_633), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_634), .Y(n_636) );
BUFx3_ASAP7_75t_L g637 ( .A(n_636), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_637), .A2(n_630), .B1(n_635), .B2(n_627), .C(n_600), .Y(n_638) );
endmodule