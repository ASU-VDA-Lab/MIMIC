module fake_jpeg_13935_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_21),
.B1(n_35),
.B2(n_34),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_60),
.B1(n_45),
.B2(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_1),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_46),
.B(n_52),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_7),
.B(n_8),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_48),
.B1(n_45),
.B2(n_52),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_61),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_48),
.B1(n_39),
.B2(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_68),
.B1(n_10),
.B2(n_11),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_78),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_42),
.B(n_39),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_74),
.C(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_83),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_4),
.C(n_5),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_7),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_9),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_9),
.B(n_10),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_93),
.C(n_96),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_91),
.B(n_94),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_8),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_68),
.B1(n_64),
.B2(n_11),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_12),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_15),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_86),
.B1(n_79),
.B2(n_22),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_108),
.B(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_86),
.C(n_20),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_109),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_33),
.B1(n_37),
.B2(n_101),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_106),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_116),
.B(n_92),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_110),
.C(n_105),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_121),
.Y(n_122)
);


endmodule