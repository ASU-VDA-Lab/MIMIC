module fake_aes_8775_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
BUFx6f_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OR2x6_ASAP7_75t_L g5 ( .A(n_2), .B(n_1), .Y(n_5) );
AOI22xp33_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
A2O1A1Ixp33_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_1), .C(n_2), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_6), .B(n_5), .Y(n_9) );
O2A1O1Ixp33_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_6), .B(n_5), .C(n_0), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_5), .Y(n_11) );
OAI211xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_8), .B(n_9), .C(n_3), .Y(n_12) );
NAND4xp25_ASAP7_75t_SL g13 ( .A(n_11), .B(n_9), .C(n_5), .D(n_0), .Y(n_13) );
OR5x1_ASAP7_75t_L g14 ( .A(n_13), .B(n_3), .C(n_5), .D(n_12), .E(n_1), .Y(n_14) );
AOI22xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_3), .B1(n_9), .B2(n_13), .Y(n_15) );
endmodule