module fake_jpeg_30297_n_118 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_32),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_26),
.C(n_16),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_23),
.B1(n_17),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_23),
.B1(n_30),
.B2(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_12),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_3),
.B(n_4),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_64),
.B(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_27),
.B(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_7),
.B1(n_44),
.B2(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_59),
.B1(n_61),
.B2(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_79),
.B1(n_55),
.B2(n_50),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_75),
.B1(n_55),
.B2(n_56),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_30),
.C(n_6),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_79),
.C(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_76),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_7),
.B1(n_44),
.B2(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_44),
.A3(n_54),
.B1(n_46),
.B2(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_56),
.C(n_50),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_67),
.C(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_66),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_55),
.B1(n_50),
.B2(n_56),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_92),
.B1(n_80),
.B2(n_76),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_97),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_99),
.B1(n_69),
.B2(n_89),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_78),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_85),
.B1(n_88),
.B2(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_93),
.C(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_96),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_89),
.B(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_106),
.B(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_110),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_113),
.B(n_115),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_102),
.Y(n_118)
);


endmodule