module fake_jpeg_21176_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_29),
.B1(n_18),
.B2(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_63),
.B(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_36),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_75),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_24),
.B1(n_32),
.B2(n_16),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_20),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_39),
.B(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

NOR4xp25_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_17),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_39),
.B1(n_35),
.B2(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_43),
.B1(n_47),
.B2(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_25),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_58),
.B1(n_76),
.B2(n_68),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_101),
.B(n_75),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_94),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_59),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_59),
.B1(n_79),
.B2(n_83),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_55),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_30),
.B1(n_23),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_74),
.B1(n_72),
.B2(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_109),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_122),
.B(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_121),
.B1(n_125),
.B2(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_134),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_82),
.B1(n_58),
.B2(n_62),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_110),
.B1(n_95),
.B2(n_105),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_57),
.B1(n_63),
.B2(n_30),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_77),
.C(n_61),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_128),
.C(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_57),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_132),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_20),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_23),
.B1(n_30),
.B2(n_26),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_133),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_133),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_143),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_89),
.B(n_101),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_95),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_134),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_101),
.B1(n_86),
.B2(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_154),
.B1(n_155),
.B2(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_93),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_116),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_103),
.B1(n_108),
.B2(n_97),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_87),
.B1(n_107),
.B2(n_23),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_87),
.B(n_4),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_132),
.B(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_11),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_174),
.B(n_148),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_126),
.C(n_116),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_175),
.C(n_135),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_146),
.B1(n_139),
.B2(n_138),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_166),
.B(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_120),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_141),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_20),
.B1(n_77),
.B2(n_61),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_176),
.B1(n_156),
.B2(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_154),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_136),
.C(n_149),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_178),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_135),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_181),
.C(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_138),
.B1(n_148),
.B2(n_147),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_168),
.B(n_170),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_147),
.C(n_61),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_7),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.C(n_163),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_12),
.C(n_14),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_190),
.A2(n_169),
.B1(n_165),
.B2(n_162),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_177),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_170),
.B1(n_171),
.B2(n_166),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_158),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_192),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_196),
.Y(n_212)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_188),
.C(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_209),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_181),
.B(n_189),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_213),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_191),
.B1(n_193),
.B2(n_198),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_210),
.B1(n_207),
.B2(n_208),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_14),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_214),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_191),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_220),
.B(n_222),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_15),
.B(n_8),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_219),
.C(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_214),
.A3(n_213),
.B1(n_9),
.B2(n_10),
.C1(n_8),
.C2(n_7),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_224),
.B(n_227),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_8),
.B(n_9),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_9),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_10),
.Y(n_231)
);


endmodule