module fake_ariane_1233_n_74 (n_8, n_7, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_74);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_74;

wire n_66;
wire n_56;
wire n_60;
wire n_24;
wire n_22;
wire n_71;
wire n_43;
wire n_49;
wire n_27;
wire n_48;
wire n_29;
wire n_64;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_62;
wire n_47;
wire n_32;
wire n_28;
wire n_37;
wire n_58;
wire n_65;
wire n_51;
wire n_67;
wire n_45;
wire n_34;
wire n_69;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_68;
wire n_73;
wire n_72;
wire n_33;
wire n_44;
wire n_40;
wire n_39;
wire n_30;
wire n_63;
wire n_42;
wire n_59;
wire n_57;
wire n_31;
wire n_53;
wire n_70;
wire n_23;
wire n_61;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx6p67_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_13),
.B(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_4),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_15),
.Y(n_46)
);

AOI21x1_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_27),
.B(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

O2A1O1Ixp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_26),
.B(n_22),
.C(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_38),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_59),
.B(n_55),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_SL g65 ( 
.A(n_64),
.B(n_61),
.C(n_46),
.Y(n_65)
);

OAI211xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_44),
.B(n_62),
.C(n_58),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_24),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.C(n_47),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_28),
.B1(n_31),
.B2(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_31),
.B(n_28),
.Y(n_73)
);

OR2x6_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);


endmodule