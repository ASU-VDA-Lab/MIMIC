module fake_jpeg_32064_n_146 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_67),
.Y(n_73)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_51),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_79),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_64),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_49),
.Y(n_88)
);

NAND2x1p5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_58),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_60),
.B(n_69),
.Y(n_85)
);

NOR2x1p5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_55),
.B1(n_51),
.B2(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_93),
.B1(n_100),
.B2(n_86),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_95),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_69),
.B(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_54),
.B1(n_56),
.B2(n_53),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_61),
.B1(n_52),
.B2(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_99),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_24),
.B1(n_42),
.B2(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_1),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_80),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_110),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_7),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_8),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_9),
.C(n_11),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_16),
.C(n_18),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_9),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_45),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_14),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_25),
.B(n_27),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_15),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_29),
.C(n_30),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_128),
.A3(n_35),
.B1(n_36),
.B2(n_37),
.C1(n_38),
.C2(n_34),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_102),
.B1(n_109),
.B2(n_101),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_127),
.B(n_114),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_20),
.B(n_23),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_32),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_115),
.C(n_129),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_109),
.B1(n_104),
.B2(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_133),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_134),
.B(n_135),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_115),
.B1(n_124),
.B2(n_125),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_122),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_133),
.C(n_138),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_139),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_130),
.Y(n_146)
);


endmodule