module real_jpeg_18690_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_1),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_1),
.B(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_3),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_3),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_4),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_6),
.B(n_105),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_6),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_6),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_6),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_6),
.B(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_6),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_6),
.B(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_6),
.B(n_512),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_7),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_7),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_7),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_7),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_7),
.B(n_220),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_8),
.Y(n_102)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_8),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g458 ( 
.A(n_8),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_9),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_9),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_9),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_9),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_9),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_9),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_9),
.A2(n_10),
.B1(n_288),
.B2(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_10),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_10),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g307 ( 
.A(n_10),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_10),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_10),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_10),
.B(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_11),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_12),
.B(n_121),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_12),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_12),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_12),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_12),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_12),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_12),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_12),
.B(n_458),
.Y(n_457)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_13),
.Y(n_321)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_14),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_14),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_14),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_15),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_15),
.B(n_89),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_15),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_15),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_15),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_15),
.B(n_425),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_15),
.B(n_509),
.Y(n_508)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_16),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g463 ( 
.A(n_16),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_16),
.Y(n_497)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_17),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_260),
.B(n_529),
.C(n_536),
.D(n_538),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_230),
.C(n_250),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_183),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_26),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_148),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_27),
.B(n_148),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_110),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_28),
.B(n_111),
.C(n_124),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_78),
.C(n_93),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_30),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_49),
.C(n_63),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_31),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_43),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_33),
.A2(n_41),
.B1(n_114),
.B2(n_118),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_33),
.B(n_42),
.C(n_43),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_33),
.B(n_307),
.C(n_309),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_33),
.A2(n_41),
.B1(n_307),
.B2(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_35),
.Y(n_350)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_36),
.Y(n_483)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_96),
.C(n_100),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_37),
.A2(n_42),
.B1(n_100),
.B2(n_101),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_37),
.B(n_219),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_37),
.B(n_359),
.Y(n_422)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_41),
.B(n_114),
.C(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_44),
.B(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_46),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_47),
.Y(n_347)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_49),
.B(n_63),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_60),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_169)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_53),
.Y(n_310)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_53),
.Y(n_481)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_60),
.A2(n_61),
.B1(n_114),
.B2(n_118),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_61),
.B(n_114),
.C(n_295),
.Y(n_352)
);

XNOR2x1_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_72),
.C(n_76),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_64),
.B(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_64),
.B(n_138),
.C(n_225),
.Y(n_253)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_72),
.A2(n_77),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_75),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_77),
.B(n_138),
.C(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_93),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_88),
.B2(n_92),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_84),
.C(n_88),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_172),
.C(n_176),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_82),
.B(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_87),
.Y(n_283)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_88),
.A2(n_92),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_88),
.B(n_226),
.C(n_256),
.Y(n_537)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_106),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g180 ( 
.A1(n_94),
.A2(n_95),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_96),
.A2(n_225),
.B1(n_226),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_96),
.Y(n_256)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_100),
.B(n_159),
.C(n_163),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_100),
.A2(n_101),
.B1(n_163),
.B2(n_164),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_100),
.B(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_101),
.B(n_429),
.Y(n_465)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_102),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_102),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_103),
.A2(n_253),
.B(n_537),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_105),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_107),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_171),
.C(n_177),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_107),
.A2(n_108),
.B1(n_177),
.B2(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_107),
.B(n_141),
.C(n_144),
.Y(n_235)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_124),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_122),
.C(n_123),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_114),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_118),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_118),
.B(n_134),
.C(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_139),
.B2(n_140),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_127),
.B(n_128),
.C(n_139),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_129),
.Y(n_244)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_134),
.A2(n_138),
.B1(n_225),
.B2(n_226),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_134),
.A2(n_138),
.B1(n_199),
.B2(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_137),
.Y(n_308)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_151),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_170),
.C(n_180),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_155),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_168),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_156),
.B(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_158),
.B(n_168),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_160),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_160),
.B(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_163),
.A2(n_164),
.B1(n_302),
.B2(n_303),
.Y(n_326)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_164),
.B(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_165),
.Y(n_318)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_180),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

OR2x6_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_184),
.B(n_186),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_193),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_187),
.B(n_190),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_193),
.B(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_206),
.C(n_211),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_194),
.A2(n_195),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_203),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_196),
.B(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_198),
.A2(n_203),
.B1(n_204),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_198),
.Y(n_387)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_199),
.Y(n_342)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_399)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_222),
.C(n_225),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_213),
.A2(n_214),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_215),
.A2(n_219),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_215),
.Y(n_358)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_216),
.Y(n_431)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_218),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_219),
.Y(n_359)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_221),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_224),
.Y(n_427)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_227),
.Y(n_379)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g530 ( 
.A1(n_231),
.A2(n_251),
.B(n_531),
.C(n_534),
.D(n_535),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_249),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_232),
.B(n_249),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_235),
.C(n_248),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_247),
.B2(n_248),
.Y(n_234)
);

CKINVDCx12_ASAP7_75t_R g247 ( 
.A(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_243),
.C(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_240),
.Y(n_245)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_252),
.B(n_259),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_252),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.CI(n_258),
.CON(n_252),
.SN(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

NAND2x1_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_412),
.Y(n_260)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_389),
.B(n_405),
.C(n_406),
.D(n_411),
.Y(n_261)
);

OAI21x1_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_365),
.B(n_388),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_336),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g528 ( 
.A(n_264),
.B(n_336),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_297),
.C(n_322),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_265),
.B(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_277),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_266),
.B(n_278),
.C(n_294),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.C(n_272),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_267),
.B(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_268),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_420)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_294),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_284),
.B(n_287),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_287),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_297),
.A2(n_298),
.B1(n_322),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_311),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_305),
.B2(n_306),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_300),
.B(n_306),
.C(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_307),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_316),
.C(n_319),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.C(n_327),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_323),
.B(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_327),
.Y(n_418)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.C(n_334),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_328),
.B(n_334),
.Y(n_470)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_331),
.B(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_354),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_355),
.C(n_364),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_353),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_352),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_348),
.B1(n_349),
.B2(n_351),
.Y(n_344)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_345),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_345),
.A2(n_349),
.B(n_352),
.C(n_381),
.Y(n_380)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_369),
.C(n_370),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_364),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_362),
.C(n_363),
.Y(n_374)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_361),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_365),
.B(n_528),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_367),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_391),
.C(n_392),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_384),
.B2(n_385),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_375)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_395),
.C(n_396),
.Y(n_394)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_385),
.Y(n_392)
);

NAND4xp25_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_406),
.C(n_413),
.D(n_527),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_393),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_397),
.Y(n_393)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_394),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_401),
.B1(n_403),
.B2(n_404),
.Y(n_397)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_398),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_399),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_401),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_403),
.C(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_409),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_435),
.B(n_526),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_432),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_415),
.B(n_432),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.C(n_421),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_416),
.A2(n_417),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_419),
.B(n_421),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.C(n_428),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_422),
.A2(n_423),
.B1(n_424),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_422),
.Y(n_473)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_428),
.B(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_520),
.B(n_525),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_474),
.B(n_519),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_466),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_438),
.B(n_466),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_455),
.C(n_464),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_439),
.A2(n_440),
.B1(n_485),
.B2(n_487),
.Y(n_484)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_450),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_448),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_448),
.C(n_450),
.Y(n_468)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_455),
.A2(n_464),
.B1(n_465),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_455),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_456),
.A2(n_457),
.B1(n_459),
.B2(n_460),
.Y(n_477)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_468),
.B(n_469),
.C(n_471),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_488),
.B(n_518),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_484),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_476),
.B(n_484),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.C(n_482),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_501),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_482),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_485),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_489),
.A2(n_503),
.B(n_517),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_500),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_490),
.B(n_500),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_498),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_498),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_507),
.B(n_516),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_505),
.B(n_506),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_511),
.Y(n_507)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_521),
.B(n_522),
.Y(n_525)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_537),
.Y(n_536)
);


endmodule