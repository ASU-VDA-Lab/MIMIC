module fake_netlist_6_4873_n_20644 (n_5643, n_2542, n_1671, n_2817, n_801, n_4452, n_2576, n_5172, n_4649, n_1674, n_5315, n_741, n_1351, n_5254, n_1212, n_208, n_5362, n_4251, n_2157, n_5019, n_2332, n_3849, n_578, n_5138, n_4388, n_4395, n_1061, n_3089, n_783, n_5653, n_4978, n_5409, n_5301, n_188, n_1854, n_3088, n_3257, n_1342, n_4829, n_5393, n_1387, n_3222, n_677, n_4699, n_1151, n_4686, n_2317, n_5524, n_442, n_5345, n_1975, n_1930, n_3706, n_5818, n_2179, n_5963, n_5055, n_1547, n_3376, n_4868, n_893, n_3801, n_5267, n_4249, n_5950, n_1192, n_3564, n_1844, n_1555, n_5548, n_5057, n_3030, n_830, n_65, n_5838, n_5725, n_447, n_2838, n_5229, n_5325, n_3427, n_852, n_5101, n_2628, n_3071, n_2926, n_1078, n_544, n_5900, n_4273, n_5545, n_35, n_2321, n_2019, n_5102, n_3345, n_2074, n_2919, n_4501, n_2129, n_4724, n_945, n_5598, n_4997, n_2399, n_4843, n_1232, n_4696, n_4347, n_5259, n_5819, n_2480, n_3877, n_3929, n_3048, n_1455, n_5279, n_2786, n_5894, n_5930, n_5239, n_567, n_1781, n_1971, n_5354, n_5332, n_2004, n_1106, n_4814, n_953, n_3979, n_5908, n_3077, n_2873, n_3452, n_3107, n_155, n_4956, n_454, n_1421, n_3664, n_1936, n_5337, n_5129, n_5420, n_1660, n_5070, n_3047, n_4414, n_112, n_713, n_1400, n_2625, n_4646, n_2843, n_3760, n_6015, n_48, n_1560, n_4262, n_734, n_1088, n_1894, n_3347, n_5136, n_907, n_6, n_5638, n_4110, n_1658, n_4950, n_4729, n_4268, n_1967, n_3999, n_3928, n_2613, n_3535, n_4751, n_44, n_2708, n_1648, n_5151, n_1911, n_2011, n_5684, n_5729, n_281, n_564, n_5680, n_279, n_686, n_4102, n_1641, n_3871, n_2735, n_4662, n_4671, n_3959, n_2268, n_1367, n_5504, n_1336, n_5522, n_5828, n_4314, n_2080, n_323, n_5099, n_1381, n_331, n_1699, n_2093, n_4296, n_102, n_2770, n_608, n_2101, n_4507, n_32, n_5902, n_512, n_3484, n_4677, n_792, n_5063, n_1328, n_2917, n_2616, n_5275, n_5306, n_3923, n_3900, n_3488, n_939, n_2811, n_3732, n_2832, n_4226, n_5493, n_1762, n_1910, n_1075, n_3980, n_2998, n_5346, n_4366, n_3446, n_5252, n_5309, n_237, n_1895, n_4294, n_4698, n_4445, n_4810, n_3859, n_2692, n_175, n_3914, n_4456, n_3397, n_3575, n_2469, n_3927, n_5452, n_3888, n_764, n_5476, n_2764, n_2895, n_733, n_2922, n_3882, n_4856, n_3492, n_4369, n_30, n_2068, n_4331, n_4972, n_1290, n_4993, n_5536, n_2072, n_1354, n_586, n_423, n_4375, n_1701, n_6055, n_2678, n_3935, n_5130, n_4291, n_88, n_5532, n_5897, n_1726, n_4613, n_2434, n_2878, n_3012, n_3875, n_5609, n_1167, n_2428, n_4717, n_4877, n_3247, n_871, n_5922, n_210, n_2641, n_5658, n_4731, n_3052, n_178, n_355, n_5046, n_2749, n_3298, n_2254, n_5058, n_1926, n_3273, n_4467, n_1747, n_195, n_5667, n_780, n_2624, n_5865, n_2350, n_5042, n_5305, n_4681, n_4072, n_4752, n_4220, n_835, n_928, n_5281, n_2092, n_1654, n_1750, n_1462, n_2514, n_604, n_5314, n_1588, n_3942, n_3997, n_26, n_2468, n_4381, n_5144, n_515, n_2096, n_3968, n_4466, n_4418, n_3434, n_4510, n_5795, n_4473, n_6043, n_5552, n_5226, n_514, n_687, n_890, n_5457, n_2812, n_190, n_4518, n_1709, n_2393, n_2657, n_5291, n_2921, n_2136, n_2409, n_2252, n_3237, n_949, n_3500, n_3834, n_4589, n_2075, n_2972, n_3542, n_91, n_2763, n_2762, n_3192, n_760, n_1546, n_4394, n_2279, n_161, n_6010, n_1296, n_3352, n_3073, n_5343, n_2150, n_1294, n_3696, n_1420, n_4082, n_595, n_1779, n_524, n_4921, n_1858, n_4329, n_5135, n_3021, n_2558, n_1164, n_4697, n_4288, n_4289, n_3763, n_2712, n_5529, n_3733, n_6042, n_1487, n_3614, n_874, n_382, n_5183, n_2145, n_898, n_4964, n_5957, n_4228, n_3423, n_925, n_1932, n_1101, n_15, n_4636, n_4322, n_3644, n_1249, n_4946, n_2706, n_4767, n_4287, n_2693, n_4137, n_1127, n_1512, n_1451, n_320, n_639, n_963, n_2767, n_4576, n_5929, n_4615, n_5787, n_1139, n_3179, n_1018, n_3400, n_1521, n_1366, n_4000, n_5445, n_2897, n_4389, n_3970, n_5342, n_5501, n_4345, n_996, n_532, n_173, n_1376, n_413, n_4664, n_2170, n_4156, n_948, n_6033, n_977, n_536, n_3158, n_1788, n_4873, n_2643, n_5748, n_3782, n_1835, n_3470, n_5076, n_581, n_5870, n_4713, n_4098, n_5026, n_4476, n_432, n_3700, n_4995, n_3166, n_3104, n_3435, n_842, n_5636, n_2239, n_4310, n_1432, n_5212, n_989, n_2689, n_1473, n_5286, n_2191, n_1246, n_4528, n_5811, n_899, n_1035, n_4914, n_4939, n_499, n_1426, n_3418, n_705, n_11, n_1004, n_1529, n_5530, n_2473, n_5397, n_4634, n_2069, n_2362, n_4096, n_2539, n_2698, n_4123, n_5595, n_3119, n_5427, n_3735, n_2297, n_4379, n_486, n_5388, n_4718, n_1448, n_5901, n_5962, n_3631, n_5599, n_648, n_2445, n_5324, n_2057, n_2103, n_3770, n_2772, n_4440, n_4402, n_927, n_5052, n_4541, n_5009, n_4872, n_929, n_4551, n_2857, n_5326, n_1183, n_4627, n_4079, n_2494, n_5300, n_3342, n_998, n_5035, n_717, n_1383, n_3390, n_3656, n_1424, n_1000, n_3025, n_2137, n_1626, n_1507, n_2482, n_3810, n_552, n_4798, n_2532, n_1388, n_3006, n_216, n_912, n_5010, n_2296, n_3633, n_5352, n_5089, n_2849, n_1201, n_1398, n_884, n_5394, n_4592, n_1395, n_2199, n_2661, n_731, n_5359, n_1955, n_931, n_474, n_312, n_1791, n_66, n_958, n_5137, n_100, n_3331, n_5104, n_1897, n_2064, n_5741, n_2773, n_5405, n_5288, n_589, n_3606, n_1310, n_819, n_1334, n_3591, n_2788, n_964, n_4756, n_2797, n_4746, n_124, n_3892, n_4970, n_4069, n_211, n_2748, n_5194, n_1834, n_2331, n_2292, n_3441, n_3534, n_5952, n_3964, n_2416, n_311, n_5947, n_1877, n_3944, n_1939, n_2030, n_1769, n_5985, n_556, n_2209, n_3605, n_1602, n_4633, n_3306, n_276, n_3026, n_221, n_4584, n_3090, n_5232, n_3724, n_4276, n_5116, n_2990, n_3847, n_1773, n_5001, n_2552, n_1053, n_5176, n_4428, n_1533, n_3323, n_4, n_266, n_2274, n_5761, n_518, n_4618, n_4679, n_1745, n_914, n_3479, n_4496, n_317, n_4805, n_1679, n_90, n_3454, n_2160, n_5760, n_2146, n_2131, n_488, n_5472, n_3547, n_5679, n_2575, n_5100, n_5973, n_4410, n_1933, n_1179, n_324, n_3816, n_4807, n_4411, n_3214, n_1243, n_301, n_2928, n_5166, n_1917, n_1580, n_2822, n_36, n_4180, n_1281, n_3109, n_3354, n_2572, n_1520, n_3126, n_3663, n_2863, n_1419, n_3299, n_5688, n_351, n_5740, n_259, n_1731, n_5820, n_5648, n_2135, n_5745, n_4707, n_1645, n_1832, n_4676, n_5180, n_858, n_2049, n_5182, n_956, n_5534, n_663, n_4880, n_3566, n_2781, n_4126, n_410, n_2829, n_1696, n_3845, n_1594, n_664, n_1869, n_3804, n_4207, n_5196, n_2016, n_5171, n_4470, n_580, n_4813, n_5542, n_1030, n_3901, n_1937, n_465, n_1790, n_5261, n_4014, n_4704, n_341, n_1744, n_828, n_2142, n_4252, n_607, n_4028, n_2448, n_5949, n_4048, n_4596, n_4444, n_5255, n_3756, n_3406, n_820, n_951, n_952, n_3919, n_2263, n_5185, n_974, n_4952, n_2656, n_5023, n_2375, n_5906, n_1934, n_628, n_5660, n_1434, n_1573, n_3981, n_3973, n_2756, n_5334, n_6024, n_807, n_4761, n_1275, n_2884, n_485, n_67, n_1510, n_5783, n_3120, n_5821, n_3797, n_238, n_2024, n_1595, n_4770, n_202, n_1749, n_3474, n_2549, n_4690, n_1669, n_1024, n_3864, n_5556, n_4932, n_5456, n_248, n_2302, n_1667, n_1037, n_5143, n_3592, n_468, n_5500, n_4230, n_2637, n_1639, n_183, n_3967, n_3195, n_466, n_2526, n_4274, n_5215, n_3277, n_2548, n_5386, n_991, n_4189, n_3817, n_340, n_1108, n_3659, n_2559, n_2177, n_39, n_2595, n_5003, n_4827, n_1601, n_1960, n_2694, n_3648, n_1686, n_6059, n_3042, n_6065, n_5094, n_4610, n_4472, n_5433, n_6075, n_3228, n_3657, n_96, n_3081, n_1430, n_1316, n_1287, n_5618, n_1586, n_2264, n_3464, n_380, n_3723, n_1190, n_397, n_4380, n_5978, n_4990, n_4996, n_5247, n_4398, n_2498, n_4515, n_1891, n_5031, n_1213, n_6006, n_2235, n_4193, n_3570, n_5082, n_1673, n_5338, n_3828, n_172, n_2392, n_3424, n_4131, n_239, n_97, n_2298, n_2326, n_1539, n_490, n_3594, n_5689, n_1043, n_4090, n_4165, n_2305, n_2120, n_80, n_4626, n_6048, n_4144, n_2964, n_352, n_2169, n_3485, n_4077, n_5931, n_2371, n_1361, n_662, n_3262, n_4008, n_3356, n_5221, n_5641, n_1642, n_3210, n_937, n_4689, n_1682, n_4547, n_5731, n_3329, n_330, n_3826, n_4905, n_1406, n_4601, n_962, n_3647, n_3681, n_1883, n_4300, n_1288, n_1186, n_4623, n_5007, n_3320, n_2518, n_5883, n_5754, n_3988, n_1720, n_3476, n_4842, n_204, n_482, n_5629, n_3439, n_4135, n_2688, n_394, n_1845, n_1489, n_942, n_2798, n_2852, n_1524, n_1964, n_1920, n_2753, n_1496, n_3292, n_2007, n_2039, n_5434, n_5934, n_1225, n_1544, n_1485, n_1846, n_3437, n_4111, n_533, n_3712, n_4608, n_879, n_2310, n_2506, n_4859, n_94, n_2626, n_5880, n_1567, n_4037, n_3562, n_5852, n_2973, n_5218, n_41, n_3665, n_273, n_3007, n_3528, n_5960, n_4571, n_3698, n_5358, n_3355, n_2454, n_2114, n_3174, n_5321, n_1066, n_1948, n_157, n_4215, n_2154, n_6073, n_1484, n_5290, n_4185, n_3752, n_2283, n_5145, n_4219, n_1229, n_1373, n_3958, n_3985, n_2427, n_4196, n_1447, n_4774, n_2056, n_5210, n_4242, n_5109, n_3389, n_4232, n_4190, n_4902, n_3000, n_5149, n_5571, n_2680, n_1047, n_3375, n_3899, n_1385, n_3713, n_1931, n_502, n_2668, n_1257, n_3197, n_4987, n_2128, n_5512, n_4736, n_2398, n_1725, n_3743, n_834, n_5033, n_2695, n_4035, n_3818, n_3124, n_1741, n_1002, n_1949, n_3759, n_545, n_2671, n_4516, n_2715, n_1804, n_251, n_2508, n_3511, n_2054, n_6025, n_1337, n_1477, n_2614, n_4492, n_2833, n_2758, n_5607, n_3694, n_2937, n_4789, n_5999, n_4376, n_1001, n_2241, n_4708, n_4657, n_1690, n_5341, n_1191, n_1076, n_4512, n_1378, n_855, n_1377, n_695, n_4081, n_1542, n_4542, n_4462, n_1716, n_278, n_4931, n_4536, n_5562, n_3303, n_978, n_4324, n_384, n_1976, n_4382, n_2905, n_1291, n_749, n_1824, n_3954, n_5911, n_2122, n_5622, n_2140, n_3503, n_3160, n_1065, n_5577, n_1255, n_568, n_5124, n_143, n_3951, n_823, n_1074, n_698, n_3569, n_739, n_3874, n_2528, n_5123, n_4639, n_5413, n_1338, n_1097, n_3027, n_781, n_4083, n_1810, n_182, n_5915, n_573, n_1583, n_4480, n_1730, n_2295, n_2746, n_389, n_814, n_5779, n_1643, n_2020, n_4171, n_3652, n_222, n_4023, n_1105, n_721, n_1461, n_742, n_691, n_3617, n_2076, n_6019, n_3567, n_377, n_1598, n_4344, n_2935, n_4705, n_4046, n_3807, n_918, n_1114, n_56, n_763, n_4027, n_3154, n_1227, n_2485, n_3898, n_3520, n_191, n_6036, n_4391, n_946, n_1303, n_4095, n_2881, n_1116, n_1570, n_1702, n_1219, n_3551, n_4947, n_3064, n_1780, n_3897, n_1689, n_8, n_5591, n_3372, n_1944, n_1347, n_795, n_1221, n_6013, n_1245, n_3215, n_448, n_3853, n_4740, n_4631, n_1561, n_1112, n_5518, n_2081, n_2168, n_5068, n_234, n_5847, n_6049, n_1460, n_911, n_82, n_27, n_5159, n_2862, n_472, n_2615, n_4068, n_4625, n_2474, n_3703, n_2437, n_2444, n_25, n_3962, n_2743, n_4766, n_4863, n_2267, n_3035, n_668, n_4166, n_1821, n_1058, n_3378, n_3745, n_3362, n_4744, n_103, n_4188, n_5357, n_2934, n_3667, n_3523, n_2222, n_712, n_3176, n_5541, n_5568, n_31, n_2505, n_334, n_4817, n_4115, n_2999, n_2014, n_1239, n_3697, n_1584, n_470, n_3680, n_5381, n_2408, n_5723, n_5918, n_3468, n_5045, n_1972, n_4383, n_4491, n_5696, n_455, n_363, n_4486, n_1816, n_393, n_503, n_5848, n_3024, n_4612, n_5673, n_5443, n_2531, n_5163, n_307, n_4529, n_500, n_3361, n_714, n_3478, n_3936, n_1349, n_291, n_2723, n_5485, n_5823, n_2800, n_3496, n_5473, n_4390, n_3096, n_2651, n_2095, n_3239, n_3161, n_2799, n_5537, n_3902, n_4062, n_3295, n_4396, n_1998, n_1574, n_3101, n_240, n_756, n_1981, n_4233, n_1606, n_3374, n_2640, n_253, n_1552, n_2918, n_583, n_3288, n_4307, n_3992, n_3876, n_249, n_3125, n_4293, n_941, n_3552, n_1031, n_115, n_849, n_4684, n_3116, n_4091, n_1753, n_5027, n_3095, n_2471, n_4412, n_2807, n_1921, n_3618, n_4580, n_1055, n_2217, n_2197, n_4758, n_5630, n_4781, n_4148, n_2461, n_271, n_206, n_4057, n_633, n_1170, n_5379, n_5335, n_308, n_3444, n_1040, n_3059, n_2634, n_1761, n_5424, n_1890, n_3017, n_1805, n_2477, n_5505, n_5868, n_2308, n_2333, n_3001, n_1089, n_3795, n_3852, n_1365, n_4138, n_5289, n_5018, n_3815, n_3896, n_5274, n_3274, n_5401, n_4457, n_4093, n_1616, n_1862, n_5989, n_339, n_434, n_64, n_288, n_4928, n_5769, n_4794, n_722, n_5613, n_5612, n_2223, n_4197, n_4482, n_629, n_1621, n_2547, n_2415, n_5073, n_827, n_4834, n_4762, n_192, n_5581, n_3113, n_992, n_3813, n_3660, n_3766, n_1613, n_1458, n_5303, n_1027, n_3266, n_3574, n_1189, n_223, n_4154, n_4907, n_5077, n_5034, n_726, n_50, n_4504, n_365, n_3844, n_1237, n_2534, n_4975, n_3741, n_5375, n_2451, n_5370, n_2243, n_4815, n_4898, n_5601, n_5784, n_3443, n_509, n_4819, n_1209, n_5248, n_1708, n_805, n_396, n_350, n_78, n_2051, n_4370, n_2359, n_5112, n_480, n_142, n_1402, n_1691, n_3332, n_4134, n_1238, n_2570, n_4092, n_4645, n_3668, n_2491, n_1264, n_4755, n_4359, n_4960, n_4087, n_1700, n_5635, n_4933, n_5091, n_3487, n_4591, n_5528, n_287, n_4302, n_5111, n_3340, n_230, n_5227, n_461, n_873, n_3946, n_2989, n_5778, n_3395, n_4474, n_5665, n_2509, n_2513, n_3757, n_5363, n_4178, n_5165, n_1704, n_2247, n_250, n_1711, n_4884, n_1579, n_3275, n_836, n_522, n_3678, n_3440, n_2094, n_1511, n_2356, n_1422, n_1772, n_4692, n_616, n_3165, n_1119, n_5788, n_1433, n_1902, n_1842, n_1620, n_2739, n_1735, n_3890, n_1541, n_1300, n_641, n_3750, n_1313, n_3607, n_3316, n_516, n_2418, n_2864, n_4311, n_1180, n_2703, n_3371, n_4722, n_4606, n_3261, n_666, n_4187, n_940, n_2058, n_405, n_213, n_2660, n_5317, n_1094, n_5430, n_5942, n_4962, n_4563, n_494, n_5056, n_4820, n_2394, n_5540, n_3532, n_5716, n_3948, n_2124, n_4619, n_381, n_5762, n_4327, n_1961, n_5211, n_5336, n_3765, n_5447, n_4125, n_5036, n_4221, n_3297, n_976, n_3067, n_2155, n_2686, n_5327, n_2364, n_4392, n_2996, n_3803, n_2085, n_917, n_5014, n_5747, n_3639, n_5192, n_4334, n_659, n_3351, n_808, n_5519, n_4047, n_5753, n_3413, n_1193, n_5233, n_3412, n_3791, n_3164, n_4575, n_551, n_699, n_4320, n_3884, n_5808, n_451, n_5436, n_5139, n_757, n_594, n_5231, n_2190, n_6068, n_3438, n_166, n_4141, n_5193, n_2850, n_572, n_1481, n_1441, n_3373, n_5789, n_92, n_2104, n_513, n_3883, n_5961, n_261, n_5866, n_3728, n_2925, n_4499, n_121, n_5822, n_433, n_5195, n_3949, n_5726, n_2792, n_219, n_5364, n_3315, n_263, n_5533, n_3798, n_788, n_1543, n_1599, n_329, n_4257, n_4458, n_2674, n_5103, n_4641, n_4720, n_4893, n_61, n_3857, n_1876, n_4107, n_243, n_1873, n_3630, n_3518, n_1866, n_117, n_2130, n_1330, n_1413, n_3714, n_2228, n_5039, n_2455, n_2876, n_4772, n_5953, n_3099, n_5198, n_4468, n_5718, n_4161, n_1663, n_4172, n_3403, n_2714, n_2245, n_4961, n_4454, n_1107, n_2457, n_3294, n_4119, n_6001, n_3686, n_4502, n_5958, n_318, n_2971, n_1713, n_715, n_4277, n_4526, n_1265, n_3490, n_4849, n_530, n_277, n_4319, n_3369, n_618, n_199, n_5792, n_3581, n_3069, n_6023, n_2028, n_3715, n_1069, n_612, n_3725, n_3933, n_5554, n_1175, n_2311, n_429, n_1012, n_3691, n_5553, n_4485, n_4066, n_903, n_4146, n_5711, n_1802, n_1504, n_4340, n_5790, n_286, n_254, n_3961, n_4855, n_1801, n_2347, n_3917, n_47, n_816, n_1188, n_2206, n_4004, n_2967, n_5404, n_2916, n_5739, n_4292, n_5972, n_2467, n_5549, n_267, n_3145, n_1124, n_1624, n_3983, n_4940, n_5444, n_3538, n_3280, n_5757, n_1515, n_961, n_4356, n_3510, n_2824, n_593, n_637, n_2377, n_701, n_950, n_3009, n_5824, n_3719, n_2525, n_4361, n_5488, n_3827, n_891, n_5154, n_2067, n_3889, n_2687, n_1630, n_2887, n_4245, n_4136, n_3526, n_2194, n_2619, n_5329, n_4367, n_5637, n_1987, n_507, n_968, n_2271, n_1008, n_2583, n_4560, n_2606, n_4899, n_5728, n_5471, n_1033, n_462, n_1052, n_2794, n_5164, n_2391, n_304, n_2431, n_5843, n_125, n_2078, n_2932, n_1767, n_3431, n_3450, n_449, n_4663, n_2893, n_1208, n_5484, n_2954, n_2728, n_1072, n_815, n_3421, n_3183, n_2493, n_4802, n_2705, n_5523, n_1067, n_3405, n_5423, n_255, n_284, n_1952, n_5074, n_4044, n_3436, n_1026, n_1880, n_3442, n_3366, n_2631, n_38, n_289, n_3937, n_1293, n_3159, n_4701, n_108, n_794, n_727, n_894, n_685, n_353, n_3240, n_3576, n_1863, n_3385, n_4851, n_3293, n_872, n_3922, n_86, n_5204, n_5333, n_847, n_644, n_682, n_851, n_4991, n_5594, n_72, n_2554, n_5422, n_1513, n_1913, n_4934, n_837, n_5087, n_5526, n_5292, n_2517, n_2713, n_5000, n_2765, n_5403, n_2590, n_5551, n_3150, n_2060, n_4479, n_2608, n_4011, n_5131, n_1959, n_3133, n_5257, n_765, n_1492, n_1340, n_4688, n_4753, n_4058, n_631, n_2262, n_3611, n_3082, n_4848, n_5059, n_156, n_5887, n_843, n_2604, n_2407, n_1277, n_2816, n_3799, n_2574, n_4475, n_5242, n_5219, n_2675, n_5631, n_3537, n_4443, n_3887, n_6008, n_1022, n_614, n_5854, n_2667, n_5460, n_4587, n_1615, n_4114, n_1474, n_1571, n_2948, n_1577, n_2119, n_947, n_1117, n_1992, n_5686, n_5899, n_3223, n_3140, n_3185, n_4749, n_2605, n_5155, n_118, n_926, n_3654, n_1849, n_2848, n_919, n_1698, n_4100, n_4264, n_5981, n_3788, n_89, n_4891, n_5937, n_777, n_1299, n_5339, n_3837, n_2718, n_1436, n_1384, n_3325, n_2238, n_6040, n_4085, n_4464, n_4624, n_4818, n_4659, n_3600, n_18, n_5217, n_5465, n_5015, n_4339, n_1178, n_98, n_2338, n_3324, n_796, n_1195, n_184, n_1811, n_1857, n_3987, n_1519, n_6039, n_2144, n_1284, n_1604, n_4487, n_4889, n_4866, n_1142, n_623, n_1048, n_5721, n_3638, n_4816, n_2110, n_5719, n_1502, n_5773, n_1659, n_5482, n_3393, n_6012, n_3451, n_1418, n_1250, n_292, n_4937, n_5277, n_3615, n_3072, n_3087, n_2053, n_2259, n_2121, n_4222, n_4874, n_4401, n_889, n_2710, n_6064, n_3142, n_4015, n_1966, n_5793, n_477, n_1110, n_4709, n_2213, n_4976, n_2389, n_2132, n_2892, n_4120, n_1564, n_5578, n_4658, n_231, n_2860, n_2330, n_40, n_5296, n_1457, n_505, n_3718, n_5893, n_1787, n_537, n_1993, n_2281, n_2617, n_2776, n_1466, n_10, n_1919, n_5742, n_5207, n_3705, n_3211, n_3909, n_5676, n_546, n_386, n_1220, n_6051, n_1893, n_2301, n_4665, n_3582, n_4223, n_2387, n_5674, n_3270, n_5539, n_2846, n_5282, n_970, n_2488, n_1980, n_5464, n_2237, n_1060, n_1951, n_444, n_4362, n_1252, n_3311, n_3913, n_1223, n_511, n_5121, n_6026, n_6070, n_1286, n_2115, n_4430, n_3302, n_4348, n_5013, n_1597, n_4489, n_4839, n_2596, n_3163, n_775, n_4404, n_1153, n_5589, n_439, n_1531, n_2828, n_453, n_2384, n_4261, n_4204, n_759, n_2724, n_426, n_2585, n_5628, n_4825, n_2352, n_1625, n_3986, n_5006, n_4513, n_4006, n_2226, n_2801, n_1901, n_3869, n_2556, n_4747, n_1647, n_5251, n_3753, n_2306, n_1614, n_1892, n_3742, n_3683, n_4801, n_401, n_3260, n_2550, n_3175, n_3736, n_5475, n_5807, n_4448, n_1096, n_2227, n_5216, n_3284, n_4869, n_427, n_2159, n_4386, n_688, n_1077, n_2315, n_4132, n_2995, n_5273, n_1437, n_4844, n_4438, n_4836, n_5439, n_4955, n_4149, n_5936, n_4355, n_501, n_2276, n_3234, n_856, n_2803, n_379, n_1668, n_2777, n_3202, n_2830, n_3220, n_1129, n_602, n_2181, n_6069, n_171, n_2911, n_169, n_4655, n_1429, n_5706, n_2826, n_3429, n_2379, n_326, n_587, n_3554, n_1593, n_1202, n_1635, n_5431, n_4067, n_4357, n_28, n_3462, n_2851, n_4374, n_5132, n_106, n_358, n_160, n_2420, n_5627, n_5774, n_3722, n_186, n_4400, n_4846, n_5798, n_2984, n_575, n_5187, n_5875, n_4024, n_1508, n_5621, n_5608, n_732, n_2983, n_2240, n_392, n_2538, n_724, n_3250, n_1042, n_4582, n_1728, n_557, n_1871, n_4860, n_845, n_140, n_5844, n_3414, n_1549, n_4870, n_768, n_3651, n_2102, n_2563, n_4989, n_3449, n_1683, n_1916, n_2598, n_597, n_280, n_1187, n_4304, n_4558, n_1403, n_4488, n_3767, n_2544, n_3550, n_4211, n_1206, n_4016, n_5867, n_621, n_750, n_5508, n_4656, n_3839, n_2823, n_5597, n_4915, n_4328, n_1057, n_2785, n_235, n_5515, n_1997, n_5662, n_2636, n_3131, n_710, n_1818, n_3730, n_1298, n_5862, n_4397, n_3399, n_2088, n_1611, n_5050, n_2740, n_746, n_4808, n_5697, n_3416, n_3498, n_5767, n_2401, n_101, n_1589, n_4712, n_2309, n_2900, n_2957, n_1740, n_2737, n_3994, n_5462, n_1497, n_133, n_5980, n_3672, n_5318, n_3533, n_1622, n_4725, n_6022, n_4406, n_1694, n_1535, n_3382, n_3132, n_5498, n_2571, n_3138, n_20, n_5053, n_2171, n_2988, n_4908, n_3136, n_1350, n_4109, n_4192, n_4824, n_2037, n_2808, n_4567, n_5150, n_782, n_809, n_3819, n_4778, n_5477, n_1797, n_5175, n_986, n_2050, n_4595, n_2164, n_4174, n_402, n_1870, n_1171, n_460, n_5987, n_5179, n_1827, n_4904, n_2187, n_1152, n_450, n_3544, n_4150, n_2904, n_5988, n_5585, n_6058, n_711, n_3105, n_2872, n_3692, n_4616, n_4982, n_370, n_1695, n_2046, n_2272, n_2760, n_1979, n_4643, n_2738, n_972, n_5348, n_1332, n_5480, n_4323, n_624, n_2346, n_4831, n_936, n_3045, n_3821, n_885, n_83, n_2342, n_2167, n_2970, n_3676, n_4896, n_2882, n_3666, n_3675, n_4017, n_4260, n_4916, n_2541, n_2940, n_5904, n_4739, n_599, n_6062, n_105, n_1974, n_4122, n_934, n_4209, n_2768, n_3858, n_1341, n_5284, n_4298, n_2314, n_3502, n_5461, n_3003, n_4128, n_543, n_5147, n_4271, n_4644, n_1355, n_2258, n_5503, n_325, n_5845, n_5945, n_804, n_2390, n_959, n_2562, n_4716, n_4312, n_1343, n_1522, n_76, n_2734, n_1782, n_5600, n_5755, n_707, n_1900, n_5048, n_6053, n_3246, n_1548, n_3381, n_1155, n_2195, n_3208, n_4944, n_5245, n_4343, n_4715, n_4935, n_4694, n_4672, n_5054, n_2962, n_5448, n_2939, n_5749, n_1672, n_1925, n_4407, n_737, n_4045, n_3517, n_2945, n_4598, n_3061, n_3893, n_3932, n_21, n_3469, n_2960, n_5993, n_138, n_3258, n_4524, n_3143, n_6020, n_333, n_4084, n_3149, n_3365, n_3379, n_24, n_459, n_4850, n_4424, n_3008, n_1751, n_2840, n_285, n_3939, n_4776, n_1375, n_3972, n_4153, n_85, n_3506, n_1650, n_1962, n_3855, n_1928, n_3091, n_4317, n_4723, n_4269, n_5418, n_4088, n_3398, n_5685, n_2761, n_2793, n_3776, n_3711, n_4235, n_5459, n_1019, n_4143, n_4170, n_729, n_876, n_774, n_3642, n_2845, n_4650, n_438, n_4719, n_5173, n_1860, n_5016, n_1904, n_2874, n_1200, n_2588, n_479, n_1353, n_1777, n_4967, n_3308, n_1113, n_1600, n_2253, n_2366, n_4912, n_4799, n_2261, n_4423, n_5086, n_5283, n_2210, n_4735, n_3602, n_187, n_3300, n_2978, n_2516, n_1050, n_1411, n_5170, n_2827, n_1177, n_3515, n_1150, n_566, n_1023, n_2951, n_1118, n_194, n_2949, n_1807, n_5028, n_5839, n_1814, n_1631, n_1879, n_256, n_440, n_3806, n_5514, n_2931, n_209, n_367, n_2569, n_3866, n_5351, n_5909, n_671, n_4543, n_740, n_703, n_4157, n_4229, n_5293, n_3865, n_4073, n_1324, n_3629, n_1435, n_5400, n_3920, n_969, n_4892, n_3255, n_1401, n_1516, n_3846, n_180, n_3512, n_5201, n_2029, n_5890, n_4439, n_1394, n_1326, n_4783, n_1379, n_214, n_935, n_4910, n_1130, n_3083, n_676, n_832, n_3049, n_5389, n_5142, n_3830, n_3679, n_5891, n_3541, n_74, n_3117, n_5935, n_4930, n_372, n_111, n_314, n_378, n_5623, n_338, n_1283, n_2385, n_4112, n_506, n_360, n_2149, n_2396, n_4557, n_4917, n_895, n_2450, n_3739, n_4432, n_2284, n_4352, n_4416, n_4593, n_344, n_2769, n_4465, n_3622, n_5114, n_4980, n_1392, n_5693, n_4495, n_5117, n_1924, n_5663, n_525, n_2463, n_3363, n_1677, n_5990, n_611, n_3721, n_3062, n_2679, n_5024, n_4559, n_838, n_3969, n_129, n_3336, n_4160, n_4231, n_2952, n_5647, n_1017, n_4256, n_2779, n_4938, n_5396, n_5203, n_109, n_445, n_930, n_2620, n_5162, n_1945, n_5426, n_1656, n_5803, n_2112, n_1464, n_2430, n_653, n_1414, n_5285, n_2721, n_944, n_4335, n_2034, n_576, n_270, n_2683, n_563, n_5365, n_2744, n_1011, n_4521, n_1566, n_626, n_990, n_3204, n_1104, n_5715, n_4920, n_498, n_870, n_5395, n_1253, n_366, n_5709, n_1693, n_3256, n_348, n_3802, n_376, n_2118, n_2111, n_390, n_2915, n_1148, n_2188, n_1989, n_2802, n_3643, n_2425, n_4265, n_2950, n_5634, n_5672, n_719, n_3060, n_3098, n_4105, n_1851, n_1090, n_4861, n_5799, n_4064, n_4926, n_1518, n_1362, n_3123, n_3380, n_5617, n_1829, n_5266, n_5580, n_1450, n_4828, n_1638, n_3038, n_570, n_1789, n_620, n_519, n_2523, n_5450, n_2413, n_3769, n_1482, n_5310, n_3863, n_3669, n_3130, n_4316, n_5722, n_4640, n_5122, n_5390, n_1710, n_2161, n_1301, n_2805, n_5593, n_33, n_4769, n_5764, n_2282, n_4628, n_2047, n_5385, n_1609, n_3344, n_5237, n_2334, n_5133, n_409, n_1763, n_5322, n_3989, n_2490, n_4460, n_4108, n_635, n_3786, n_3841, n_4254, n_1996, n_2867, n_1442, n_2726, n_4303, n_5853, n_5982, n_1158, n_2248, n_5011, n_5917, n_2662, n_4909, n_3147, n_753, n_3925, n_3180, n_2795, n_3472, n_5376, n_5106, n_269, n_359, n_1479, n_4768, n_1675, n_3717, n_5561, n_5410, n_571, n_2215, n_404, n_158, n_1884, n_665, n_2055, n_5156, n_2553, n_149, n_632, n_2038, n_4447, n_4826, n_3445, n_373, n_87, n_1833, n_3903, n_5998, n_1494, n_2325, n_1850, n_5304, n_3854, n_3235, n_5378, n_6028, n_1417, n_3673, n_4281, n_5916, n_681, n_4648, n_3094, n_412, n_965, n_1428, n_1576, n_1856, n_2077, n_5691, n_1059, n_4951, n_422, n_4957, n_3079, n_165, n_4360, n_540, n_4039, n_457, n_3070, n_3800, n_4566, n_3263, n_4853, n_1748, n_3504, n_531, n_4272, n_2930, n_5615, n_1025, n_3111, n_336, n_12, n_1885, n_5269, n_3054, n_1538, n_1240, n_5468, n_1, n_4730, n_5399, n_1234, n_5262, n_3254, n_3684, n_4670, n_4882, n_4620, n_3152, n_4738, n_3579, n_5421, n_3335, n_4177, n_3783, n_700, n_1307, n_3178, n_4127, n_5206, n_1003, n_5713, n_5256, n_168, n_2353, n_4099, n_4517, n_77, n_4168, n_5188, n_1738, n_4490, n_1575, n_1923, n_2260, n_3952, n_5550, n_3911, n_1688, n_4285, n_3465, n_1743, n_2997, n_1991, n_2386, n_5161, n_5373, n_1724, n_3708, n_4078, n_3046, n_2956, n_5573, n_1553, n_5939, n_5509, n_5382, n_5659, n_3619, n_1415, n_5881, n_1370, n_1786, n_4198, n_2382, n_3754, n_2291, n_415, n_1371, n_383, n_2886, n_2974, n_4213, n_200, n_2184, n_2982, n_1803, n_4065, n_5863, n_229, n_2645, n_3904, n_1393, n_1517, n_1867, n_2630, n_1444, n_1603, n_2470, n_4446, n_1263, n_4417, n_5466, n_4733, n_4764, n_1261, n_3879, n_2286, n_4743, n_2018, n_3080, n_1903, n_1143, n_5955, n_658, n_1874, n_2865, n_2825, n_2013, n_2044, n_3023, n_3232, n_693, n_1056, n_758, n_5851, n_2256, n_943, n_4060, n_5110, n_4879, n_5796, n_42, n_772, n_2806, n_770, n_3028, n_3662, n_2981, n_3076, n_886, n_343, n_3624, n_1345, n_1820, n_4556, n_539, n_45, n_4117, n_4687, n_2836, n_638, n_1404, n_5492, n_5995, n_2378, n_887, n_5905, n_2655, n_4600, n_126, n_1467, n_4250, n_5829, n_3906, n_224, n_4954, n_5191, n_1231, n_2599, n_3963, n_3368, n_9, n_2370, n_2612, n_2591, n_4881, n_1815, n_2214, n_4253, n_407, n_913, n_5734, n_2593, n_4255, n_867, n_4071, n_3568, n_1230, n_3850, n_5770, n_1333, n_2496, n_5705, n_3313, n_4605, n_3189, n_5525, n_163, n_1644, n_2725, n_2277, n_4691, n_1558, n_1732, n_2300, n_3943, n_4305, n_824, n_4297, n_6052, n_2907, n_577, n_5374, n_5575, n_1843, n_619, n_5675, n_4227, n_521, n_2778, n_395, n_1909, n_5020, n_606, n_5297, n_1123, n_1309, n_2961, n_916, n_3934, n_4033, n_4415, n_483, n_1970, n_630, n_2059, n_2669, n_4094, n_4765, n_2546, n_3193, n_2522, n_476, n_4364, n_1957, n_4354, n_4732, n_3912, n_3118, n_5959, n_3720, n_1907, n_2529, n_264, n_860, n_1530, n_4745, n_938, n_1302, n_5642, n_4581, n_549, n_4377, n_2143, n_905, n_4792, n_1680, n_3842, n_322, n_993, n_689, n_2031, n_4878, n_1605, n_3514, n_4979, n_1988, n_558, n_2654, n_3036, n_5302, n_966, n_4511, n_2908, n_3357, n_692, n_5639, n_5781, n_1233, n_3895, n_487, n_241, n_4520, n_5299, n_3455, n_4118, n_4503, n_2176, n_2459, n_1111, n_3599, n_5543, n_1251, n_5361, n_2711, n_4199, n_5885, n_1912, n_5356, n_4441, n_1982, n_3872, n_3772, n_5458, n_1312, n_5668, n_5038, n_268, n_1760, n_5330, n_4585, n_2664, n_5, n_1664, n_1722, n_5463, n_3022, n_247, n_5489, n_1165, n_5892, n_4773, n_5654, n_2008, n_6009, n_2192, n_3281, n_2345, n_328, n_1386, n_4427, n_5923, n_5113, n_5479, n_3549, n_5714, n_2804, n_2453, n_2676, n_5510, n_3940, n_4822, n_1214, n_690, n_850, n_5692, n_4800, n_1157, n_3453, n_5555, n_3410, n_1752, n_1813, n_3768, n_4958, n_2810, n_4043, n_2319, n_5441, n_825, n_6066, n_3785, n_2963, n_5366, n_2602, n_55, n_3873, n_2980, n_696, n_4886, n_1082, n_1317, n_3227, n_2733, n_3289, n_4055, n_2178, n_5968, n_2644, n_2036, n_3326, n_4200, n_3460, n_2411, n_1796, n_2082, n_3519, n_678, n_5078, n_3707, n_283, n_3578, n_909, n_4737, n_590, n_4925, n_4116, n_5415, n_362, n_22, n_5419, n_1990, n_3805, n_2943, n_5205, n_1634, n_3252, n_627, n_3253, n_1465, n_342, n_2622, n_2658, n_2665, n_2133, n_1712, n_4603, n_1523, n_1627, n_5080, n_5976, n_3128, n_1527, n_495, n_5732, n_5372, n_2691, n_840, n_2913, n_4471, n_2230, n_1969, n_2690, n_5208, n_1565, n_1493, n_5690, n_2573, n_2646, n_2535, n_1364, n_3078, n_2436, n_615, n_3838, n_5371, n_4651, n_3941, n_3793, n_4854, n_5071, n_3789, n_605, n_1514, n_5801, n_6047, n_3037, n_1646, n_3729, n_4994, n_2537, n_4483, n_5347, n_5168, n_4661, n_1308, n_4988, n_3171, n_3608, n_4540, n_2097, n_79, n_3459, n_2853, n_1808, n_3053, n_3358, n_6021, n_3499, n_4284, n_1005, n_1947, n_3426, n_4971, n_5656, n_1469, n_5125, n_5857, n_2650, n_5652, n_987, n_5499, n_720, n_153, n_3229, n_3348, n_1707, n_656, n_5228, n_797, n_2933, n_2717, n_1723, n_1878, n_189, n_738, n_2012, n_3497, n_5066, n_2842, n_3580, n_2335, n_529, n_2307, n_3704, n_684, n_5507, n_1809, n_5569, n_4280, n_1181, n_37, n_5190, n_3173, n_3677, n_3996, n_1049, n_4097, n_1666, n_803, n_4218, n_5392, n_1717, n_1817, n_2449, n_3880, n_3685, n_2868, n_2231, n_3609, n_1228, n_5455, n_417, n_5442, n_5948, n_4459, n_4545, n_272, n_2896, n_3019, n_2639, n_3471, n_5511, n_2898, n_69, n_5295, n_2368, n_53, n_458, n_4175, n_5490, n_16, n_3200, n_4771, n_3259, n_2524, n_3167, n_2460, n_5836, n_3867, n_3593, n_4455, n_1073, n_252, n_4514, n_5834, n_3191, n_5584, n_4140, n_2481, n_3561, n_4806, n_2682, n_3032, n_5160, n_2877, n_5098, n_1021, n_811, n_683, n_1207, n_5707, n_5140, n_4992, n_5197, n_5497, n_880, n_3505, n_3540, n_3577, n_2432, n_150, n_1478, n_4796, n_3598, n_4442, n_2581, n_1363, n_3641, n_3777, n_4203, n_767, n_1837, n_2218, n_4533, n_831, n_5481, n_3590, n_2435, n_5344, n_954, n_4419, n_5308, n_1410, n_5184, n_5794, n_1382, n_5408, n_1736, n_4053, n_1483, n_3848, n_1372, n_3327, n_1719, n_319, n_2701, n_2511, n_4167, n_1427, n_2745, n_1080, n_5271, n_123, n_562, n_5964, n_6004, n_2323, n_2784, n_5494, n_162, n_5234, n_4431, n_2421, n_1136, n_4387, n_2618, n_3265, n_2464, n_128, n_1125, n_3755, n_4042, n_5128, n_2224, n_2329, n_1092, n_441, n_5467, n_4299, n_4890, n_146, n_1784, n_3571, n_193, n_1775, n_2410, n_1093, n_1783, n_2929, n_4176, n_5827, n_5199, n_296, n_651, n_3407, n_5992, n_217, n_5313, n_1185, n_3856, n_4236, n_3425, n_215, n_3894, n_3127, n_1831, n_2621, n_3623, n_5312, n_5079, n_54, n_1453, n_2502, n_3646, n_5513, n_5614, n_497, n_4830, n_4706, n_1315, n_5225, n_4570, n_2754, n_1224, n_2783, n_3188, n_1459, n_2462, n_3243, n_1135, n_2889, n_4034, n_4056, n_4622, n_3960, n_1470, n_4887, n_2732, n_4693, n_4206, n_2249, n_1091, n_2000, n_3862, n_4267, n_5835, n_2270, n_1425, n_5049, n_983, n_5846, n_906, n_1390, n_2289, n_1733, n_2955, n_5592, n_2158, n_4609, n_1855, n_3051, n_3367, n_385, n_1687, n_1439, n_2328, n_2859, n_2202, n_1331, n_613, n_736, n_5278, n_3314, n_3525, n_2100, n_5157, n_2993, n_4754, n_3016, n_4647, n_1134, n_3688, n_4003, n_5708, n_554, n_1995, n_3751, n_5223, n_4894, n_5474, n_4113, n_1889, n_4760, n_5649, n_435, n_1905, n_3466, n_762, n_5704, n_4983, n_1778, n_5956, n_5287, n_1079, n_2139, n_419, n_5083, n_4509, n_6007, n_2875, n_1103, n_3907, n_3338, n_144, n_4217, n_4906, n_2219, n_1203, n_3636, n_2327, n_999, n_5516, n_1254, n_2841, n_4897, n_3539, n_3291, n_4399, n_2304, n_2487, n_5698, n_3276, n_2597, n_3194, n_5084, n_5771, n_3572, n_349, n_3886, n_4710, n_4420, n_443, n_892, n_3637, n_4574, n_1468, n_2855, n_1859, n_2156, n_1718, n_5174, n_4234, n_5538, n_4101, n_3548, n_5017, n_1768, n_3974, n_198, n_1847, n_3634, n_1397, n_3236, n_901, n_2755, n_3141, n_923, n_5096, n_1841, n_4660, n_5241, n_1623, n_1015, n_3112, n_4797, n_3108, n_4270, n_5428, n_4151, n_4945, n_3417, n_5677, n_4124, n_5570, n_73, n_785, n_5153, n_609, n_4611, n_5927, n_5435, n_2337, n_1356, n_3213, n_4333, n_127, n_3820, n_5200, n_2607, n_2890, n_1168, n_5115, n_1943, n_5566, n_3249, n_1320, n_2722, n_1452, n_2854, n_2499, n_4152, n_5487, n_302, n_5486, n_137, n_1596, n_5092, n_5244, n_1734, n_3172, n_4832, n_2902, n_5889, n_3217, n_1983, n_5391, n_1938, n_2472, n_3394, n_1715, n_3536, n_1443, n_1272, n_2894, n_3957, n_3710, n_4195, n_5849, n_4554, n_3040, n_3279, n_5240, n_2402, n_2225, n_1081, n_5951, n_1692, n_1084, n_5912, n_1864, n_2006, n_3402, n_3475, n_3501, n_374, n_1705, n_3905, n_4680, n_3013, n_921, n_579, n_2789, n_5152, n_5265, n_2257, n_4927, n_5574, n_4258, n_1828, n_2699, n_2200, n_650, n_1940, n_4548, n_4862, n_1405, n_2376, n_5469, n_456, n_3878, n_2670, n_313, n_2700, n_5910, n_5895, n_1041, n_5804, n_565, n_3134, n_5965, n_1569, n_3115, n_1062, n_896, n_4553, n_3278, n_2084, n_4875, n_5682, n_5387, n_654, n_5557, n_411, n_2458, n_1222, n_3050, n_2673, n_2456, n_2527, n_2635, n_1637, n_3307, n_1407, n_1795, n_2871, n_420, n_4321, n_4183, n_164, n_5681, n_1271, n_4901, n_1545, n_4821, n_4145, n_3121, n_1640, n_4040, n_2406, n_806, n_584, n_2141, n_5316, n_244, n_548, n_282, n_5703, n_833, n_523, n_345, n_3930, n_4943, n_799, n_3044, n_4757, n_2196, n_2629, n_2809, n_787, n_2172, n_4682, n_5564, n_5620, n_4530, n_1528, n_1146, n_2021, n_4942, n_159, n_1086, n_5406, n_2125, n_2561, n_652, n_4604, n_1906, n_3305, n_2992, n_5724, n_1241, n_3157, n_4841, n_1758, n_3221, n_3267, n_2422, n_1914, n_1318, n_5806, n_4338, n_3457, n_306, n_3762, n_5738, n_3005, n_3151, n_3411, n_4840, n_1029, n_4519, n_3779, n_2388, n_5355, n_3984, n_5320, n_5353, n_1706, n_5186, n_5710, n_1498, n_2417, n_1210, n_5093, n_1556, n_4052, n_5979, n_3558, n_1984, n_2236, n_5438, n_6044, n_4326, n_1269, n_2083, n_2834, n_5517, n_3207, n_5605, n_2441, n_3401, n_3242, n_3613, n_655, n_4726, n_1045, n_5907, n_786, n_1559, n_6045, n_1872, n_19, n_29, n_75, n_5040, n_6063, n_1325, n_3761, n_4315, n_2888, n_2923, n_1727, n_4301, n_151, n_3744, n_4788, n_2041, n_1360, n_5977, n_3814, n_3781, n_1908, n_2484, n_2126, n_6003, n_3843, n_1098, n_5746, n_2045, n_817, n_5451, n_3687, n_2216, n_5402, n_3543, n_3621, n_6031, n_2903, n_3216, n_332, n_3808, n_398, n_4365, n_6060, n_1882, n_3726, n_1007, n_1929, n_2369, n_1592, n_2719, n_591, n_3758, n_5417, n_2587, n_3199, n_680, n_3339, n_4923, n_2400, n_5864, n_1953, n_4741, n_3343, n_2752, n_4885, n_751, n_5432, n_1399, n_4550, n_4652, n_2358, n_5453, n_3658, n_4900, n_2163, n_2186, n_2815, n_3034, n_4408, n_4577, n_4748, n_643, n_5842, n_400, n_337, n_5814, n_2814, n_5253, n_5209, n_789, n_3231, n_4212, n_2979, n_5699, n_181, n_5531, n_5765, n_2953, n_327, n_4295, n_5943, n_2946, n_2500, n_3430, n_2269, n_1729, n_5777, n_4225, n_300, n_747, n_2565, n_5495, n_1389, n_535, n_3583, n_3860, n_3851, n_5655, n_5064, n_5610, n_3015, n_2175, n_601, n_2182, n_4009, n_1848, n_5002, n_5759, n_1506, n_119, n_3473, n_1652, n_6035, n_957, n_1994, n_2566, n_387, n_744, n_971, n_2702, n_3241, n_2906, n_4342, n_4568, n_1205, n_6061, n_5559, n_1258, n_2438, n_2914, n_5786, n_3100, n_2180, n_2858, n_5377, n_3573, n_1016, n_4106, n_5737, n_1501, n_3604, n_4373, n_197, n_4711, n_3068, n_2685, n_1083, n_5768, n_3553, n_2275, n_2465, n_2568, n_2022, n_3811, n_910, n_3494, n_1721, n_1737, n_3486, n_4086, n_752, n_908, n_1028, n_2106, n_2265, n_5350, n_5470, n_2032, n_4812, n_4409, n_5872, n_5858, n_4629, n_4638, n_708, n_1973, n_3181, n_5700, n_1500, n_6037, n_3699, n_854, n_4913, n_2312, n_5874, n_904, n_709, n_1266, n_2242, n_3328, n_185, n_3868, n_1276, n_4266, n_2466, n_2530, n_5873, n_1085, n_2042, n_771, n_475, n_924, n_298, n_1582, n_492, n_5588, n_2318, n_3286, n_4012, n_1149, n_3170, n_265, n_3645, n_5075, n_3682, n_3304, n_2592, n_4968, n_3771, n_2666, n_1585, n_1799, n_2564, n_5085, n_5736, n_4259, n_2433, n_829, n_2035, n_3422, n_4572, n_859, n_3086, n_2033, n_406, n_4104, n_4845, n_1770, n_878, n_5120, n_130, n_3285, n_4208, n_981, n_5928, n_4089, n_5478, n_6016, n_1144, n_2071, n_3219, n_3702, n_2233, n_4779, n_481, n_3233, n_4599, n_997, n_4437, n_5222, n_3310, n_1306, n_3264, n_2010, n_1198, n_4061, n_2174, n_436, n_3881, n_4508, n_4727, n_4594, n_2426, n_2478, n_1133, n_95, n_4429, n_4642, n_4051, n_1051, n_4865, n_1039, n_2043, n_1480, n_6056, n_5832, n_3206, n_1305, n_2363, n_2578, n_4562, n_553, n_3383, n_4903, n_3709, n_3738, n_4186, n_5812, n_2540, n_973, n_5743, n_3610, n_4998, n_3330, n_2065, n_2879, n_967, n_4522, n_2001, n_4341, n_679, n_1629, n_5368, n_4263, n_225, n_1260, n_1819, n_309, n_3555, n_915, n_5971, n_812, n_1131, n_3155, n_1006, n_3110, n_1632, n_5933, n_257, n_1888, n_1311, n_4780, n_670, n_2697, n_3908, n_4973, n_3467, n_1887, n_1587, n_3916, n_3527, n_4803, n_2512, n_3950, n_6030, n_1242, n_2086, n_2927, n_4750, n_3039, n_1226, n_3740, n_5996, n_2166, n_2899, n_3186, n_640, n_1322, n_1958, n_315, n_5903, n_5986, n_1197, n_3065, n_2632, n_4984, n_2579, n_2105, n_135, n_1423, n_3387, n_364, n_5782, n_3420, n_5041, n_1915, n_4275, n_4283, n_4959, n_900, n_4426, n_2912, n_60, n_2659, n_4425, n_3409, n_4449, n_2116, n_2320, n_1013, n_1259, n_2183, n_3002, n_51, n_649, n_1612, n_4809, n_1199, n_3392, n_6050, n_625, n_226, n_68, n_212, n_3773, n_2003, n_1038, n_1581, n_3301, n_1357, n_4241, n_1853, n_798, n_2324, n_5563, n_245, n_1348, n_2977, n_1739, n_5840, n_1380, n_2847, n_2557, n_1009, n_62, n_2405, n_4050, n_1160, n_883, n_2647, n_1032, n_2336, n_1247, n_5717, n_6017, n_2521, n_1099, n_471, n_424, n_4578, n_2211, n_4777, n_5720, n_369, n_2672, n_4702, n_2299, n_4179, n_4895, n_5871, n_141, n_1285, n_1985, n_5898, n_1172, n_4026, n_71, n_4531, n_3282, n_1590, n_3626, n_1532, n_2313, n_5072, n_3106, n_1140, n_1670, n_2344, n_2365, n_4666, n_3031, n_4029, n_375, n_2447, n_4617, n_2340, n_4010, n_5896, n_1649, n_4555, n_5882, n_5940, n_5650, n_4969, n_6057, n_5105, n_1572, n_4308, n_5021, n_3463, n_428, n_5263, n_2510, n_1954, n_822, n_2791, n_4325, n_3251, n_4602, n_5044, n_5134, n_2212, n_3063, n_1163, n_2729, n_2582, n_1798, n_1550, n_491, n_3998, n_1591, n_3632, n_3122, n_5567, n_1344, n_2730, n_2495, n_371, n_5249, n_2090, n_2603, n_538, n_3829, n_4164, n_2173, n_5625, n_1471, n_4919, n_3737, n_5969, n_3655, n_493, n_3825, n_2880, n_3225, n_2108, n_5158, n_1211, n_5022, n_5670, n_1280, n_6041, n_3296, n_5276, n_58, n_1445, n_2551, n_1526, n_5047, n_196, n_2985, n_1978, n_574, n_3792, n_4202, n_1446, n_14, n_3938, n_4791, n_3507, n_5879, n_4403, n_5238, n_5855, n_3269, n_3531, n_473, n_1054, n_559, n_1956, n_4139, n_4549, n_1986, n_2397, n_3931, n_4349, n_5141, n_2113, n_1918, n_3603, n_5429, n_813, n_3822, n_4163, n_818, n_5535, n_645, n_3812, n_3910, n_2633, n_2207, n_4948, n_5268, n_2696, n_3482, n_4080, n_6002, n_2198, n_3319, n_541, n_2073, n_2273, n_3748, n_3272, n_4941, n_5506, n_5298, n_2, n_3396, n_4393, n_1162, n_4372, n_821, n_1068, n_982, n_5640, n_408, n_932, n_2831, n_4318, n_4158, n_3317, n_3978, n_5560, n_2123, n_1697, n_979, n_4074, n_3716, n_4795, n_5544, n_4918, n_3824, n_5067, n_5744, n_4013, n_5384, n_4544, n_3248, n_354, n_5841, n_134, n_2941, n_1278, n_547, n_5108, n_4032, n_1064, n_1396, n_634, n_2355, n_4147, n_136, n_4477, n_3168, n_2751, n_4337, n_4130, n_5941, n_2009, n_1793, n_3601, n_5611, n_3092, n_1289, n_3055, n_3966, n_2866, n_4742, n_1014, n_3734, n_1703, n_2580, n_882, n_3649, n_2821, n_1875, n_1865, n_5701, n_3746, n_6067, n_3384, n_1950, n_1563, n_3419, n_1297, n_1662, n_4478, n_1359, n_2818, n_5367, n_3794, n_674, n_3921, n_922, n_1335, n_1927, n_4838, n_5970, n_5202, n_702, n_4965, n_347, n_3346, n_1896, n_2965, n_3058, n_3861, n_675, n_1540, n_1977, n_3891, n_2193, n_4523, n_1655, n_242, n_6011, n_1886, n_4371, n_2994, n_5502, n_3428, n_3153, n_4552, n_3689, n_877, n_5850, n_4673, n_2519, n_728, n_3415, n_1063, n_4607, n_4041, n_2947, n_3918, n_5876, n_5521, n_1965, n_4837, n_2476, n_598, n_437, n_4169, n_697, n_3271, n_295, n_5088, n_4248, n_388, n_484, n_2976, n_2152, n_2652, n_1825, n_1757, n_170, n_1792, n_5856, n_1412, n_2497, n_3809, n_3139, n_4070, n_3545, n_3885, n_1369, n_881, n_3993, n_4685, n_63, n_4031, n_5837, n_148, n_4675, n_2663, n_5825, n_4018, n_5491, n_2987, n_694, n_2938, n_3780, n_5496, n_5802, n_297, n_3337, n_4002, n_3209, n_5178, n_1044, n_2165, n_5547, n_1391, n_131, n_2750, n_2775, n_1295, n_3477, n_2349, n_5596, n_6074, n_2684, n_5983, n_3146, n_1495, n_1438, n_3953, n_4588, n_1100, n_585, n_4653, n_4435, n_5604, n_1756, n_1128, n_5411, n_673, n_4019, n_1071, n_1968, n_4728, n_4999, n_4385, n_4922, n_865, n_3616, n_5815, n_4191, n_5695, n_6027, n_2870, n_59, n_2151, n_1839, n_2341, n_1765, n_3727, n_5235, n_2707, n_826, n_4350, n_3747, n_1714, n_104, n_718, n_5331, n_4330, n_542, n_5311, n_305, n_2089, n_3522, n_2747, n_3924, n_791, n_4621, n_4216, n_5797, n_510, n_4240, n_3491, n_5572, n_1488, n_704, n_2148, n_4162, n_5565, n_2339, n_2861, n_1999, n_2731, n_622, n_5520, n_147, n_3353, n_3018, n_3975, n_5800, n_5984, n_1838, n_2638, n_4785, n_4683, n_1766, n_1776, n_2002, n_2138, n_4021, n_2414, n_3014, n_1771, n_2316, n_4103, n_5060, n_3148, n_4022, n_4986, n_5888, n_5669, n_5772, n_145, n_2208, n_4775, n_5884, n_4864, n_5758, n_4674, n_4481, n_1304, n_294, n_3775, n_4669, n_2134, n_1176, n_425, n_5603, n_1431, n_3312, n_3835, n_4286, n_5763, n_2958, n_3731, n_1822, n_2936, n_3224, n_2489, n_6029, n_1087, n_657, n_5751, n_2771, n_3020, n_5264, n_4525, n_5924, n_1505, n_290, n_5712, n_3557, n_2610, n_3129, n_3620, n_478, n_107, n_3832, n_2520, n_4484, n_3693, n_446, n_4497, n_1568, n_2372, n_1490, n_526, n_2251, n_3674, n_2959, n_2501, n_3203, n_5694, n_4871, n_293, n_1070, n_2403, n_2837, n_4700, n_4883, n_1665, n_4306, n_154, n_4224, n_2127, n_3341, n_6005, n_4453, n_3559, n_5449, n_4005, n_3546, n_1358, n_3661, n_4564, n_5146, n_3056, n_745, n_2424, n_3201, n_3447, n_3971, n_5926, n_716, n_1475, n_1774, n_2354, n_3103, n_4573, n_5398, n_5860, n_2589, n_4535, n_755, n_527, n_2442, n_3627, n_3480, n_1368, n_1137, n_3612, n_4695, n_2545, n_3509, n_5919, n_4368, n_2966, n_2294, n_1942, n_1314, n_600, n_3196, n_864, n_5319, n_2504, n_2623, n_399, n_1440, n_5270, n_2063, n_1534, n_5005, n_6014, n_1339, n_2475, n_5181, n_403, n_723, n_3144, n_3244, n_596, n_1141, n_1268, n_3287, n_3322, n_1755, n_5043, n_2025, n_2357, n_5583, n_4654, n_3640, n_642, n_995, n_1159, n_3481, n_2250, n_3033, n_303, n_5775, n_2374, n_416, n_1681, n_6034, n_520, n_418, n_4597, n_113, n_3364, n_3226, n_2780, n_4020, n_5220, n_1618, n_4867, n_5061, n_1653, n_4063, n_4237, n_2601, n_5029, n_5127, n_6071, n_2920, n_773, n_920, n_99, n_1374, n_2648, n_3212, n_13, n_1169, n_1617, n_3370, n_3386, n_335, n_4721, n_463, n_3093, n_848, n_120, n_274, n_4247, n_3169, n_3205, n_1881, n_1267, n_1806, n_2023, n_2204, n_2720, n_496, n_4614, n_177, n_3360, n_2087, n_1636, n_3956, n_4001, n_1323, n_2627, n_4422, n_960, n_778, n_3004, n_3870, n_5177, n_5483, n_3625, n_1764, n_4632, n_1610, n_3084, n_5785, n_2343, n_793, n_5967, n_4546, n_4583, n_4963, n_3749, n_2942, n_4966, n_5780, n_4714, n_5037, n_2515, n_316, n_1551, n_4847, n_4054, n_2555, n_3586, n_3653, n_5966, n_2201, n_725, n_3349, n_4668, n_5213, n_4635, n_0, n_368, n_994, n_5735, n_2278, n_1020, n_1273, n_4214, n_3448, n_617, n_2924, n_1036, n_3595, n_1138, n_5752, n_1661, n_5360, n_421, n_3991, n_3516, n_3926, n_1095, n_1270, n_4405, n_610, n_4413, n_1852, n_4036, n_4759, n_2153, n_3670, n_2381, n_2052, n_179, n_4667, n_5081, n_517, n_4182, n_667, n_3230, n_1279, n_1115, n_1499, n_504, n_1409, n_5877, n_6018, n_5189, n_1503, n_2819, n_3041, n_4637, n_2423, n_603, n_1657, n_1126, n_2412, n_5869, n_2439, n_2404, n_1182, n_3635, n_5118, n_4155, n_4238, n_3011, n_2061, n_2757, n_4977, n_167, n_5632, n_5582, n_5425, n_5886, n_1216, n_2716, n_6032, n_2452, n_3650, n_5446, n_3010, n_3043, n_5224, n_4590, n_2543, n_5090, n_3137, n_2486, n_3560, n_3177, n_4929, n_5678, n_122, n_2220, n_2577, n_34, n_1262, n_3238, n_218, n_3529, n_70, n_4835, n_2232, n_4038, n_2790, n_4565, n_5414, n_4159, n_3784, n_5437, n_220, n_4586, n_1608, n_2373, n_1472, n_3628, n_5454, n_800, n_4734, n_1491, n_1840, n_4434, n_5307, n_2244, n_4290, n_2586, n_1684, n_2446, n_1346, n_1352, n_5407, n_2017, n_3029, n_3597, n_5913, n_1046, n_2560, n_2704, n_1145, n_1121, n_1102, n_1963, n_258, n_3790, n_2766, n_260, n_356, n_3318, n_4833, n_5062, n_5230, n_5944, n_152, n_4888, n_776, n_321, n_1823, n_2479, n_3350, n_6000, n_2782, n_3977, n_227, n_3588, n_4279, n_5008, n_1456, n_5004, n_5294, n_23, n_5974, n_2229, n_4133, n_4527, n_2288, n_6046, n_2099, n_5323, n_3388, n_4790, n_1946, n_4181, n_3184, n_5810, n_4561, n_4461, n_464, n_3245, n_3075, n_4007, n_4949, n_2642, n_4239, n_2383, n_5991, n_4184, n_1676, n_1830, n_2351, n_1319, n_5069, n_2986, n_5702, n_2536, n_3915, n_139, n_1633, n_3489, n_2835, n_5243, n_1416, n_5914, n_2820, n_2293, n_5250, n_3074, n_3102, n_5590, n_2026, n_1282, n_5260, n_550, n_3321, n_2567, n_5809, n_2322, n_275, n_2727, n_3377, n_560, n_4782, n_1321, n_2533, n_569, n_3530, n_2869, n_4378, n_5349, n_1235, n_2759, n_2361, n_1292, n_2266, n_4876, n_346, n_3, n_5813, n_790, n_5833, n_2611, n_2901, n_4358, n_5616, n_5805, n_2653, n_49, n_299, n_1248, n_902, n_2189, n_2246, n_4469, n_5169, n_431, n_5816, n_3156, n_672, n_1941, n_3483, n_5416, n_706, n_1794, n_1236, n_4493, n_4924, n_743, n_766, n_430, n_1746, n_3524, n_489, n_2885, n_636, n_110, n_3097, n_660, n_2062, n_4539, n_2975, n_4421, n_6072, n_2839, n_2856, n_4793, n_4498, n_2070, n_1607, n_1454, n_4953, n_2348, n_2944, n_3831, n_869, n_1154, n_646, n_528, n_391, n_1329, n_5167, n_5661, n_5830, n_5932, n_3589, n_262, n_897, n_846, n_2066, n_841, n_1476, n_3391, n_508, n_1800, n_1463, n_3458, n_4505, n_3190, n_1562, n_5558, n_1826, n_5687, n_57, n_5383, n_5126, n_1759, n_5051, n_52, n_5587, n_5236, n_853, n_875, n_5012, n_1678, n_661, n_3787, n_1256, n_3585, n_3565, n_4450, n_5954, n_7, n_5025, n_933, n_4173, n_3135, n_5651, n_4630, n_1217, n_5645, n_3990, n_310, n_1628, n_5766, n_2109, n_988, n_2796, n_2507, n_84, n_5878, n_5671, n_4534, n_1536, n_1204, n_1132, n_233, n_1327, n_955, n_246, n_2787, n_2969, n_2395, n_1554, n_4494, n_5412, n_769, n_2380, n_4786, n_1120, n_555, n_4579, n_669, n_2290, n_4811, n_2048, n_176, n_114, n_2005, n_4857, n_3432, n_2736, n_2883, n_1408, n_4282, n_1196, n_3493, n_863, n_3774, n_5733, n_2910, n_748, n_3268, n_1785, n_1147, n_1754, n_3057, n_3701, n_5148, n_2584, n_1812, n_866, n_2287, n_452, n_5791, n_5727, n_761, n_5946, n_5997, n_2492, n_3778, n_5328, n_5657, n_174, n_1173, n_4974, n_5975, n_4911, n_4436, n_5119, n_4569, n_1174, n_3334, n_5938, n_5602, n_647, n_5097, n_844, n_17, n_4985, n_2117, n_2234, n_3823, n_4384, n_2741, n_3114, n_888, n_2203, n_2255, n_3584, n_5246, n_236, n_4858, n_4678, n_2649, n_3556, n_3836, n_5579, n_414, n_1922, n_5750, n_4823, n_5831, n_4309, n_4363, n_1215, n_93, n_839, n_5107, n_3456, n_5095, n_779, n_1537, n_2205, n_4243, n_4025, n_3404, n_1122, n_5666, n_4059, n_1509, n_4121, n_3290, n_1109, n_4313, n_3309, n_3671, n_4142, n_2015, n_3982, n_2609, n_1161, n_5546, n_3796, n_232, n_3840, n_46, n_3461, n_3408, n_4246, n_3513, n_3690, n_1184, n_2483, n_4532, n_228, n_1525, n_3995, n_4076, n_2594, n_5994, n_4244, n_2147, n_592, n_2503, n_4049, n_1156, n_2600, n_984, n_5626, n_3508, n_132, n_868, n_4353, n_735, n_4787, n_5633, n_469, n_1218, n_5664, n_5921, n_3596, n_4537, n_4346, n_4351, n_357, n_2429, n_985, n_2440, n_6054, n_3521, n_802, n_561, n_980, n_2681, n_1651, n_2360, n_3764, n_4784, n_4075, n_116, n_5340, n_3947, n_1244, n_1685, n_3066, n_2844, n_2303, n_1619, n_2285, n_5280, n_4451, n_4332, n_810, n_1194, n_4538, n_4506, n_2742, n_3695, n_3976, n_3563, n_2367, n_201, n_3198, n_3495, n_1034, n_5925, n_2909, n_754, n_5369, n_975, n_43, n_5730, n_5576, n_3359, n_5272, n_467, n_3187, n_3218, n_582, n_861, n_857, n_2107, n_2040, n_2968, n_4201, n_4336, n_2221, n_588, n_5646, n_5624, n_4852, n_1010, n_4210, n_4981, n_1166, n_5440, n_2891, n_2709, n_534, n_1578, n_1861, n_3955, n_1557, n_2280, n_3945, n_730, n_5817, n_5214, n_203, n_1898, n_2443, n_4936, n_4205, n_2162, n_1868, n_207, n_2079, n_4763, n_3587, n_4278, n_5586, n_3433, n_4463, n_205, n_2185, n_6038, n_5861, n_1836, n_3833, n_2774, n_3162, n_1274, n_1486, n_3333, n_4129, n_5258, n_81, n_5032, n_1899, n_784, n_4804, n_5619, n_3965, n_5859, n_5380, n_4500, n_5065, n_862, n_5776, n_2098, n_3085, n_4433, n_5606, n_5644, n_2813, n_1935, n_5826, n_2027, n_2091, n_5920, n_2991, n_5030, n_4194, n_1449, n_4703, n_361, n_2419, n_5683, n_2677, n_3182, n_5756, n_3283, n_5527, n_1742, n_4030, n_20644);

input n_5643;
input n_2542;
input n_1671;
input n_2817;
input n_801;
input n_4452;
input n_2576;
input n_5172;
input n_4649;
input n_1674;
input n_5315;
input n_741;
input n_1351;
input n_5254;
input n_1212;
input n_208;
input n_5362;
input n_4251;
input n_2157;
input n_5019;
input n_2332;
input n_3849;
input n_578;
input n_5138;
input n_4388;
input n_4395;
input n_1061;
input n_3089;
input n_783;
input n_5653;
input n_4978;
input n_5409;
input n_5301;
input n_188;
input n_1854;
input n_3088;
input n_3257;
input n_1342;
input n_4829;
input n_5393;
input n_1387;
input n_3222;
input n_677;
input n_4699;
input n_1151;
input n_4686;
input n_2317;
input n_5524;
input n_442;
input n_5345;
input n_1975;
input n_1930;
input n_3706;
input n_5818;
input n_2179;
input n_5963;
input n_5055;
input n_1547;
input n_3376;
input n_4868;
input n_893;
input n_3801;
input n_5267;
input n_4249;
input n_5950;
input n_1192;
input n_3564;
input n_1844;
input n_1555;
input n_5548;
input n_5057;
input n_3030;
input n_830;
input n_65;
input n_5838;
input n_5725;
input n_447;
input n_2838;
input n_5229;
input n_5325;
input n_3427;
input n_852;
input n_5101;
input n_2628;
input n_3071;
input n_2926;
input n_1078;
input n_544;
input n_5900;
input n_4273;
input n_5545;
input n_35;
input n_2321;
input n_2019;
input n_5102;
input n_3345;
input n_2074;
input n_2919;
input n_4501;
input n_2129;
input n_4724;
input n_945;
input n_5598;
input n_4997;
input n_2399;
input n_4843;
input n_1232;
input n_4696;
input n_4347;
input n_5259;
input n_5819;
input n_2480;
input n_3877;
input n_3929;
input n_3048;
input n_1455;
input n_5279;
input n_2786;
input n_5894;
input n_5930;
input n_5239;
input n_567;
input n_1781;
input n_1971;
input n_5354;
input n_5332;
input n_2004;
input n_1106;
input n_4814;
input n_953;
input n_3979;
input n_5908;
input n_3077;
input n_2873;
input n_3452;
input n_3107;
input n_155;
input n_4956;
input n_454;
input n_1421;
input n_3664;
input n_1936;
input n_5337;
input n_5129;
input n_5420;
input n_1660;
input n_5070;
input n_3047;
input n_4414;
input n_112;
input n_713;
input n_1400;
input n_2625;
input n_4646;
input n_2843;
input n_3760;
input n_6015;
input n_48;
input n_1560;
input n_4262;
input n_734;
input n_1088;
input n_1894;
input n_3347;
input n_5136;
input n_907;
input n_6;
input n_5638;
input n_4110;
input n_1658;
input n_4950;
input n_4729;
input n_4268;
input n_1967;
input n_3999;
input n_3928;
input n_2613;
input n_3535;
input n_4751;
input n_44;
input n_2708;
input n_1648;
input n_5151;
input n_1911;
input n_2011;
input n_5684;
input n_5729;
input n_281;
input n_564;
input n_5680;
input n_279;
input n_686;
input n_4102;
input n_1641;
input n_3871;
input n_2735;
input n_4662;
input n_4671;
input n_3959;
input n_2268;
input n_1367;
input n_5504;
input n_1336;
input n_5522;
input n_5828;
input n_4314;
input n_2080;
input n_323;
input n_5099;
input n_1381;
input n_331;
input n_1699;
input n_2093;
input n_4296;
input n_102;
input n_2770;
input n_608;
input n_2101;
input n_4507;
input n_32;
input n_5902;
input n_512;
input n_3484;
input n_4677;
input n_792;
input n_5063;
input n_1328;
input n_2917;
input n_2616;
input n_5275;
input n_5306;
input n_3923;
input n_3900;
input n_3488;
input n_939;
input n_2811;
input n_3732;
input n_2832;
input n_4226;
input n_5493;
input n_1762;
input n_1910;
input n_1075;
input n_3980;
input n_2998;
input n_5346;
input n_4366;
input n_3446;
input n_5252;
input n_5309;
input n_237;
input n_1895;
input n_4294;
input n_4698;
input n_4445;
input n_4810;
input n_3859;
input n_2692;
input n_175;
input n_3914;
input n_4456;
input n_3397;
input n_3575;
input n_2469;
input n_3927;
input n_5452;
input n_3888;
input n_764;
input n_5476;
input n_2764;
input n_2895;
input n_733;
input n_2922;
input n_3882;
input n_4856;
input n_3492;
input n_4369;
input n_30;
input n_2068;
input n_4331;
input n_4972;
input n_1290;
input n_4993;
input n_5536;
input n_2072;
input n_1354;
input n_586;
input n_423;
input n_4375;
input n_1701;
input n_6055;
input n_2678;
input n_3935;
input n_5130;
input n_4291;
input n_88;
input n_5532;
input n_5897;
input n_1726;
input n_4613;
input n_2434;
input n_2878;
input n_3012;
input n_3875;
input n_5609;
input n_1167;
input n_2428;
input n_4717;
input n_4877;
input n_3247;
input n_871;
input n_5922;
input n_210;
input n_2641;
input n_5658;
input n_4731;
input n_3052;
input n_178;
input n_355;
input n_5046;
input n_2749;
input n_3298;
input n_2254;
input n_5058;
input n_1926;
input n_3273;
input n_4467;
input n_1747;
input n_195;
input n_5667;
input n_780;
input n_2624;
input n_5865;
input n_2350;
input n_5042;
input n_5305;
input n_4681;
input n_4072;
input n_4752;
input n_4220;
input n_835;
input n_928;
input n_5281;
input n_2092;
input n_1654;
input n_1750;
input n_1462;
input n_2514;
input n_604;
input n_5314;
input n_1588;
input n_3942;
input n_3997;
input n_26;
input n_2468;
input n_4381;
input n_5144;
input n_515;
input n_2096;
input n_3968;
input n_4466;
input n_4418;
input n_3434;
input n_4510;
input n_5795;
input n_4473;
input n_6043;
input n_5552;
input n_5226;
input n_514;
input n_687;
input n_890;
input n_5457;
input n_2812;
input n_190;
input n_4518;
input n_1709;
input n_2393;
input n_2657;
input n_5291;
input n_2921;
input n_2136;
input n_2409;
input n_2252;
input n_3237;
input n_949;
input n_3500;
input n_3834;
input n_4589;
input n_2075;
input n_2972;
input n_3542;
input n_91;
input n_2763;
input n_2762;
input n_3192;
input n_760;
input n_1546;
input n_4394;
input n_2279;
input n_161;
input n_6010;
input n_1296;
input n_3352;
input n_3073;
input n_5343;
input n_2150;
input n_1294;
input n_3696;
input n_1420;
input n_4082;
input n_595;
input n_1779;
input n_524;
input n_4921;
input n_1858;
input n_4329;
input n_5135;
input n_3021;
input n_2558;
input n_1164;
input n_4697;
input n_4288;
input n_4289;
input n_3763;
input n_2712;
input n_5529;
input n_3733;
input n_6042;
input n_1487;
input n_3614;
input n_874;
input n_382;
input n_5183;
input n_2145;
input n_898;
input n_4964;
input n_5957;
input n_4228;
input n_3423;
input n_925;
input n_1932;
input n_1101;
input n_15;
input n_4636;
input n_4322;
input n_3644;
input n_1249;
input n_4946;
input n_2706;
input n_4767;
input n_4287;
input n_2693;
input n_4137;
input n_1127;
input n_1512;
input n_1451;
input n_320;
input n_639;
input n_963;
input n_2767;
input n_4576;
input n_5929;
input n_4615;
input n_5787;
input n_1139;
input n_3179;
input n_1018;
input n_3400;
input n_1521;
input n_1366;
input n_4000;
input n_5445;
input n_2897;
input n_4389;
input n_3970;
input n_5342;
input n_5501;
input n_4345;
input n_996;
input n_532;
input n_173;
input n_1376;
input n_413;
input n_4664;
input n_2170;
input n_4156;
input n_948;
input n_6033;
input n_977;
input n_536;
input n_3158;
input n_1788;
input n_4873;
input n_2643;
input n_5748;
input n_3782;
input n_1835;
input n_3470;
input n_5076;
input n_581;
input n_5870;
input n_4713;
input n_4098;
input n_5026;
input n_4476;
input n_432;
input n_3700;
input n_4995;
input n_3166;
input n_3104;
input n_3435;
input n_842;
input n_5636;
input n_2239;
input n_4310;
input n_1432;
input n_5212;
input n_989;
input n_2689;
input n_1473;
input n_5286;
input n_2191;
input n_1246;
input n_4528;
input n_5811;
input n_899;
input n_1035;
input n_4914;
input n_4939;
input n_499;
input n_1426;
input n_3418;
input n_705;
input n_11;
input n_1004;
input n_1529;
input n_5530;
input n_2473;
input n_5397;
input n_4634;
input n_2069;
input n_2362;
input n_4096;
input n_2539;
input n_2698;
input n_4123;
input n_5595;
input n_3119;
input n_5427;
input n_3735;
input n_2297;
input n_4379;
input n_486;
input n_5388;
input n_4718;
input n_1448;
input n_5901;
input n_5962;
input n_3631;
input n_5599;
input n_648;
input n_2445;
input n_5324;
input n_2057;
input n_2103;
input n_3770;
input n_2772;
input n_4440;
input n_4402;
input n_927;
input n_5052;
input n_4541;
input n_5009;
input n_4872;
input n_929;
input n_4551;
input n_2857;
input n_5326;
input n_1183;
input n_4627;
input n_4079;
input n_2494;
input n_5300;
input n_3342;
input n_998;
input n_5035;
input n_717;
input n_1383;
input n_3390;
input n_3656;
input n_1424;
input n_1000;
input n_3025;
input n_2137;
input n_1626;
input n_1507;
input n_2482;
input n_3810;
input n_552;
input n_4798;
input n_2532;
input n_1388;
input n_3006;
input n_216;
input n_912;
input n_5010;
input n_2296;
input n_3633;
input n_5352;
input n_5089;
input n_2849;
input n_1201;
input n_1398;
input n_884;
input n_5394;
input n_4592;
input n_1395;
input n_2199;
input n_2661;
input n_731;
input n_5359;
input n_1955;
input n_931;
input n_474;
input n_312;
input n_1791;
input n_66;
input n_958;
input n_5137;
input n_100;
input n_3331;
input n_5104;
input n_1897;
input n_2064;
input n_5741;
input n_2773;
input n_5405;
input n_5288;
input n_589;
input n_3606;
input n_1310;
input n_819;
input n_1334;
input n_3591;
input n_2788;
input n_964;
input n_4756;
input n_2797;
input n_4746;
input n_124;
input n_3892;
input n_4970;
input n_4069;
input n_211;
input n_2748;
input n_5194;
input n_1834;
input n_2331;
input n_2292;
input n_3441;
input n_3534;
input n_5952;
input n_3964;
input n_2416;
input n_311;
input n_5947;
input n_1877;
input n_3944;
input n_1939;
input n_2030;
input n_1769;
input n_5985;
input n_556;
input n_2209;
input n_3605;
input n_1602;
input n_4633;
input n_3306;
input n_276;
input n_3026;
input n_221;
input n_4584;
input n_3090;
input n_5232;
input n_3724;
input n_4276;
input n_5116;
input n_2990;
input n_3847;
input n_1773;
input n_5001;
input n_2552;
input n_1053;
input n_5176;
input n_4428;
input n_1533;
input n_3323;
input n_4;
input n_266;
input n_2274;
input n_5761;
input n_518;
input n_4618;
input n_4679;
input n_1745;
input n_914;
input n_3479;
input n_4496;
input n_317;
input n_4805;
input n_1679;
input n_90;
input n_3454;
input n_2160;
input n_5760;
input n_2146;
input n_2131;
input n_488;
input n_5472;
input n_3547;
input n_5679;
input n_2575;
input n_5100;
input n_5973;
input n_4410;
input n_1933;
input n_1179;
input n_324;
input n_3816;
input n_4807;
input n_4411;
input n_3214;
input n_1243;
input n_301;
input n_2928;
input n_5166;
input n_1917;
input n_1580;
input n_2822;
input n_36;
input n_4180;
input n_1281;
input n_3109;
input n_3354;
input n_2572;
input n_1520;
input n_3126;
input n_3663;
input n_2863;
input n_1419;
input n_3299;
input n_5688;
input n_351;
input n_5740;
input n_259;
input n_1731;
input n_5820;
input n_5648;
input n_2135;
input n_5745;
input n_4707;
input n_1645;
input n_1832;
input n_4676;
input n_5180;
input n_858;
input n_2049;
input n_5182;
input n_956;
input n_5534;
input n_663;
input n_4880;
input n_3566;
input n_2781;
input n_4126;
input n_410;
input n_2829;
input n_1696;
input n_3845;
input n_1594;
input n_664;
input n_1869;
input n_3804;
input n_4207;
input n_5196;
input n_2016;
input n_5171;
input n_4470;
input n_580;
input n_4813;
input n_5542;
input n_1030;
input n_3901;
input n_1937;
input n_465;
input n_1790;
input n_5261;
input n_4014;
input n_4704;
input n_341;
input n_1744;
input n_828;
input n_2142;
input n_4252;
input n_607;
input n_4028;
input n_2448;
input n_5949;
input n_4048;
input n_4596;
input n_4444;
input n_5255;
input n_3756;
input n_3406;
input n_820;
input n_951;
input n_952;
input n_3919;
input n_2263;
input n_5185;
input n_974;
input n_4952;
input n_2656;
input n_5023;
input n_2375;
input n_5906;
input n_1934;
input n_628;
input n_5660;
input n_1434;
input n_1573;
input n_3981;
input n_3973;
input n_2756;
input n_5334;
input n_6024;
input n_807;
input n_4761;
input n_1275;
input n_2884;
input n_485;
input n_67;
input n_1510;
input n_5783;
input n_3120;
input n_5821;
input n_3797;
input n_238;
input n_2024;
input n_1595;
input n_4770;
input n_202;
input n_1749;
input n_3474;
input n_2549;
input n_4690;
input n_1669;
input n_1024;
input n_3864;
input n_5556;
input n_4932;
input n_5456;
input n_248;
input n_2302;
input n_1667;
input n_1037;
input n_5143;
input n_3592;
input n_468;
input n_5500;
input n_4230;
input n_2637;
input n_1639;
input n_183;
input n_3967;
input n_3195;
input n_466;
input n_2526;
input n_4274;
input n_5215;
input n_3277;
input n_2548;
input n_5386;
input n_991;
input n_4189;
input n_3817;
input n_340;
input n_1108;
input n_3659;
input n_2559;
input n_2177;
input n_39;
input n_2595;
input n_5003;
input n_4827;
input n_1601;
input n_1960;
input n_2694;
input n_3648;
input n_1686;
input n_6059;
input n_3042;
input n_6065;
input n_5094;
input n_4610;
input n_4472;
input n_5433;
input n_6075;
input n_3228;
input n_3657;
input n_96;
input n_3081;
input n_1430;
input n_1316;
input n_1287;
input n_5618;
input n_1586;
input n_2264;
input n_3464;
input n_380;
input n_3723;
input n_1190;
input n_397;
input n_4380;
input n_5978;
input n_4990;
input n_4996;
input n_5247;
input n_4398;
input n_2498;
input n_4515;
input n_1891;
input n_5031;
input n_1213;
input n_6006;
input n_2235;
input n_4193;
input n_3570;
input n_5082;
input n_1673;
input n_5338;
input n_3828;
input n_172;
input n_2392;
input n_3424;
input n_4131;
input n_239;
input n_97;
input n_2298;
input n_2326;
input n_1539;
input n_490;
input n_3594;
input n_5689;
input n_1043;
input n_4090;
input n_4165;
input n_2305;
input n_2120;
input n_80;
input n_4626;
input n_6048;
input n_4144;
input n_2964;
input n_352;
input n_2169;
input n_3485;
input n_4077;
input n_5931;
input n_2371;
input n_1361;
input n_662;
input n_3262;
input n_4008;
input n_3356;
input n_5221;
input n_5641;
input n_1642;
input n_3210;
input n_937;
input n_4689;
input n_1682;
input n_4547;
input n_5731;
input n_3329;
input n_330;
input n_3826;
input n_4905;
input n_1406;
input n_4601;
input n_962;
input n_3647;
input n_3681;
input n_1883;
input n_4300;
input n_1288;
input n_1186;
input n_4623;
input n_5007;
input n_3320;
input n_2518;
input n_5883;
input n_5754;
input n_3988;
input n_1720;
input n_3476;
input n_4842;
input n_204;
input n_482;
input n_5629;
input n_3439;
input n_4135;
input n_2688;
input n_394;
input n_1845;
input n_1489;
input n_942;
input n_2798;
input n_2852;
input n_1524;
input n_1964;
input n_1920;
input n_2753;
input n_1496;
input n_3292;
input n_2007;
input n_2039;
input n_5434;
input n_5934;
input n_1225;
input n_1544;
input n_1485;
input n_1846;
input n_3437;
input n_4111;
input n_533;
input n_3712;
input n_4608;
input n_879;
input n_2310;
input n_2506;
input n_4859;
input n_94;
input n_2626;
input n_5880;
input n_1567;
input n_4037;
input n_3562;
input n_5852;
input n_2973;
input n_5218;
input n_41;
input n_3665;
input n_273;
input n_3007;
input n_3528;
input n_5960;
input n_4571;
input n_3698;
input n_5358;
input n_3355;
input n_2454;
input n_2114;
input n_3174;
input n_5321;
input n_1066;
input n_1948;
input n_157;
input n_4215;
input n_2154;
input n_6073;
input n_1484;
input n_5290;
input n_4185;
input n_3752;
input n_2283;
input n_5145;
input n_4219;
input n_1229;
input n_1373;
input n_3958;
input n_3985;
input n_2427;
input n_4196;
input n_1447;
input n_4774;
input n_2056;
input n_5210;
input n_4242;
input n_5109;
input n_3389;
input n_4232;
input n_4190;
input n_4902;
input n_3000;
input n_5149;
input n_5571;
input n_2680;
input n_1047;
input n_3375;
input n_3899;
input n_1385;
input n_3713;
input n_1931;
input n_502;
input n_2668;
input n_1257;
input n_3197;
input n_4987;
input n_2128;
input n_5512;
input n_4736;
input n_2398;
input n_1725;
input n_3743;
input n_834;
input n_5033;
input n_2695;
input n_4035;
input n_3818;
input n_3124;
input n_1741;
input n_1002;
input n_1949;
input n_3759;
input n_545;
input n_2671;
input n_4516;
input n_2715;
input n_1804;
input n_251;
input n_2508;
input n_3511;
input n_2054;
input n_6025;
input n_1337;
input n_1477;
input n_2614;
input n_4492;
input n_2833;
input n_2758;
input n_5607;
input n_3694;
input n_2937;
input n_4789;
input n_5999;
input n_4376;
input n_1001;
input n_2241;
input n_4708;
input n_4657;
input n_1690;
input n_5341;
input n_1191;
input n_1076;
input n_4512;
input n_1378;
input n_855;
input n_1377;
input n_695;
input n_4081;
input n_1542;
input n_4542;
input n_4462;
input n_1716;
input n_278;
input n_4931;
input n_4536;
input n_5562;
input n_3303;
input n_978;
input n_4324;
input n_384;
input n_1976;
input n_4382;
input n_2905;
input n_1291;
input n_749;
input n_1824;
input n_3954;
input n_5911;
input n_2122;
input n_5622;
input n_2140;
input n_3503;
input n_3160;
input n_1065;
input n_5577;
input n_1255;
input n_568;
input n_5124;
input n_143;
input n_3951;
input n_823;
input n_1074;
input n_698;
input n_3569;
input n_739;
input n_3874;
input n_2528;
input n_5123;
input n_4639;
input n_5413;
input n_1338;
input n_1097;
input n_3027;
input n_781;
input n_4083;
input n_1810;
input n_182;
input n_5915;
input n_573;
input n_1583;
input n_4480;
input n_1730;
input n_2295;
input n_2746;
input n_389;
input n_814;
input n_5779;
input n_1643;
input n_2020;
input n_4171;
input n_3652;
input n_222;
input n_4023;
input n_1105;
input n_721;
input n_1461;
input n_742;
input n_691;
input n_3617;
input n_2076;
input n_6019;
input n_3567;
input n_377;
input n_1598;
input n_4344;
input n_2935;
input n_4705;
input n_4046;
input n_3807;
input n_918;
input n_1114;
input n_56;
input n_763;
input n_4027;
input n_3154;
input n_1227;
input n_2485;
input n_3898;
input n_3520;
input n_191;
input n_6036;
input n_4391;
input n_946;
input n_1303;
input n_4095;
input n_2881;
input n_1116;
input n_1570;
input n_1702;
input n_1219;
input n_3551;
input n_4947;
input n_3064;
input n_1780;
input n_3897;
input n_1689;
input n_8;
input n_5591;
input n_3372;
input n_1944;
input n_1347;
input n_795;
input n_1221;
input n_6013;
input n_1245;
input n_3215;
input n_448;
input n_3853;
input n_4740;
input n_4631;
input n_1561;
input n_1112;
input n_5518;
input n_2081;
input n_2168;
input n_5068;
input n_234;
input n_5847;
input n_6049;
input n_1460;
input n_911;
input n_82;
input n_27;
input n_5159;
input n_2862;
input n_472;
input n_2615;
input n_4068;
input n_4625;
input n_2474;
input n_3703;
input n_2437;
input n_2444;
input n_25;
input n_3962;
input n_2743;
input n_4766;
input n_4863;
input n_2267;
input n_3035;
input n_668;
input n_4166;
input n_1821;
input n_1058;
input n_3378;
input n_3745;
input n_3362;
input n_4744;
input n_103;
input n_4188;
input n_5357;
input n_2934;
input n_3667;
input n_3523;
input n_2222;
input n_712;
input n_3176;
input n_5541;
input n_5568;
input n_31;
input n_2505;
input n_334;
input n_4817;
input n_4115;
input n_2999;
input n_2014;
input n_1239;
input n_3697;
input n_1584;
input n_470;
input n_3680;
input n_5381;
input n_2408;
input n_5723;
input n_5918;
input n_3468;
input n_5045;
input n_1972;
input n_4383;
input n_4491;
input n_5696;
input n_455;
input n_363;
input n_4486;
input n_1816;
input n_393;
input n_503;
input n_5848;
input n_3024;
input n_4612;
input n_5673;
input n_5443;
input n_2531;
input n_5163;
input n_307;
input n_4529;
input n_500;
input n_3361;
input n_714;
input n_3478;
input n_3936;
input n_1349;
input n_291;
input n_2723;
input n_5485;
input n_5823;
input n_2800;
input n_3496;
input n_5473;
input n_4390;
input n_3096;
input n_2651;
input n_2095;
input n_3239;
input n_3161;
input n_2799;
input n_5537;
input n_3902;
input n_4062;
input n_3295;
input n_4396;
input n_1998;
input n_1574;
input n_3101;
input n_240;
input n_756;
input n_1981;
input n_4233;
input n_1606;
input n_3374;
input n_2640;
input n_253;
input n_1552;
input n_2918;
input n_583;
input n_3288;
input n_4307;
input n_3992;
input n_3876;
input n_249;
input n_3125;
input n_4293;
input n_941;
input n_3552;
input n_1031;
input n_115;
input n_849;
input n_4684;
input n_3116;
input n_4091;
input n_1753;
input n_5027;
input n_3095;
input n_2471;
input n_4412;
input n_2807;
input n_1921;
input n_3618;
input n_4580;
input n_1055;
input n_2217;
input n_2197;
input n_4758;
input n_5630;
input n_4781;
input n_4148;
input n_2461;
input n_271;
input n_206;
input n_4057;
input n_633;
input n_1170;
input n_5379;
input n_5335;
input n_308;
input n_3444;
input n_1040;
input n_3059;
input n_2634;
input n_1761;
input n_5424;
input n_1890;
input n_3017;
input n_1805;
input n_2477;
input n_5505;
input n_5868;
input n_2308;
input n_2333;
input n_3001;
input n_1089;
input n_3795;
input n_3852;
input n_1365;
input n_4138;
input n_5289;
input n_5018;
input n_3815;
input n_3896;
input n_5274;
input n_3274;
input n_5401;
input n_4457;
input n_4093;
input n_1616;
input n_1862;
input n_5989;
input n_339;
input n_434;
input n_64;
input n_288;
input n_4928;
input n_5769;
input n_4794;
input n_722;
input n_5613;
input n_5612;
input n_2223;
input n_4197;
input n_4482;
input n_629;
input n_1621;
input n_2547;
input n_2415;
input n_5073;
input n_827;
input n_4834;
input n_4762;
input n_192;
input n_5581;
input n_3113;
input n_992;
input n_3813;
input n_3660;
input n_3766;
input n_1613;
input n_1458;
input n_5303;
input n_1027;
input n_3266;
input n_3574;
input n_1189;
input n_223;
input n_4154;
input n_4907;
input n_5077;
input n_5034;
input n_726;
input n_50;
input n_4504;
input n_365;
input n_3844;
input n_1237;
input n_2534;
input n_4975;
input n_3741;
input n_5375;
input n_2451;
input n_5370;
input n_2243;
input n_4815;
input n_4898;
input n_5601;
input n_5784;
input n_3443;
input n_509;
input n_4819;
input n_1209;
input n_5248;
input n_1708;
input n_805;
input n_396;
input n_350;
input n_78;
input n_2051;
input n_4370;
input n_2359;
input n_5112;
input n_480;
input n_142;
input n_1402;
input n_1691;
input n_3332;
input n_4134;
input n_1238;
input n_2570;
input n_4092;
input n_4645;
input n_3668;
input n_2491;
input n_1264;
input n_4755;
input n_4359;
input n_4960;
input n_4087;
input n_1700;
input n_5635;
input n_4933;
input n_5091;
input n_3487;
input n_4591;
input n_5528;
input n_287;
input n_4302;
input n_5111;
input n_3340;
input n_230;
input n_5227;
input n_461;
input n_873;
input n_3946;
input n_2989;
input n_5778;
input n_3395;
input n_4474;
input n_5665;
input n_2509;
input n_2513;
input n_3757;
input n_5363;
input n_4178;
input n_5165;
input n_1704;
input n_2247;
input n_250;
input n_1711;
input n_4884;
input n_1579;
input n_3275;
input n_836;
input n_522;
input n_3678;
input n_3440;
input n_2094;
input n_1511;
input n_2356;
input n_1422;
input n_1772;
input n_4692;
input n_616;
input n_3165;
input n_1119;
input n_5788;
input n_1433;
input n_1902;
input n_1842;
input n_1620;
input n_2739;
input n_1735;
input n_3890;
input n_1541;
input n_1300;
input n_641;
input n_3750;
input n_1313;
input n_3607;
input n_3316;
input n_516;
input n_2418;
input n_2864;
input n_4311;
input n_1180;
input n_2703;
input n_3371;
input n_4722;
input n_4606;
input n_3261;
input n_666;
input n_4187;
input n_940;
input n_2058;
input n_405;
input n_213;
input n_2660;
input n_5317;
input n_1094;
input n_5430;
input n_5942;
input n_4962;
input n_4563;
input n_494;
input n_5056;
input n_4820;
input n_2394;
input n_5540;
input n_3532;
input n_5716;
input n_3948;
input n_2124;
input n_4619;
input n_381;
input n_5762;
input n_4327;
input n_1961;
input n_5211;
input n_5336;
input n_3765;
input n_5447;
input n_4125;
input n_5036;
input n_4221;
input n_3297;
input n_976;
input n_3067;
input n_2155;
input n_2686;
input n_5327;
input n_2364;
input n_4392;
input n_2996;
input n_3803;
input n_2085;
input n_917;
input n_5014;
input n_5747;
input n_3639;
input n_5192;
input n_4334;
input n_659;
input n_3351;
input n_808;
input n_5519;
input n_4047;
input n_5753;
input n_3413;
input n_1193;
input n_5233;
input n_3412;
input n_3791;
input n_3164;
input n_4575;
input n_551;
input n_699;
input n_4320;
input n_3884;
input n_5808;
input n_451;
input n_5436;
input n_5139;
input n_757;
input n_594;
input n_5231;
input n_2190;
input n_6068;
input n_3438;
input n_166;
input n_4141;
input n_5193;
input n_2850;
input n_572;
input n_1481;
input n_1441;
input n_3373;
input n_5789;
input n_92;
input n_2104;
input n_513;
input n_3883;
input n_5961;
input n_261;
input n_5866;
input n_3728;
input n_2925;
input n_4499;
input n_121;
input n_5822;
input n_433;
input n_5195;
input n_3949;
input n_5726;
input n_2792;
input n_219;
input n_5364;
input n_3315;
input n_263;
input n_5533;
input n_3798;
input n_788;
input n_1543;
input n_1599;
input n_329;
input n_4257;
input n_4458;
input n_2674;
input n_5103;
input n_4641;
input n_4720;
input n_4893;
input n_61;
input n_3857;
input n_1876;
input n_4107;
input n_243;
input n_1873;
input n_3630;
input n_3518;
input n_1866;
input n_117;
input n_2130;
input n_1330;
input n_1413;
input n_3714;
input n_2228;
input n_5039;
input n_2455;
input n_2876;
input n_4772;
input n_5953;
input n_3099;
input n_5198;
input n_4468;
input n_5718;
input n_4161;
input n_1663;
input n_4172;
input n_3403;
input n_2714;
input n_2245;
input n_4961;
input n_4454;
input n_1107;
input n_2457;
input n_3294;
input n_4119;
input n_6001;
input n_3686;
input n_4502;
input n_5958;
input n_318;
input n_2971;
input n_1713;
input n_715;
input n_4277;
input n_4526;
input n_1265;
input n_3490;
input n_4849;
input n_530;
input n_277;
input n_4319;
input n_3369;
input n_618;
input n_199;
input n_5792;
input n_3581;
input n_3069;
input n_6023;
input n_2028;
input n_3715;
input n_1069;
input n_612;
input n_3725;
input n_3933;
input n_5554;
input n_1175;
input n_2311;
input n_429;
input n_1012;
input n_3691;
input n_5553;
input n_4485;
input n_4066;
input n_903;
input n_4146;
input n_5711;
input n_1802;
input n_1504;
input n_4340;
input n_5790;
input n_286;
input n_254;
input n_3961;
input n_4855;
input n_1801;
input n_2347;
input n_3917;
input n_47;
input n_816;
input n_1188;
input n_2206;
input n_4004;
input n_2967;
input n_5404;
input n_2916;
input n_5739;
input n_4292;
input n_5972;
input n_2467;
input n_5549;
input n_267;
input n_3145;
input n_1124;
input n_1624;
input n_3983;
input n_4940;
input n_5444;
input n_3538;
input n_3280;
input n_5757;
input n_1515;
input n_961;
input n_4356;
input n_3510;
input n_2824;
input n_593;
input n_637;
input n_2377;
input n_701;
input n_950;
input n_3009;
input n_5824;
input n_3719;
input n_2525;
input n_4361;
input n_5488;
input n_3827;
input n_891;
input n_5154;
input n_2067;
input n_3889;
input n_2687;
input n_1630;
input n_2887;
input n_4245;
input n_4136;
input n_3526;
input n_2194;
input n_2619;
input n_5329;
input n_4367;
input n_5637;
input n_1987;
input n_507;
input n_968;
input n_2271;
input n_1008;
input n_2583;
input n_4560;
input n_2606;
input n_4899;
input n_5728;
input n_5471;
input n_1033;
input n_462;
input n_1052;
input n_2794;
input n_5164;
input n_2391;
input n_304;
input n_2431;
input n_5843;
input n_125;
input n_2078;
input n_2932;
input n_1767;
input n_3431;
input n_3450;
input n_449;
input n_4663;
input n_2893;
input n_1208;
input n_5484;
input n_2954;
input n_2728;
input n_1072;
input n_815;
input n_3421;
input n_3183;
input n_2493;
input n_4802;
input n_2705;
input n_5523;
input n_1067;
input n_3405;
input n_5423;
input n_255;
input n_284;
input n_1952;
input n_5074;
input n_4044;
input n_3436;
input n_1026;
input n_1880;
input n_3442;
input n_3366;
input n_2631;
input n_38;
input n_289;
input n_3937;
input n_1293;
input n_3159;
input n_4701;
input n_108;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_3240;
input n_3576;
input n_1863;
input n_3385;
input n_4851;
input n_3293;
input n_872;
input n_3922;
input n_86;
input n_5204;
input n_5333;
input n_847;
input n_644;
input n_682;
input n_851;
input n_4991;
input n_5594;
input n_72;
input n_2554;
input n_5422;
input n_1513;
input n_1913;
input n_4934;
input n_837;
input n_5087;
input n_5526;
input n_5292;
input n_2517;
input n_2713;
input n_5000;
input n_2765;
input n_5403;
input n_2590;
input n_5551;
input n_3150;
input n_2060;
input n_4479;
input n_2608;
input n_4011;
input n_5131;
input n_1959;
input n_3133;
input n_5257;
input n_765;
input n_1492;
input n_1340;
input n_4688;
input n_4753;
input n_4058;
input n_631;
input n_2262;
input n_3611;
input n_3082;
input n_4848;
input n_5059;
input n_156;
input n_5887;
input n_843;
input n_2604;
input n_2407;
input n_1277;
input n_2816;
input n_3799;
input n_2574;
input n_4475;
input n_5242;
input n_5219;
input n_2675;
input n_5631;
input n_3537;
input n_4443;
input n_3887;
input n_6008;
input n_1022;
input n_614;
input n_5854;
input n_2667;
input n_5460;
input n_4587;
input n_1615;
input n_4114;
input n_1474;
input n_1571;
input n_2948;
input n_1577;
input n_2119;
input n_947;
input n_1117;
input n_1992;
input n_5686;
input n_5899;
input n_3223;
input n_3140;
input n_3185;
input n_4749;
input n_2605;
input n_5155;
input n_118;
input n_926;
input n_3654;
input n_1849;
input n_2848;
input n_919;
input n_1698;
input n_4100;
input n_4264;
input n_5981;
input n_3788;
input n_89;
input n_4891;
input n_5937;
input n_777;
input n_1299;
input n_5339;
input n_3837;
input n_2718;
input n_1436;
input n_1384;
input n_3325;
input n_2238;
input n_6040;
input n_4085;
input n_4464;
input n_4624;
input n_4818;
input n_4659;
input n_3600;
input n_18;
input n_5217;
input n_5465;
input n_5015;
input n_4339;
input n_1178;
input n_98;
input n_2338;
input n_3324;
input n_796;
input n_1195;
input n_184;
input n_1811;
input n_1857;
input n_3987;
input n_1519;
input n_6039;
input n_2144;
input n_1284;
input n_1604;
input n_4487;
input n_4889;
input n_4866;
input n_1142;
input n_623;
input n_1048;
input n_5721;
input n_3638;
input n_4816;
input n_2110;
input n_5719;
input n_1502;
input n_5773;
input n_1659;
input n_5482;
input n_3393;
input n_6012;
input n_3451;
input n_1418;
input n_1250;
input n_292;
input n_4937;
input n_5277;
input n_3615;
input n_3072;
input n_3087;
input n_2053;
input n_2259;
input n_2121;
input n_4222;
input n_4874;
input n_4401;
input n_889;
input n_2710;
input n_6064;
input n_3142;
input n_4015;
input n_1966;
input n_5793;
input n_477;
input n_1110;
input n_4709;
input n_2213;
input n_4976;
input n_2389;
input n_2132;
input n_2892;
input n_4120;
input n_1564;
input n_5578;
input n_4658;
input n_231;
input n_2860;
input n_2330;
input n_40;
input n_5296;
input n_1457;
input n_505;
input n_3718;
input n_5893;
input n_1787;
input n_537;
input n_1993;
input n_2281;
input n_2617;
input n_2776;
input n_1466;
input n_10;
input n_1919;
input n_5742;
input n_5207;
input n_3705;
input n_3211;
input n_3909;
input n_5676;
input n_546;
input n_386;
input n_1220;
input n_6051;
input n_1893;
input n_2301;
input n_4665;
input n_3582;
input n_4223;
input n_2387;
input n_5674;
input n_3270;
input n_5539;
input n_2846;
input n_5282;
input n_970;
input n_2488;
input n_1980;
input n_5464;
input n_2237;
input n_1060;
input n_1951;
input n_444;
input n_4362;
input n_1252;
input n_3311;
input n_3913;
input n_1223;
input n_511;
input n_5121;
input n_6026;
input n_6070;
input n_1286;
input n_2115;
input n_4430;
input n_3302;
input n_4348;
input n_5013;
input n_1597;
input n_4489;
input n_4839;
input n_2596;
input n_3163;
input n_775;
input n_4404;
input n_1153;
input n_5589;
input n_439;
input n_1531;
input n_2828;
input n_453;
input n_2384;
input n_4261;
input n_4204;
input n_759;
input n_2724;
input n_426;
input n_2585;
input n_5628;
input n_4825;
input n_2352;
input n_1625;
input n_3986;
input n_5006;
input n_4513;
input n_4006;
input n_2226;
input n_2801;
input n_1901;
input n_3869;
input n_2556;
input n_4747;
input n_1647;
input n_5251;
input n_3753;
input n_2306;
input n_1614;
input n_1892;
input n_3742;
input n_3683;
input n_4801;
input n_401;
input n_3260;
input n_2550;
input n_3175;
input n_3736;
input n_5475;
input n_5807;
input n_4448;
input n_1096;
input n_2227;
input n_5216;
input n_3284;
input n_4869;
input n_427;
input n_2159;
input n_4386;
input n_688;
input n_1077;
input n_2315;
input n_4132;
input n_2995;
input n_5273;
input n_1437;
input n_4844;
input n_4438;
input n_4836;
input n_5439;
input n_4955;
input n_4149;
input n_5936;
input n_4355;
input n_501;
input n_2276;
input n_3234;
input n_856;
input n_2803;
input n_379;
input n_1668;
input n_2777;
input n_3202;
input n_2830;
input n_3220;
input n_1129;
input n_602;
input n_2181;
input n_6069;
input n_171;
input n_2911;
input n_169;
input n_4655;
input n_1429;
input n_5706;
input n_2826;
input n_3429;
input n_2379;
input n_326;
input n_587;
input n_3554;
input n_1593;
input n_1202;
input n_1635;
input n_5431;
input n_4067;
input n_4357;
input n_28;
input n_3462;
input n_2851;
input n_4374;
input n_5132;
input n_106;
input n_358;
input n_160;
input n_2420;
input n_5627;
input n_5774;
input n_3722;
input n_186;
input n_4400;
input n_4846;
input n_5798;
input n_2984;
input n_575;
input n_5187;
input n_5875;
input n_4024;
input n_1508;
input n_5621;
input n_5608;
input n_732;
input n_2983;
input n_2240;
input n_392;
input n_2538;
input n_724;
input n_3250;
input n_1042;
input n_4582;
input n_1728;
input n_557;
input n_1871;
input n_4860;
input n_845;
input n_140;
input n_5844;
input n_3414;
input n_1549;
input n_4870;
input n_768;
input n_3651;
input n_2102;
input n_2563;
input n_4989;
input n_3449;
input n_1683;
input n_1916;
input n_2598;
input n_597;
input n_280;
input n_1187;
input n_4304;
input n_4558;
input n_1403;
input n_4488;
input n_3767;
input n_2544;
input n_3550;
input n_4211;
input n_1206;
input n_4016;
input n_5867;
input n_621;
input n_750;
input n_5508;
input n_4656;
input n_3839;
input n_2823;
input n_5597;
input n_4915;
input n_4328;
input n_1057;
input n_2785;
input n_235;
input n_5515;
input n_1997;
input n_5662;
input n_2636;
input n_3131;
input n_710;
input n_1818;
input n_3730;
input n_1298;
input n_5862;
input n_4397;
input n_3399;
input n_2088;
input n_1611;
input n_5050;
input n_2740;
input n_746;
input n_4808;
input n_5697;
input n_3416;
input n_3498;
input n_5767;
input n_2401;
input n_101;
input n_1589;
input n_4712;
input n_2309;
input n_2900;
input n_2957;
input n_1740;
input n_2737;
input n_3994;
input n_5462;
input n_1497;
input n_133;
input n_5980;
input n_3672;
input n_5318;
input n_3533;
input n_1622;
input n_4725;
input n_6022;
input n_4406;
input n_1694;
input n_1535;
input n_3382;
input n_3132;
input n_5498;
input n_2571;
input n_3138;
input n_20;
input n_5053;
input n_2171;
input n_2988;
input n_4908;
input n_3136;
input n_1350;
input n_4109;
input n_4192;
input n_4824;
input n_2037;
input n_2808;
input n_4567;
input n_5150;
input n_782;
input n_809;
input n_3819;
input n_4778;
input n_5477;
input n_1797;
input n_5175;
input n_986;
input n_2050;
input n_4595;
input n_2164;
input n_4174;
input n_402;
input n_1870;
input n_1171;
input n_460;
input n_5987;
input n_5179;
input n_1827;
input n_4904;
input n_2187;
input n_1152;
input n_450;
input n_3544;
input n_4150;
input n_2904;
input n_5988;
input n_5585;
input n_6058;
input n_711;
input n_3105;
input n_2872;
input n_3692;
input n_4616;
input n_4982;
input n_370;
input n_1695;
input n_2046;
input n_2272;
input n_2760;
input n_1979;
input n_4643;
input n_2738;
input n_972;
input n_5348;
input n_1332;
input n_5480;
input n_4323;
input n_624;
input n_2346;
input n_4831;
input n_936;
input n_3045;
input n_3821;
input n_885;
input n_83;
input n_2342;
input n_2167;
input n_2970;
input n_3676;
input n_4896;
input n_2882;
input n_3666;
input n_3675;
input n_4017;
input n_4260;
input n_4916;
input n_2541;
input n_2940;
input n_5904;
input n_4739;
input n_599;
input n_6062;
input n_105;
input n_1974;
input n_4122;
input n_934;
input n_4209;
input n_2768;
input n_3858;
input n_1341;
input n_5284;
input n_4298;
input n_2314;
input n_3502;
input n_5461;
input n_3003;
input n_4128;
input n_543;
input n_5147;
input n_4271;
input n_4644;
input n_1355;
input n_2258;
input n_5503;
input n_325;
input n_5845;
input n_5945;
input n_804;
input n_2390;
input n_959;
input n_2562;
input n_4716;
input n_4312;
input n_1343;
input n_1522;
input n_76;
input n_2734;
input n_1782;
input n_5600;
input n_5755;
input n_707;
input n_1900;
input n_5048;
input n_6053;
input n_3246;
input n_1548;
input n_3381;
input n_1155;
input n_2195;
input n_3208;
input n_4944;
input n_5245;
input n_4343;
input n_4715;
input n_4935;
input n_4694;
input n_4672;
input n_5054;
input n_2962;
input n_5448;
input n_2939;
input n_5749;
input n_1672;
input n_1925;
input n_4407;
input n_737;
input n_4045;
input n_3517;
input n_2945;
input n_4598;
input n_3061;
input n_3893;
input n_3932;
input n_21;
input n_3469;
input n_2960;
input n_5993;
input n_138;
input n_3258;
input n_4524;
input n_3143;
input n_6020;
input n_333;
input n_4084;
input n_3149;
input n_3365;
input n_3379;
input n_24;
input n_459;
input n_4850;
input n_4424;
input n_3008;
input n_1751;
input n_2840;
input n_285;
input n_3939;
input n_4776;
input n_1375;
input n_3972;
input n_4153;
input n_85;
input n_3506;
input n_1650;
input n_1962;
input n_3855;
input n_1928;
input n_3091;
input n_4317;
input n_4723;
input n_4269;
input n_5418;
input n_4088;
input n_3398;
input n_5685;
input n_2761;
input n_2793;
input n_3776;
input n_3711;
input n_4235;
input n_5459;
input n_1019;
input n_4143;
input n_4170;
input n_729;
input n_876;
input n_774;
input n_3642;
input n_2845;
input n_4650;
input n_438;
input n_4719;
input n_5173;
input n_1860;
input n_5016;
input n_1904;
input n_2874;
input n_1200;
input n_2588;
input n_479;
input n_1353;
input n_1777;
input n_4967;
input n_3308;
input n_1113;
input n_1600;
input n_2253;
input n_2366;
input n_4912;
input n_4799;
input n_2261;
input n_4423;
input n_5086;
input n_5283;
input n_2210;
input n_4735;
input n_3602;
input n_187;
input n_3300;
input n_2978;
input n_2516;
input n_1050;
input n_1411;
input n_5170;
input n_2827;
input n_1177;
input n_3515;
input n_1150;
input n_566;
input n_1023;
input n_2951;
input n_1118;
input n_194;
input n_2949;
input n_1807;
input n_5028;
input n_5839;
input n_1814;
input n_1631;
input n_1879;
input n_256;
input n_440;
input n_3806;
input n_5514;
input n_2931;
input n_209;
input n_367;
input n_2569;
input n_3866;
input n_5351;
input n_5909;
input n_671;
input n_4543;
input n_740;
input n_703;
input n_4157;
input n_4229;
input n_5293;
input n_3865;
input n_4073;
input n_1324;
input n_3629;
input n_1435;
input n_5400;
input n_3920;
input n_969;
input n_4892;
input n_3255;
input n_1401;
input n_1516;
input n_3846;
input n_180;
input n_3512;
input n_5201;
input n_2029;
input n_5890;
input n_4439;
input n_1394;
input n_1326;
input n_4783;
input n_1379;
input n_214;
input n_935;
input n_4910;
input n_1130;
input n_3083;
input n_676;
input n_832;
input n_3049;
input n_5389;
input n_5142;
input n_3830;
input n_3679;
input n_5891;
input n_3541;
input n_74;
input n_3117;
input n_5935;
input n_4930;
input n_372;
input n_111;
input n_314;
input n_378;
input n_5623;
input n_338;
input n_1283;
input n_2385;
input n_4112;
input n_506;
input n_360;
input n_2149;
input n_2396;
input n_4557;
input n_4917;
input n_895;
input n_2450;
input n_3739;
input n_4432;
input n_2284;
input n_4352;
input n_4416;
input n_4593;
input n_344;
input n_2769;
input n_4465;
input n_3622;
input n_5114;
input n_4980;
input n_1392;
input n_5693;
input n_4495;
input n_5117;
input n_1924;
input n_5663;
input n_525;
input n_2463;
input n_3363;
input n_1677;
input n_5990;
input n_611;
input n_3721;
input n_3062;
input n_2679;
input n_5024;
input n_4559;
input n_838;
input n_3969;
input n_129;
input n_3336;
input n_4160;
input n_4231;
input n_2952;
input n_5647;
input n_1017;
input n_4256;
input n_2779;
input n_4938;
input n_5396;
input n_5203;
input n_109;
input n_445;
input n_930;
input n_2620;
input n_5162;
input n_1945;
input n_5426;
input n_1656;
input n_5803;
input n_2112;
input n_1464;
input n_2430;
input n_653;
input n_1414;
input n_5285;
input n_2721;
input n_944;
input n_4335;
input n_2034;
input n_576;
input n_270;
input n_2683;
input n_563;
input n_5365;
input n_2744;
input n_1011;
input n_4521;
input n_1566;
input n_626;
input n_990;
input n_3204;
input n_1104;
input n_5715;
input n_4920;
input n_498;
input n_870;
input n_5395;
input n_1253;
input n_366;
input n_5709;
input n_1693;
input n_3256;
input n_348;
input n_3802;
input n_376;
input n_2118;
input n_2111;
input n_390;
input n_2915;
input n_1148;
input n_2188;
input n_1989;
input n_2802;
input n_3643;
input n_2425;
input n_4265;
input n_2950;
input n_5634;
input n_5672;
input n_719;
input n_3060;
input n_3098;
input n_4105;
input n_1851;
input n_1090;
input n_4861;
input n_5799;
input n_4064;
input n_4926;
input n_1518;
input n_1362;
input n_3123;
input n_3380;
input n_5617;
input n_1829;
input n_5266;
input n_5580;
input n_1450;
input n_4828;
input n_1638;
input n_3038;
input n_570;
input n_1789;
input n_620;
input n_519;
input n_2523;
input n_5450;
input n_2413;
input n_3769;
input n_1482;
input n_5310;
input n_3863;
input n_3669;
input n_3130;
input n_4316;
input n_5722;
input n_4640;
input n_5122;
input n_5390;
input n_1710;
input n_2161;
input n_1301;
input n_2805;
input n_5593;
input n_33;
input n_4769;
input n_5764;
input n_2282;
input n_4628;
input n_2047;
input n_5385;
input n_1609;
input n_3344;
input n_5237;
input n_2334;
input n_5133;
input n_409;
input n_1763;
input n_5322;
input n_3989;
input n_2490;
input n_4460;
input n_4108;
input n_635;
input n_3786;
input n_3841;
input n_4254;
input n_1996;
input n_2867;
input n_1442;
input n_2726;
input n_4303;
input n_5853;
input n_5982;
input n_1158;
input n_2248;
input n_5011;
input n_5917;
input n_2662;
input n_4909;
input n_3147;
input n_753;
input n_3925;
input n_3180;
input n_2795;
input n_3472;
input n_5376;
input n_5106;
input n_269;
input n_359;
input n_1479;
input n_4768;
input n_1675;
input n_3717;
input n_5561;
input n_5410;
input n_571;
input n_2215;
input n_404;
input n_158;
input n_1884;
input n_665;
input n_2055;
input n_5156;
input n_2553;
input n_149;
input n_632;
input n_2038;
input n_4447;
input n_4826;
input n_3445;
input n_373;
input n_87;
input n_1833;
input n_3903;
input n_5998;
input n_1494;
input n_2325;
input n_1850;
input n_5304;
input n_3854;
input n_3235;
input n_5378;
input n_6028;
input n_1417;
input n_3673;
input n_4281;
input n_5916;
input n_681;
input n_4648;
input n_3094;
input n_412;
input n_965;
input n_1428;
input n_1576;
input n_1856;
input n_2077;
input n_5691;
input n_1059;
input n_4951;
input n_422;
input n_4957;
input n_3079;
input n_165;
input n_4360;
input n_540;
input n_4039;
input n_457;
input n_3070;
input n_3800;
input n_4566;
input n_3263;
input n_4853;
input n_1748;
input n_3504;
input n_531;
input n_4272;
input n_2930;
input n_5615;
input n_1025;
input n_3111;
input n_336;
input n_12;
input n_1885;
input n_5269;
input n_3054;
input n_1538;
input n_1240;
input n_5468;
input n_1;
input n_4730;
input n_5399;
input n_1234;
input n_5262;
input n_3254;
input n_3684;
input n_4670;
input n_4882;
input n_4620;
input n_3152;
input n_4738;
input n_3579;
input n_5421;
input n_3335;
input n_4177;
input n_3783;
input n_700;
input n_1307;
input n_3178;
input n_4127;
input n_5206;
input n_1003;
input n_5713;
input n_5256;
input n_168;
input n_2353;
input n_4099;
input n_4517;
input n_77;
input n_4168;
input n_5188;
input n_1738;
input n_4490;
input n_1575;
input n_1923;
input n_2260;
input n_3952;
input n_5550;
input n_3911;
input n_1688;
input n_4285;
input n_3465;
input n_1743;
input n_2997;
input n_1991;
input n_2386;
input n_5161;
input n_5373;
input n_1724;
input n_3708;
input n_4078;
input n_3046;
input n_2956;
input n_5573;
input n_1553;
input n_5939;
input n_5509;
input n_5382;
input n_5659;
input n_3619;
input n_1415;
input n_5881;
input n_1370;
input n_1786;
input n_4198;
input n_2382;
input n_3754;
input n_2291;
input n_415;
input n_1371;
input n_383;
input n_2886;
input n_2974;
input n_4213;
input n_200;
input n_2184;
input n_2982;
input n_1803;
input n_4065;
input n_5863;
input n_229;
input n_2645;
input n_3904;
input n_1393;
input n_1517;
input n_1867;
input n_2630;
input n_1444;
input n_1603;
input n_2470;
input n_4446;
input n_1263;
input n_4417;
input n_5466;
input n_4733;
input n_4764;
input n_1261;
input n_3879;
input n_2286;
input n_4743;
input n_2018;
input n_3080;
input n_1903;
input n_1143;
input n_5955;
input n_658;
input n_1874;
input n_2865;
input n_2825;
input n_2013;
input n_2044;
input n_3023;
input n_3232;
input n_693;
input n_1056;
input n_758;
input n_5851;
input n_2256;
input n_943;
input n_4060;
input n_5110;
input n_4879;
input n_5796;
input n_42;
input n_772;
input n_2806;
input n_770;
input n_3028;
input n_3662;
input n_2981;
input n_3076;
input n_886;
input n_343;
input n_3624;
input n_1345;
input n_1820;
input n_4556;
input n_539;
input n_45;
input n_4117;
input n_4687;
input n_2836;
input n_638;
input n_1404;
input n_5492;
input n_5995;
input n_2378;
input n_887;
input n_5905;
input n_2655;
input n_4600;
input n_126;
input n_1467;
input n_4250;
input n_5829;
input n_3906;
input n_224;
input n_4954;
input n_5191;
input n_1231;
input n_2599;
input n_3963;
input n_3368;
input n_9;
input n_2370;
input n_2612;
input n_2591;
input n_4881;
input n_1815;
input n_2214;
input n_4253;
input n_407;
input n_913;
input n_5734;
input n_2593;
input n_4255;
input n_867;
input n_4071;
input n_3568;
input n_1230;
input n_3850;
input n_5770;
input n_1333;
input n_2496;
input n_5705;
input n_3313;
input n_4605;
input n_3189;
input n_5525;
input n_163;
input n_1644;
input n_2725;
input n_2277;
input n_4691;
input n_1558;
input n_1732;
input n_2300;
input n_3943;
input n_4305;
input n_824;
input n_4297;
input n_6052;
input n_2907;
input n_577;
input n_5374;
input n_5575;
input n_1843;
input n_619;
input n_5675;
input n_4227;
input n_521;
input n_2778;
input n_395;
input n_1909;
input n_5020;
input n_606;
input n_5297;
input n_1123;
input n_1309;
input n_2961;
input n_916;
input n_3934;
input n_4033;
input n_4415;
input n_483;
input n_1970;
input n_630;
input n_2059;
input n_2669;
input n_4094;
input n_4765;
input n_2546;
input n_3193;
input n_2522;
input n_476;
input n_4364;
input n_1957;
input n_4354;
input n_4732;
input n_3912;
input n_3118;
input n_5959;
input n_3720;
input n_1907;
input n_2529;
input n_264;
input n_860;
input n_1530;
input n_4745;
input n_938;
input n_1302;
input n_5642;
input n_4581;
input n_549;
input n_4377;
input n_2143;
input n_905;
input n_4792;
input n_1680;
input n_3842;
input n_322;
input n_993;
input n_689;
input n_2031;
input n_4878;
input n_1605;
input n_3514;
input n_4979;
input n_1988;
input n_558;
input n_2654;
input n_3036;
input n_5302;
input n_966;
input n_4511;
input n_2908;
input n_3357;
input n_692;
input n_5639;
input n_5781;
input n_1233;
input n_3895;
input n_487;
input n_241;
input n_4520;
input n_5299;
input n_3455;
input n_4118;
input n_4503;
input n_2176;
input n_2459;
input n_1111;
input n_3599;
input n_5543;
input n_1251;
input n_5361;
input n_2711;
input n_4199;
input n_5885;
input n_1912;
input n_5356;
input n_4441;
input n_1982;
input n_3872;
input n_3772;
input n_5458;
input n_1312;
input n_5668;
input n_5038;
input n_268;
input n_1760;
input n_5330;
input n_4585;
input n_2664;
input n_5;
input n_1664;
input n_1722;
input n_5463;
input n_3022;
input n_247;
input n_5489;
input n_1165;
input n_5892;
input n_4773;
input n_5654;
input n_2008;
input n_6009;
input n_2192;
input n_3281;
input n_2345;
input n_328;
input n_1386;
input n_4427;
input n_5923;
input n_5113;
input n_5479;
input n_3549;
input n_5714;
input n_2804;
input n_2453;
input n_2676;
input n_5510;
input n_3940;
input n_4822;
input n_1214;
input n_690;
input n_850;
input n_5692;
input n_4800;
input n_1157;
input n_3453;
input n_5555;
input n_3410;
input n_1752;
input n_1813;
input n_3768;
input n_4958;
input n_2810;
input n_4043;
input n_2319;
input n_5441;
input n_825;
input n_6066;
input n_3785;
input n_2963;
input n_5366;
input n_2602;
input n_55;
input n_3873;
input n_2980;
input n_696;
input n_4886;
input n_1082;
input n_1317;
input n_3227;
input n_2733;
input n_3289;
input n_4055;
input n_2178;
input n_5968;
input n_2644;
input n_2036;
input n_3326;
input n_4200;
input n_3460;
input n_2411;
input n_1796;
input n_2082;
input n_3519;
input n_678;
input n_5078;
input n_3707;
input n_283;
input n_3578;
input n_909;
input n_4737;
input n_590;
input n_4925;
input n_4116;
input n_5415;
input n_362;
input n_22;
input n_5419;
input n_1990;
input n_3805;
input n_2943;
input n_5205;
input n_1634;
input n_3252;
input n_627;
input n_3253;
input n_1465;
input n_342;
input n_2622;
input n_2658;
input n_2665;
input n_2133;
input n_1712;
input n_4603;
input n_1523;
input n_1627;
input n_5080;
input n_5976;
input n_3128;
input n_1527;
input n_495;
input n_5732;
input n_5372;
input n_2691;
input n_840;
input n_2913;
input n_4471;
input n_2230;
input n_1969;
input n_2690;
input n_5208;
input n_1565;
input n_1493;
input n_5690;
input n_2573;
input n_2646;
input n_2535;
input n_1364;
input n_3078;
input n_2436;
input n_615;
input n_3838;
input n_5371;
input n_4651;
input n_3941;
input n_3793;
input n_4854;
input n_5071;
input n_3789;
input n_605;
input n_1514;
input n_5801;
input n_6047;
input n_3037;
input n_1646;
input n_3729;
input n_4994;
input n_2537;
input n_4483;
input n_5347;
input n_5168;
input n_4661;
input n_1308;
input n_4988;
input n_3171;
input n_3608;
input n_4540;
input n_2097;
input n_79;
input n_3459;
input n_2853;
input n_1808;
input n_3053;
input n_3358;
input n_6021;
input n_3499;
input n_4284;
input n_1005;
input n_1947;
input n_3426;
input n_4971;
input n_5656;
input n_1469;
input n_5125;
input n_5857;
input n_2650;
input n_5652;
input n_987;
input n_5499;
input n_720;
input n_153;
input n_3229;
input n_3348;
input n_1707;
input n_656;
input n_5228;
input n_797;
input n_2933;
input n_2717;
input n_1723;
input n_1878;
input n_189;
input n_738;
input n_2012;
input n_3497;
input n_5066;
input n_2842;
input n_3580;
input n_2335;
input n_529;
input n_2307;
input n_3704;
input n_684;
input n_5507;
input n_1809;
input n_5569;
input n_4280;
input n_1181;
input n_37;
input n_5190;
input n_3173;
input n_3677;
input n_3996;
input n_1049;
input n_4097;
input n_1666;
input n_803;
input n_4218;
input n_5392;
input n_1717;
input n_1817;
input n_2449;
input n_3880;
input n_3685;
input n_2868;
input n_2231;
input n_3609;
input n_1228;
input n_5455;
input n_417;
input n_5442;
input n_5948;
input n_4459;
input n_4545;
input n_272;
input n_2896;
input n_3019;
input n_2639;
input n_3471;
input n_5511;
input n_2898;
input n_69;
input n_5295;
input n_2368;
input n_53;
input n_458;
input n_4175;
input n_5490;
input n_16;
input n_3200;
input n_4771;
input n_3259;
input n_2524;
input n_3167;
input n_2460;
input n_5836;
input n_3867;
input n_3593;
input n_4455;
input n_1073;
input n_252;
input n_4514;
input n_5834;
input n_3191;
input n_5584;
input n_4140;
input n_2481;
input n_3561;
input n_4806;
input n_2682;
input n_3032;
input n_5160;
input n_2877;
input n_5098;
input n_1021;
input n_811;
input n_683;
input n_1207;
input n_5707;
input n_5140;
input n_4992;
input n_5197;
input n_5497;
input n_880;
input n_3505;
input n_3540;
input n_3577;
input n_2432;
input n_150;
input n_1478;
input n_4796;
input n_3598;
input n_4442;
input n_2581;
input n_1363;
input n_3641;
input n_3777;
input n_4203;
input n_767;
input n_1837;
input n_2218;
input n_4533;
input n_831;
input n_5481;
input n_3590;
input n_2435;
input n_5344;
input n_954;
input n_4419;
input n_5308;
input n_1410;
input n_5184;
input n_5794;
input n_1382;
input n_5408;
input n_1736;
input n_4053;
input n_1483;
input n_3848;
input n_1372;
input n_3327;
input n_1719;
input n_319;
input n_2701;
input n_2511;
input n_4167;
input n_1427;
input n_2745;
input n_1080;
input n_5271;
input n_123;
input n_562;
input n_5964;
input n_6004;
input n_2323;
input n_2784;
input n_5494;
input n_162;
input n_5234;
input n_4431;
input n_2421;
input n_1136;
input n_4387;
input n_2618;
input n_3265;
input n_2464;
input n_128;
input n_1125;
input n_3755;
input n_4042;
input n_5128;
input n_2224;
input n_2329;
input n_1092;
input n_441;
input n_5467;
input n_4299;
input n_4890;
input n_146;
input n_1784;
input n_3571;
input n_193;
input n_1775;
input n_2410;
input n_1093;
input n_1783;
input n_2929;
input n_4176;
input n_5827;
input n_5199;
input n_296;
input n_651;
input n_3407;
input n_5992;
input n_217;
input n_5313;
input n_1185;
input n_3856;
input n_4236;
input n_3425;
input n_215;
input n_3894;
input n_3127;
input n_1831;
input n_2621;
input n_3623;
input n_5312;
input n_5079;
input n_54;
input n_1453;
input n_2502;
input n_3646;
input n_5513;
input n_5614;
input n_497;
input n_4830;
input n_4706;
input n_1315;
input n_5225;
input n_4570;
input n_2754;
input n_1224;
input n_2783;
input n_3188;
input n_1459;
input n_2462;
input n_3243;
input n_1135;
input n_2889;
input n_4034;
input n_4056;
input n_4622;
input n_3960;
input n_1470;
input n_4887;
input n_2732;
input n_4693;
input n_4206;
input n_2249;
input n_1091;
input n_2000;
input n_3862;
input n_4267;
input n_5835;
input n_2270;
input n_1425;
input n_5049;
input n_983;
input n_5846;
input n_906;
input n_1390;
input n_2289;
input n_1733;
input n_2955;
input n_5592;
input n_2158;
input n_4609;
input n_1855;
input n_3051;
input n_3367;
input n_385;
input n_1687;
input n_1439;
input n_2328;
input n_2859;
input n_2202;
input n_1331;
input n_613;
input n_736;
input n_5278;
input n_3314;
input n_3525;
input n_2100;
input n_5157;
input n_2993;
input n_4754;
input n_3016;
input n_4647;
input n_1134;
input n_3688;
input n_4003;
input n_5708;
input n_554;
input n_1995;
input n_3751;
input n_5223;
input n_4894;
input n_5474;
input n_4113;
input n_1889;
input n_4760;
input n_5649;
input n_435;
input n_1905;
input n_3466;
input n_762;
input n_5704;
input n_4983;
input n_1778;
input n_5956;
input n_5287;
input n_1079;
input n_2139;
input n_419;
input n_5083;
input n_4509;
input n_6007;
input n_2875;
input n_1103;
input n_3907;
input n_3338;
input n_144;
input n_4217;
input n_4906;
input n_2219;
input n_1203;
input n_3636;
input n_2327;
input n_999;
input n_5516;
input n_1254;
input n_2841;
input n_4897;
input n_3539;
input n_3291;
input n_4399;
input n_2304;
input n_2487;
input n_5698;
input n_3276;
input n_2597;
input n_3194;
input n_5084;
input n_5771;
input n_3572;
input n_349;
input n_3886;
input n_4710;
input n_4420;
input n_443;
input n_892;
input n_3637;
input n_4574;
input n_1468;
input n_2855;
input n_1859;
input n_2156;
input n_1718;
input n_5174;
input n_4234;
input n_5538;
input n_4101;
input n_3548;
input n_5017;
input n_1768;
input n_3974;
input n_198;
input n_1847;
input n_3634;
input n_1397;
input n_3236;
input n_901;
input n_2755;
input n_3141;
input n_923;
input n_5096;
input n_1841;
input n_4660;
input n_5241;
input n_1623;
input n_1015;
input n_3112;
input n_4797;
input n_3108;
input n_4270;
input n_5428;
input n_4151;
input n_4945;
input n_3417;
input n_5677;
input n_4124;
input n_5570;
input n_73;
input n_785;
input n_5153;
input n_609;
input n_4611;
input n_5927;
input n_5435;
input n_2337;
input n_1356;
input n_3213;
input n_4333;
input n_127;
input n_3820;
input n_5200;
input n_2607;
input n_2890;
input n_1168;
input n_5115;
input n_1943;
input n_5566;
input n_3249;
input n_1320;
input n_2722;
input n_1452;
input n_2854;
input n_2499;
input n_4152;
input n_5487;
input n_302;
input n_5486;
input n_137;
input n_1596;
input n_5092;
input n_5244;
input n_1734;
input n_3172;
input n_4832;
input n_2902;
input n_5889;
input n_3217;
input n_1983;
input n_5391;
input n_1938;
input n_2472;
input n_3394;
input n_1715;
input n_3536;
input n_1443;
input n_1272;
input n_2894;
input n_3957;
input n_3710;
input n_4195;
input n_5849;
input n_4554;
input n_3040;
input n_3279;
input n_5240;
input n_2402;
input n_2225;
input n_1081;
input n_5951;
input n_1692;
input n_1084;
input n_5912;
input n_1864;
input n_2006;
input n_3402;
input n_3475;
input n_3501;
input n_374;
input n_1705;
input n_3905;
input n_4680;
input n_3013;
input n_921;
input n_579;
input n_2789;
input n_5152;
input n_5265;
input n_2257;
input n_4927;
input n_5574;
input n_4258;
input n_1828;
input n_2699;
input n_2200;
input n_650;
input n_1940;
input n_4548;
input n_4862;
input n_1405;
input n_2376;
input n_5469;
input n_456;
input n_3878;
input n_2670;
input n_313;
input n_2700;
input n_5910;
input n_5895;
input n_1041;
input n_5804;
input n_565;
input n_3134;
input n_5965;
input n_1569;
input n_3115;
input n_1062;
input n_896;
input n_4553;
input n_3278;
input n_2084;
input n_4875;
input n_5682;
input n_5387;
input n_654;
input n_5557;
input n_411;
input n_2458;
input n_1222;
input n_3050;
input n_2673;
input n_2456;
input n_2527;
input n_2635;
input n_1637;
input n_3307;
input n_1407;
input n_1795;
input n_2871;
input n_420;
input n_4321;
input n_4183;
input n_164;
input n_5681;
input n_1271;
input n_4901;
input n_1545;
input n_4821;
input n_4145;
input n_3121;
input n_1640;
input n_4040;
input n_2406;
input n_806;
input n_584;
input n_2141;
input n_5316;
input n_244;
input n_548;
input n_282;
input n_5703;
input n_833;
input n_523;
input n_345;
input n_3930;
input n_4943;
input n_799;
input n_3044;
input n_4757;
input n_2196;
input n_2629;
input n_2809;
input n_787;
input n_2172;
input n_4682;
input n_5564;
input n_5620;
input n_4530;
input n_1528;
input n_1146;
input n_2021;
input n_4942;
input n_159;
input n_1086;
input n_5406;
input n_2125;
input n_2561;
input n_652;
input n_4604;
input n_1906;
input n_3305;
input n_2992;
input n_5724;
input n_1241;
input n_3157;
input n_4841;
input n_1758;
input n_3221;
input n_3267;
input n_2422;
input n_1914;
input n_1318;
input n_5806;
input n_4338;
input n_3457;
input n_306;
input n_3762;
input n_5738;
input n_3005;
input n_3151;
input n_3411;
input n_4840;
input n_1029;
input n_4519;
input n_3779;
input n_2388;
input n_5355;
input n_3984;
input n_5320;
input n_5353;
input n_1706;
input n_5186;
input n_5710;
input n_1498;
input n_2417;
input n_1210;
input n_5093;
input n_1556;
input n_4052;
input n_5979;
input n_3558;
input n_1984;
input n_2236;
input n_5438;
input n_6044;
input n_4326;
input n_1269;
input n_2083;
input n_2834;
input n_5517;
input n_3207;
input n_5605;
input n_2441;
input n_3401;
input n_3242;
input n_3613;
input n_655;
input n_4726;
input n_1045;
input n_5907;
input n_786;
input n_1559;
input n_6045;
input n_1872;
input n_19;
input n_29;
input n_75;
input n_5040;
input n_6063;
input n_1325;
input n_3761;
input n_4315;
input n_2888;
input n_2923;
input n_1727;
input n_4301;
input n_151;
input n_3744;
input n_4788;
input n_2041;
input n_1360;
input n_5977;
input n_3814;
input n_3781;
input n_1908;
input n_2484;
input n_2126;
input n_6003;
input n_3843;
input n_1098;
input n_5746;
input n_2045;
input n_817;
input n_5451;
input n_3687;
input n_2216;
input n_5402;
input n_3543;
input n_3621;
input n_6031;
input n_2903;
input n_3216;
input n_332;
input n_3808;
input n_398;
input n_4365;
input n_6060;
input n_1882;
input n_3726;
input n_1007;
input n_1929;
input n_2369;
input n_1592;
input n_2719;
input n_591;
input n_3758;
input n_5417;
input n_2587;
input n_3199;
input n_680;
input n_3339;
input n_4923;
input n_2400;
input n_5864;
input n_1953;
input n_4741;
input n_3343;
input n_2752;
input n_4885;
input n_751;
input n_5432;
input n_1399;
input n_4550;
input n_4652;
input n_2358;
input n_5453;
input n_3658;
input n_4900;
input n_2163;
input n_2186;
input n_2815;
input n_3034;
input n_4408;
input n_4577;
input n_4748;
input n_643;
input n_5842;
input n_400;
input n_337;
input n_5814;
input n_2814;
input n_5253;
input n_5209;
input n_789;
input n_3231;
input n_4212;
input n_2979;
input n_5699;
input n_181;
input n_5531;
input n_5765;
input n_2953;
input n_327;
input n_4295;
input n_5943;
input n_2946;
input n_2500;
input n_3430;
input n_2269;
input n_1729;
input n_5777;
input n_4225;
input n_300;
input n_747;
input n_2565;
input n_5495;
input n_1389;
input n_535;
input n_3583;
input n_3860;
input n_3851;
input n_5655;
input n_5064;
input n_5610;
input n_3015;
input n_2175;
input n_601;
input n_2182;
input n_4009;
input n_1848;
input n_5002;
input n_5759;
input n_1506;
input n_119;
input n_3473;
input n_1652;
input n_6035;
input n_957;
input n_1994;
input n_2566;
input n_387;
input n_744;
input n_971;
input n_2702;
input n_3241;
input n_2906;
input n_4342;
input n_4568;
input n_1205;
input n_6061;
input n_5559;
input n_1258;
input n_2438;
input n_2914;
input n_5786;
input n_3100;
input n_2180;
input n_2858;
input n_5377;
input n_3573;
input n_1016;
input n_4106;
input n_5737;
input n_1501;
input n_3604;
input n_4373;
input n_197;
input n_4711;
input n_3068;
input n_2685;
input n_1083;
input n_5768;
input n_3553;
input n_2275;
input n_2465;
input n_2568;
input n_2022;
input n_3811;
input n_910;
input n_3494;
input n_1721;
input n_1737;
input n_3486;
input n_4086;
input n_752;
input n_908;
input n_1028;
input n_2106;
input n_2265;
input n_5350;
input n_5470;
input n_2032;
input n_4812;
input n_4409;
input n_5872;
input n_5858;
input n_4629;
input n_4638;
input n_708;
input n_1973;
input n_3181;
input n_5700;
input n_1500;
input n_6037;
input n_3699;
input n_854;
input n_4913;
input n_2312;
input n_5874;
input n_904;
input n_709;
input n_1266;
input n_2242;
input n_3328;
input n_185;
input n_3868;
input n_1276;
input n_4266;
input n_2466;
input n_2530;
input n_5873;
input n_1085;
input n_2042;
input n_771;
input n_475;
input n_924;
input n_298;
input n_1582;
input n_492;
input n_5588;
input n_2318;
input n_3286;
input n_4012;
input n_1149;
input n_3170;
input n_265;
input n_3645;
input n_5075;
input n_3682;
input n_3304;
input n_2592;
input n_4968;
input n_3771;
input n_2666;
input n_1585;
input n_1799;
input n_2564;
input n_5085;
input n_5736;
input n_4259;
input n_2433;
input n_829;
input n_2035;
input n_3422;
input n_4572;
input n_859;
input n_3086;
input n_2033;
input n_406;
input n_4104;
input n_4845;
input n_1770;
input n_878;
input n_5120;
input n_130;
input n_3285;
input n_4208;
input n_981;
input n_5928;
input n_4089;
input n_5478;
input n_6016;
input n_1144;
input n_2071;
input n_3219;
input n_3702;
input n_2233;
input n_4779;
input n_481;
input n_3233;
input n_4599;
input n_997;
input n_4437;
input n_5222;
input n_3310;
input n_1306;
input n_3264;
input n_2010;
input n_1198;
input n_4061;
input n_2174;
input n_436;
input n_3881;
input n_4508;
input n_4727;
input n_4594;
input n_2426;
input n_2478;
input n_1133;
input n_95;
input n_4429;
input n_4642;
input n_4051;
input n_1051;
input n_4865;
input n_1039;
input n_2043;
input n_1480;
input n_6056;
input n_5832;
input n_3206;
input n_1305;
input n_2363;
input n_2578;
input n_4562;
input n_553;
input n_3383;
input n_4903;
input n_3709;
input n_3738;
input n_4186;
input n_5812;
input n_2540;
input n_973;
input n_5743;
input n_3610;
input n_4998;
input n_3330;
input n_2065;
input n_2879;
input n_967;
input n_4522;
input n_2001;
input n_4341;
input n_679;
input n_1629;
input n_5368;
input n_4263;
input n_225;
input n_1260;
input n_1819;
input n_309;
input n_3555;
input n_915;
input n_5971;
input n_812;
input n_1131;
input n_3155;
input n_1006;
input n_3110;
input n_1632;
input n_5933;
input n_257;
input n_1888;
input n_1311;
input n_4780;
input n_670;
input n_2697;
input n_3908;
input n_4973;
input n_3467;
input n_1887;
input n_1587;
input n_3916;
input n_3527;
input n_4803;
input n_2512;
input n_3950;
input n_6030;
input n_1242;
input n_2086;
input n_2927;
input n_4750;
input n_3039;
input n_1226;
input n_3740;
input n_5996;
input n_2166;
input n_2899;
input n_3186;
input n_640;
input n_1322;
input n_1958;
input n_315;
input n_5903;
input n_5986;
input n_1197;
input n_3065;
input n_2632;
input n_4984;
input n_2579;
input n_2105;
input n_135;
input n_1423;
input n_3387;
input n_364;
input n_5782;
input n_3420;
input n_5041;
input n_1915;
input n_4275;
input n_4283;
input n_4959;
input n_900;
input n_4426;
input n_2912;
input n_60;
input n_2659;
input n_4425;
input n_3409;
input n_4449;
input n_2116;
input n_2320;
input n_1013;
input n_1259;
input n_2183;
input n_3002;
input n_51;
input n_649;
input n_1612;
input n_4809;
input n_1199;
input n_3392;
input n_6050;
input n_625;
input n_226;
input n_68;
input n_212;
input n_3773;
input n_2003;
input n_1038;
input n_1581;
input n_3301;
input n_1357;
input n_4241;
input n_1853;
input n_798;
input n_2324;
input n_5563;
input n_245;
input n_1348;
input n_2977;
input n_1739;
input n_5840;
input n_1380;
input n_2847;
input n_2557;
input n_1009;
input n_62;
input n_2405;
input n_4050;
input n_1160;
input n_883;
input n_2647;
input n_1032;
input n_2336;
input n_1247;
input n_5717;
input n_6017;
input n_2521;
input n_1099;
input n_471;
input n_424;
input n_4578;
input n_2211;
input n_4777;
input n_5720;
input n_369;
input n_2672;
input n_4702;
input n_2299;
input n_4179;
input n_4895;
input n_5871;
input n_141;
input n_1285;
input n_1985;
input n_5898;
input n_1172;
input n_4026;
input n_71;
input n_4531;
input n_3282;
input n_1590;
input n_3626;
input n_1532;
input n_2313;
input n_5072;
input n_3106;
input n_1140;
input n_1670;
input n_2344;
input n_2365;
input n_4666;
input n_3031;
input n_4029;
input n_375;
input n_2447;
input n_4617;
input n_2340;
input n_4010;
input n_5896;
input n_1649;
input n_4555;
input n_5882;
input n_5940;
input n_5650;
input n_4969;
input n_6057;
input n_5105;
input n_1572;
input n_4308;
input n_5021;
input n_3463;
input n_428;
input n_5263;
input n_2510;
input n_1954;
input n_822;
input n_2791;
input n_4325;
input n_3251;
input n_4602;
input n_5044;
input n_5134;
input n_2212;
input n_3063;
input n_1163;
input n_2729;
input n_2582;
input n_1798;
input n_1550;
input n_491;
input n_3998;
input n_1591;
input n_3632;
input n_3122;
input n_5567;
input n_1344;
input n_2730;
input n_2495;
input n_371;
input n_5249;
input n_2090;
input n_2603;
input n_538;
input n_3829;
input n_4164;
input n_2173;
input n_5625;
input n_1471;
input n_4919;
input n_3737;
input n_5969;
input n_3655;
input n_493;
input n_3825;
input n_2880;
input n_3225;
input n_2108;
input n_5158;
input n_1211;
input n_5022;
input n_5670;
input n_1280;
input n_6041;
input n_3296;
input n_5276;
input n_58;
input n_1445;
input n_2551;
input n_1526;
input n_5047;
input n_196;
input n_2985;
input n_1978;
input n_574;
input n_3792;
input n_4202;
input n_1446;
input n_14;
input n_3938;
input n_4791;
input n_3507;
input n_5879;
input n_4403;
input n_5238;
input n_5855;
input n_3269;
input n_3531;
input n_473;
input n_1054;
input n_559;
input n_1956;
input n_4139;
input n_4549;
input n_1986;
input n_2397;
input n_3931;
input n_4349;
input n_5141;
input n_2113;
input n_1918;
input n_3603;
input n_5429;
input n_813;
input n_3822;
input n_4163;
input n_818;
input n_5535;
input n_645;
input n_3812;
input n_3910;
input n_2633;
input n_2207;
input n_4948;
input n_5268;
input n_2696;
input n_3482;
input n_4080;
input n_6002;
input n_2198;
input n_3319;
input n_541;
input n_2073;
input n_2273;
input n_3748;
input n_3272;
input n_4941;
input n_5506;
input n_5298;
input n_2;
input n_3396;
input n_4393;
input n_1162;
input n_4372;
input n_821;
input n_1068;
input n_982;
input n_5640;
input n_408;
input n_932;
input n_2831;
input n_4318;
input n_4158;
input n_3317;
input n_3978;
input n_5560;
input n_2123;
input n_1697;
input n_979;
input n_4074;
input n_3716;
input n_4795;
input n_5544;
input n_4918;
input n_3824;
input n_5067;
input n_5744;
input n_4013;
input n_5384;
input n_4544;
input n_3248;
input n_354;
input n_5841;
input n_134;
input n_2941;
input n_1278;
input n_547;
input n_5108;
input n_4032;
input n_1064;
input n_1396;
input n_634;
input n_2355;
input n_4147;
input n_136;
input n_4477;
input n_3168;
input n_2751;
input n_4337;
input n_4130;
input n_5941;
input n_2009;
input n_1793;
input n_3601;
input n_5611;
input n_3092;
input n_1289;
input n_3055;
input n_3966;
input n_2866;
input n_4742;
input n_1014;
input n_3734;
input n_1703;
input n_2580;
input n_882;
input n_3649;
input n_2821;
input n_1875;
input n_1865;
input n_5701;
input n_3746;
input n_6067;
input n_3384;
input n_1950;
input n_1563;
input n_3419;
input n_1297;
input n_1662;
input n_4478;
input n_1359;
input n_2818;
input n_5367;
input n_3794;
input n_674;
input n_3921;
input n_922;
input n_1335;
input n_1927;
input n_4838;
input n_5970;
input n_5202;
input n_702;
input n_4965;
input n_347;
input n_3346;
input n_1896;
input n_2965;
input n_3058;
input n_3861;
input n_675;
input n_1540;
input n_1977;
input n_3891;
input n_2193;
input n_4523;
input n_1655;
input n_242;
input n_6011;
input n_1886;
input n_4371;
input n_2994;
input n_5502;
input n_3428;
input n_3153;
input n_4552;
input n_3689;
input n_877;
input n_5850;
input n_4673;
input n_2519;
input n_728;
input n_3415;
input n_1063;
input n_4607;
input n_4041;
input n_2947;
input n_3918;
input n_5876;
input n_5521;
input n_1965;
input n_4837;
input n_2476;
input n_598;
input n_437;
input n_4169;
input n_697;
input n_3271;
input n_295;
input n_5088;
input n_4248;
input n_388;
input n_484;
input n_2976;
input n_2152;
input n_2652;
input n_1825;
input n_1757;
input n_170;
input n_1792;
input n_5856;
input n_1412;
input n_2497;
input n_3809;
input n_3139;
input n_4070;
input n_3545;
input n_3885;
input n_1369;
input n_881;
input n_3993;
input n_4685;
input n_63;
input n_4031;
input n_5837;
input n_148;
input n_4675;
input n_2663;
input n_5825;
input n_4018;
input n_5491;
input n_2987;
input n_694;
input n_2938;
input n_3780;
input n_5496;
input n_5802;
input n_297;
input n_3337;
input n_4002;
input n_3209;
input n_5178;
input n_1044;
input n_2165;
input n_5547;
input n_1391;
input n_131;
input n_2750;
input n_2775;
input n_1295;
input n_3477;
input n_2349;
input n_5596;
input n_6074;
input n_2684;
input n_5983;
input n_3146;
input n_1495;
input n_1438;
input n_3953;
input n_4588;
input n_1100;
input n_585;
input n_4653;
input n_4435;
input n_5604;
input n_1756;
input n_1128;
input n_5411;
input n_673;
input n_4019;
input n_1071;
input n_1968;
input n_4728;
input n_4999;
input n_4385;
input n_4922;
input n_865;
input n_3616;
input n_5815;
input n_4191;
input n_5695;
input n_6027;
input n_2870;
input n_59;
input n_2151;
input n_1839;
input n_2341;
input n_1765;
input n_3727;
input n_5235;
input n_2707;
input n_826;
input n_4350;
input n_3747;
input n_1714;
input n_104;
input n_718;
input n_5331;
input n_4330;
input n_542;
input n_5311;
input n_305;
input n_2089;
input n_3522;
input n_2747;
input n_3924;
input n_791;
input n_4621;
input n_4216;
input n_5797;
input n_510;
input n_4240;
input n_3491;
input n_5572;
input n_1488;
input n_704;
input n_2148;
input n_4162;
input n_5565;
input n_2339;
input n_2861;
input n_1999;
input n_2731;
input n_622;
input n_5520;
input n_147;
input n_3353;
input n_3018;
input n_3975;
input n_5800;
input n_5984;
input n_1838;
input n_2638;
input n_4785;
input n_4683;
input n_1766;
input n_1776;
input n_2002;
input n_2138;
input n_4021;
input n_2414;
input n_3014;
input n_1771;
input n_2316;
input n_4103;
input n_5060;
input n_3148;
input n_4022;
input n_4986;
input n_5888;
input n_5669;
input n_5772;
input n_145;
input n_2208;
input n_4775;
input n_5884;
input n_4864;
input n_5758;
input n_4674;
input n_4481;
input n_1304;
input n_294;
input n_3775;
input n_4669;
input n_2134;
input n_1176;
input n_425;
input n_5603;
input n_1431;
input n_3312;
input n_3835;
input n_4286;
input n_5763;
input n_2958;
input n_3731;
input n_1822;
input n_2936;
input n_3224;
input n_2489;
input n_6029;
input n_1087;
input n_657;
input n_5751;
input n_2771;
input n_3020;
input n_5264;
input n_4525;
input n_5924;
input n_1505;
input n_290;
input n_5712;
input n_3557;
input n_2610;
input n_3129;
input n_3620;
input n_478;
input n_107;
input n_3832;
input n_2520;
input n_4484;
input n_3693;
input n_446;
input n_4497;
input n_1568;
input n_2372;
input n_1490;
input n_526;
input n_2251;
input n_3674;
input n_2959;
input n_2501;
input n_3203;
input n_5694;
input n_4871;
input n_293;
input n_1070;
input n_2403;
input n_2837;
input n_4700;
input n_4883;
input n_1665;
input n_4306;
input n_154;
input n_4224;
input n_2127;
input n_3341;
input n_6005;
input n_4453;
input n_3559;
input n_5449;
input n_4005;
input n_3546;
input n_1358;
input n_3661;
input n_4564;
input n_5146;
input n_3056;
input n_745;
input n_2424;
input n_3201;
input n_3447;
input n_3971;
input n_5926;
input n_716;
input n_1475;
input n_1774;
input n_2354;
input n_3103;
input n_4573;
input n_5398;
input n_5860;
input n_2589;
input n_4535;
input n_755;
input n_527;
input n_2442;
input n_3627;
input n_3480;
input n_1368;
input n_1137;
input n_3612;
input n_4695;
input n_2545;
input n_3509;
input n_5919;
input n_4368;
input n_2966;
input n_2294;
input n_1942;
input n_1314;
input n_600;
input n_3196;
input n_864;
input n_5319;
input n_2504;
input n_2623;
input n_399;
input n_1440;
input n_5270;
input n_2063;
input n_1534;
input n_5005;
input n_6014;
input n_1339;
input n_2475;
input n_5181;
input n_403;
input n_723;
input n_3144;
input n_3244;
input n_596;
input n_1141;
input n_1268;
input n_3287;
input n_3322;
input n_1755;
input n_5043;
input n_2025;
input n_2357;
input n_5583;
input n_4654;
input n_3640;
input n_642;
input n_995;
input n_1159;
input n_3481;
input n_2250;
input n_3033;
input n_303;
input n_5775;
input n_2374;
input n_416;
input n_1681;
input n_6034;
input n_520;
input n_418;
input n_4597;
input n_113;
input n_3364;
input n_3226;
input n_2780;
input n_4020;
input n_5220;
input n_1618;
input n_4867;
input n_5061;
input n_1653;
input n_4063;
input n_4237;
input n_2601;
input n_5029;
input n_5127;
input n_6071;
input n_2920;
input n_773;
input n_920;
input n_99;
input n_1374;
input n_2648;
input n_3212;
input n_13;
input n_1169;
input n_1617;
input n_3370;
input n_3386;
input n_335;
input n_4721;
input n_463;
input n_3093;
input n_848;
input n_120;
input n_274;
input n_4247;
input n_3169;
input n_3205;
input n_1881;
input n_1267;
input n_1806;
input n_2023;
input n_2204;
input n_2720;
input n_496;
input n_4614;
input n_177;
input n_3360;
input n_2087;
input n_1636;
input n_3956;
input n_4001;
input n_1323;
input n_2627;
input n_4422;
input n_960;
input n_778;
input n_3004;
input n_3870;
input n_5177;
input n_5483;
input n_3625;
input n_1764;
input n_4632;
input n_1610;
input n_3084;
input n_5785;
input n_2343;
input n_793;
input n_5967;
input n_4546;
input n_4583;
input n_4963;
input n_3749;
input n_2942;
input n_4966;
input n_5780;
input n_4714;
input n_5037;
input n_2515;
input n_316;
input n_1551;
input n_4847;
input n_4054;
input n_2555;
input n_3586;
input n_3653;
input n_5966;
input n_2201;
input n_725;
input n_3349;
input n_4668;
input n_5213;
input n_4635;
input n_0;
input n_368;
input n_994;
input n_5735;
input n_2278;
input n_1020;
input n_1273;
input n_4214;
input n_3448;
input n_617;
input n_2924;
input n_1036;
input n_3595;
input n_1138;
input n_5752;
input n_1661;
input n_5360;
input n_421;
input n_3991;
input n_3516;
input n_3926;
input n_1095;
input n_1270;
input n_4405;
input n_610;
input n_4413;
input n_1852;
input n_4036;
input n_4759;
input n_2153;
input n_3670;
input n_2381;
input n_2052;
input n_179;
input n_4667;
input n_5081;
input n_517;
input n_4182;
input n_667;
input n_3230;
input n_1279;
input n_1115;
input n_1499;
input n_504;
input n_1409;
input n_5877;
input n_6018;
input n_5189;
input n_1503;
input n_2819;
input n_3041;
input n_4637;
input n_2423;
input n_603;
input n_1657;
input n_1126;
input n_2412;
input n_5869;
input n_2439;
input n_2404;
input n_1182;
input n_3635;
input n_5118;
input n_4155;
input n_4238;
input n_3011;
input n_2061;
input n_2757;
input n_4977;
input n_167;
input n_5632;
input n_5582;
input n_5425;
input n_5886;
input n_1216;
input n_2716;
input n_6032;
input n_2452;
input n_3650;
input n_5446;
input n_3010;
input n_3043;
input n_5224;
input n_4590;
input n_2543;
input n_5090;
input n_3137;
input n_2486;
input n_3560;
input n_3177;
input n_4929;
input n_5678;
input n_122;
input n_2220;
input n_2577;
input n_34;
input n_1262;
input n_3238;
input n_218;
input n_3529;
input n_70;
input n_4835;
input n_2232;
input n_4038;
input n_2790;
input n_4565;
input n_5414;
input n_4159;
input n_3784;
input n_5437;
input n_220;
input n_4586;
input n_1608;
input n_2373;
input n_1472;
input n_3628;
input n_5454;
input n_800;
input n_4734;
input n_1491;
input n_1840;
input n_4434;
input n_5307;
input n_2244;
input n_4290;
input n_2586;
input n_1684;
input n_2446;
input n_1346;
input n_1352;
input n_5407;
input n_2017;
input n_3029;
input n_3597;
input n_5913;
input n_1046;
input n_2560;
input n_2704;
input n_1145;
input n_1121;
input n_1102;
input n_1963;
input n_258;
input n_3790;
input n_2766;
input n_260;
input n_356;
input n_3318;
input n_4833;
input n_5062;
input n_5230;
input n_5944;
input n_152;
input n_4888;
input n_776;
input n_321;
input n_1823;
input n_2479;
input n_3350;
input n_6000;
input n_2782;
input n_3977;
input n_227;
input n_3588;
input n_4279;
input n_5008;
input n_1456;
input n_5004;
input n_5294;
input n_23;
input n_5974;
input n_2229;
input n_4133;
input n_4527;
input n_2288;
input n_6046;
input n_2099;
input n_5323;
input n_3388;
input n_4790;
input n_1946;
input n_4181;
input n_3184;
input n_5810;
input n_4561;
input n_4461;
input n_464;
input n_3245;
input n_3075;
input n_4007;
input n_4949;
input n_2642;
input n_4239;
input n_2383;
input n_5991;
input n_4184;
input n_1676;
input n_1830;
input n_2351;
input n_1319;
input n_5069;
input n_2986;
input n_5702;
input n_2536;
input n_3915;
input n_139;
input n_1633;
input n_3489;
input n_2835;
input n_5243;
input n_1416;
input n_5914;
input n_2820;
input n_2293;
input n_5250;
input n_3074;
input n_3102;
input n_5590;
input n_2026;
input n_1282;
input n_5260;
input n_550;
input n_3321;
input n_2567;
input n_5809;
input n_2322;
input n_275;
input n_2727;
input n_3377;
input n_560;
input n_4782;
input n_1321;
input n_2533;
input n_569;
input n_3530;
input n_2869;
input n_4378;
input n_5349;
input n_1235;
input n_2759;
input n_2361;
input n_1292;
input n_2266;
input n_4876;
input n_346;
input n_3;
input n_5813;
input n_790;
input n_5833;
input n_2611;
input n_2901;
input n_4358;
input n_5616;
input n_5805;
input n_2653;
input n_49;
input n_299;
input n_1248;
input n_902;
input n_2189;
input n_2246;
input n_4469;
input n_5169;
input n_431;
input n_5816;
input n_3156;
input n_672;
input n_1941;
input n_3483;
input n_5416;
input n_706;
input n_1794;
input n_1236;
input n_4493;
input n_4924;
input n_743;
input n_766;
input n_430;
input n_1746;
input n_3524;
input n_489;
input n_2885;
input n_636;
input n_110;
input n_3097;
input n_660;
input n_2062;
input n_4539;
input n_2975;
input n_4421;
input n_6072;
input n_2839;
input n_2856;
input n_4793;
input n_4498;
input n_2070;
input n_1607;
input n_1454;
input n_4953;
input n_2348;
input n_2944;
input n_3831;
input n_869;
input n_1154;
input n_646;
input n_528;
input n_391;
input n_1329;
input n_5167;
input n_5661;
input n_5830;
input n_5932;
input n_3589;
input n_262;
input n_897;
input n_846;
input n_2066;
input n_841;
input n_1476;
input n_3391;
input n_508;
input n_1800;
input n_1463;
input n_3458;
input n_4505;
input n_3190;
input n_1562;
input n_5558;
input n_1826;
input n_5687;
input n_57;
input n_5383;
input n_5126;
input n_1759;
input n_5051;
input n_52;
input n_5587;
input n_5236;
input n_853;
input n_875;
input n_5012;
input n_1678;
input n_661;
input n_3787;
input n_1256;
input n_3585;
input n_3565;
input n_4450;
input n_5954;
input n_7;
input n_5025;
input n_933;
input n_4173;
input n_3135;
input n_5651;
input n_4630;
input n_1217;
input n_5645;
input n_3990;
input n_310;
input n_1628;
input n_5766;
input n_2109;
input n_988;
input n_2796;
input n_2507;
input n_84;
input n_5878;
input n_5671;
input n_4534;
input n_1536;
input n_1204;
input n_1132;
input n_233;
input n_1327;
input n_955;
input n_246;
input n_2787;
input n_2969;
input n_2395;
input n_1554;
input n_4494;
input n_5412;
input n_769;
input n_2380;
input n_4786;
input n_1120;
input n_555;
input n_4579;
input n_669;
input n_2290;
input n_4811;
input n_2048;
input n_176;
input n_114;
input n_2005;
input n_4857;
input n_3432;
input n_2736;
input n_2883;
input n_1408;
input n_4282;
input n_1196;
input n_3493;
input n_863;
input n_3774;
input n_5733;
input n_2910;
input n_748;
input n_3268;
input n_1785;
input n_1147;
input n_1754;
input n_3057;
input n_3701;
input n_5148;
input n_2584;
input n_1812;
input n_866;
input n_2287;
input n_452;
input n_5791;
input n_5727;
input n_761;
input n_5946;
input n_5997;
input n_2492;
input n_3778;
input n_5328;
input n_5657;
input n_174;
input n_1173;
input n_4974;
input n_5975;
input n_4911;
input n_4436;
input n_5119;
input n_4569;
input n_1174;
input n_3334;
input n_5938;
input n_5602;
input n_647;
input n_5097;
input n_844;
input n_17;
input n_4985;
input n_2117;
input n_2234;
input n_3823;
input n_4384;
input n_2741;
input n_3114;
input n_888;
input n_2203;
input n_2255;
input n_3584;
input n_5246;
input n_236;
input n_4858;
input n_4678;
input n_2649;
input n_3556;
input n_3836;
input n_5579;
input n_414;
input n_1922;
input n_5750;
input n_4823;
input n_5831;
input n_4309;
input n_4363;
input n_1215;
input n_93;
input n_839;
input n_5107;
input n_3456;
input n_5095;
input n_779;
input n_1537;
input n_2205;
input n_4243;
input n_4025;
input n_3404;
input n_1122;
input n_5666;
input n_4059;
input n_1509;
input n_4121;
input n_3290;
input n_1109;
input n_4313;
input n_3309;
input n_3671;
input n_4142;
input n_2015;
input n_3982;
input n_2609;
input n_1161;
input n_5546;
input n_3796;
input n_232;
input n_3840;
input n_46;
input n_3461;
input n_3408;
input n_4246;
input n_3513;
input n_3690;
input n_1184;
input n_2483;
input n_4532;
input n_228;
input n_1525;
input n_3995;
input n_4076;
input n_2594;
input n_5994;
input n_4244;
input n_2147;
input n_592;
input n_2503;
input n_4049;
input n_1156;
input n_2600;
input n_984;
input n_5626;
input n_3508;
input n_132;
input n_868;
input n_4353;
input n_735;
input n_4787;
input n_5633;
input n_469;
input n_1218;
input n_5664;
input n_5921;
input n_3596;
input n_4537;
input n_4346;
input n_4351;
input n_357;
input n_2429;
input n_985;
input n_2440;
input n_6054;
input n_3521;
input n_802;
input n_561;
input n_980;
input n_2681;
input n_1651;
input n_2360;
input n_3764;
input n_4784;
input n_4075;
input n_116;
input n_5340;
input n_3947;
input n_1244;
input n_1685;
input n_3066;
input n_2844;
input n_2303;
input n_1619;
input n_2285;
input n_5280;
input n_4451;
input n_4332;
input n_810;
input n_1194;
input n_4538;
input n_4506;
input n_2742;
input n_3695;
input n_3976;
input n_3563;
input n_2367;
input n_201;
input n_3198;
input n_3495;
input n_1034;
input n_5925;
input n_2909;
input n_754;
input n_5369;
input n_975;
input n_43;
input n_5730;
input n_5576;
input n_3359;
input n_5272;
input n_467;
input n_3187;
input n_3218;
input n_582;
input n_861;
input n_857;
input n_2107;
input n_2040;
input n_2968;
input n_4201;
input n_4336;
input n_2221;
input n_588;
input n_5646;
input n_5624;
input n_4852;
input n_1010;
input n_4210;
input n_4981;
input n_1166;
input n_5440;
input n_2891;
input n_2709;
input n_534;
input n_1578;
input n_1861;
input n_3955;
input n_1557;
input n_2280;
input n_3945;
input n_730;
input n_5817;
input n_5214;
input n_203;
input n_1898;
input n_2443;
input n_4936;
input n_4205;
input n_2162;
input n_1868;
input n_207;
input n_2079;
input n_4763;
input n_3587;
input n_4278;
input n_5586;
input n_3433;
input n_4463;
input n_205;
input n_2185;
input n_6038;
input n_5861;
input n_1836;
input n_3833;
input n_2774;
input n_3162;
input n_1274;
input n_1486;
input n_3333;
input n_4129;
input n_5258;
input n_81;
input n_5032;
input n_1899;
input n_784;
input n_4804;
input n_5619;
input n_3965;
input n_5859;
input n_5380;
input n_4500;
input n_5065;
input n_862;
input n_5776;
input n_2098;
input n_3085;
input n_4433;
input n_5606;
input n_5644;
input n_2813;
input n_1935;
input n_5826;
input n_2027;
input n_2091;
input n_5920;
input n_2991;
input n_5030;
input n_4194;
input n_1449;
input n_4703;
input n_361;
input n_2419;
input n_5683;
input n_2677;
input n_3182;
input n_5756;
input n_3283;
input n_5527;
input n_1742;
input n_4030;

output n_20644;

wire n_18652;
wire n_18318;
wire n_16664;
wire n_19057;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_11111;
wire n_7933;
wire n_19613;
wire n_16335;
wire n_13125;
wire n_8186;
wire n_6725;
wire n_6126;
wire n_17647;
wire n_8899;
wire n_17634;
wire n_10053;
wire n_19785;
wire n_8534;
wire n_10020;
wire n_19715;
wire n_17991;
wire n_15665;
wire n_19382;
wire n_17735;
wire n_20091;
wire n_19161;
wire n_7161;
wire n_19232;
wire n_7868;
wire n_15764;
wire n_18903;
wire n_18105;
wire n_8561;
wire n_14998;
wire n_14944;
wire n_11954;
wire n_19220;
wire n_14341;
wire n_10392;
wire n_15074;
wire n_15253;
wire n_9626;
wire n_20377;
wire n_19097;
wire n_15898;
wire n_18013;
wire n_10719;
wire n_7389;
wire n_20151;
wire n_6913;
wire n_10015;
wire n_6948;
wire n_9362;
wire n_7516;
wire n_7401;
wire n_12767;
wire n_16095;
wire n_18502;
wire n_9658;
wire n_8426;
wire n_19755;
wire n_13681;
wire n_17209;
wire n_6243;
wire n_6585;
wire n_16553;
wire n_18122;
wire n_11543;
wire n_7651;
wire n_14662;
wire n_13247;
wire n_16286;
wire n_7956;
wire n_20321;
wire n_7369;
wire n_16549;
wire n_15421;
wire n_20011;
wire n_15964;
wire n_9100;
wire n_6784;
wire n_18310;
wire n_10868;
wire n_9067;
wire n_6323;
wire n_17847;
wire n_14431;
wire n_17478;
wire n_13515;
wire n_6110;
wire n_11684;
wire n_16324;
wire n_14410;
wire n_15800;
wire n_9400;
wire n_13139;
wire n_7774;
wire n_15600;
wire n_16267;
wire n_20471;
wire n_6951;
wire n_15899;
wire n_19991;
wire n_18317;
wire n_13729;
wire n_18709;
wire n_14813;
wire n_18002;
wire n_19810;
wire n_14628;
wire n_8421;
wire n_18863;
wire n_17854;
wire n_10114;
wire n_10357;
wire n_15762;
wire n_16351;
wire n_15883;
wire n_17706;
wire n_8389;
wire n_13711;
wire n_16721;
wire n_12742;
wire n_11768;
wire n_9267;
wire n_19401;
wire n_9652;
wire n_8849;
wire n_9059;
wire n_15332;
wire n_18445;
wire n_16254;
wire n_7564;
wire n_14989;
wire n_17564;
wire n_10204;
wire n_6383;
wire n_18669;
wire n_11637;
wire n_8151;
wire n_9038;
wire n_16004;
wire n_8748;
wire n_20487;
wire n_13984;
wire n_6794;
wire n_18608;
wire n_8718;
wire n_9935;
wire n_6990;
wire n_14288;
wire n_14824;
wire n_18699;
wire n_8223;
wire n_9135;
wire n_16800;
wire n_13771;
wire n_18644;
wire n_11295;
wire n_13960;
wire n_9070;
wire n_11708;
wire n_15629;
wire n_14401;
wire n_10827;
wire n_14922;
wire n_7569;
wire n_7823;
wire n_9477;
wire n_7062;
wire n_12158;
wire n_14769;
wire n_8577;
wire n_14961;
wire n_20559;
wire n_8594;
wire n_8428;
wire n_9829;
wire n_13341;
wire n_20345;
wire n_10685;
wire n_17139;
wire n_15185;
wire n_12083;
wire n_12014;
wire n_14803;
wire n_19270;
wire n_19816;
wire n_16035;
wire n_10607;
wire n_15490;
wire n_18033;
wire n_19569;
wire n_8164;
wire n_20485;
wire n_15100;
wire n_10368;
wire n_19137;
wire n_9088;
wire n_10183;
wire n_17161;
wire n_6952;
wire n_11464;
wire n_19421;
wire n_14878;
wire n_15046;
wire n_10383;
wire n_6776;
wire n_13550;
wire n_17601;
wire n_13348;
wire n_10724;
wire n_16398;
wire n_19396;
wire n_9988;
wire n_7009;
wire n_11553;
wire n_12795;
wire n_10876;
wire n_18780;
wire n_9137;
wire n_11180;
wire n_14043;
wire n_18820;
wire n_8995;
wire n_20006;
wire n_8711;
wire n_12505;
wire n_18602;
wire n_13721;
wire n_18430;
wire n_20018;
wire n_10820;
wire n_13514;
wire n_8306;
wire n_7488;
wire n_13194;
wire n_8887;
wire n_18677;
wire n_16183;
wire n_11866;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_15659;
wire n_9578;
wire n_13109;
wire n_7438;
wire n_20003;
wire n_20224;
wire n_16631;
wire n_14355;
wire n_7337;
wire n_9489;
wire n_14123;
wire n_10728;
wire n_6357;
wire n_6800;
wire n_18962;
wire n_10655;
wire n_9797;
wire n_8332;
wire n_9478;
wire n_11379;
wire n_16627;
wire n_19571;
wire n_19659;
wire n_19944;
wire n_10670;
wire n_11981;
wire n_19181;
wire n_9351;
wire n_14556;
wire n_6839;
wire n_9189;
wire n_18888;
wire n_16528;
wire n_14701;
wire n_7098;
wire n_16587;
wire n_19933;
wire n_18936;
wire n_20502;
wire n_8921;
wire n_20404;
wire n_9356;
wire n_15880;
wire n_16499;
wire n_18328;
wire n_9175;
wire n_6508;
wire n_12013;
wire n_11835;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_7782;
wire n_13385;
wire n_6636;
wire n_16339;
wire n_13992;
wire n_17429;
wire n_19103;
wire n_13790;
wire n_10624;
wire n_13304;
wire n_14633;
wire n_15699;
wire n_11900;
wire n_6538;
wire n_12883;
wire n_8983;
wire n_10422;
wire n_9818;
wire n_16503;
wire n_18974;
wire n_12367;
wire n_17360;
wire n_13526;
wire n_12563;
wire n_7243;
wire n_13321;
wire n_15042;
wire n_15519;
wire n_14722;
wire n_13427;
wire n_9909;
wire n_19607;
wire n_8620;
wire n_19204;
wire n_15264;
wire n_13270;
wire n_10052;
wire n_10109;
wire n_18151;
wire n_19582;
wire n_10448;
wire n_11196;
wire n_16239;
wire n_11963;
wire n_16334;
wire n_8424;
wire n_9571;
wire n_16003;
wire n_12655;
wire n_7941;
wire n_16096;
wire n_18628;
wire n_11483;
wire n_15067;
wire n_19591;
wire n_19345;
wire n_13356;
wire n_14912;
wire n_19177;
wire n_8907;
wire n_11080;
wire n_20447;
wire n_17557;
wire n_14079;
wire n_15168;
wire n_9894;
wire n_8324;
wire n_15411;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7913;
wire n_15144;
wire n_14224;
wire n_10380;
wire n_6449;
wire n_18687;
wire n_6461;
wire n_18273;
wire n_14682;
wire n_9033;
wire n_15031;
wire n_12933;
wire n_15718;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_17076;
wire n_13893;
wire n_11946;
wire n_9443;
wire n_9996;
wire n_14950;
wire n_20205;
wire n_7800;
wire n_13795;
wire n_17501;
wire n_14547;
wire n_15416;
wire n_20562;
wire n_17942;
wire n_18735;
wire n_9938;
wire n_7261;
wire n_9023;
wire n_14415;
wire n_11818;
wire n_16298;
wire n_18739;
wire n_6773;
wire n_13569;
wire n_7455;
wire n_18042;
wire n_19105;
wire n_9201;
wire n_6531;
wire n_10952;
wire n_13628;
wire n_18958;
wire n_9559;
wire n_11803;
wire n_15738;
wire n_16301;
wire n_8015;
wire n_18507;
wire n_19102;
wire n_15613;
wire n_14786;
wire n_9184;
wire n_13585;
wire n_18418;
wire n_18472;
wire n_8024;
wire n_12562;
wire n_18396;
wire n_16531;
wire n_20243;
wire n_11090;
wire n_19035;
wire n_13266;
wire n_13957;
wire n_9403;
wire n_9875;
wire n_11561;
wire n_19956;
wire n_8003;
wire n_8785;
wire n_17826;
wire n_8692;
wire n_6889;
wire n_16142;
wire n_9183;
wire n_14326;
wire n_16381;
wire n_10852;
wire n_9529;
wire n_11425;
wire n_6478;
wire n_6100;
wire n_6516;
wire n_17845;
wire n_6977;
wire n_16854;
wire n_17542;
wire n_7660;
wire n_6911;
wire n_6599;
wire n_6522;
wire n_17189;
wire n_9347;
wire n_18879;
wire n_16395;
wire n_13603;
wire n_6207;
wire n_6931;
wire n_7948;
wire n_9082;
wire n_6963;
wire n_8685;
wire n_16252;
wire n_19358;
wire n_10618;
wire n_9594;
wire n_7837;
wire n_20639;
wire n_19531;
wire n_9445;
wire n_7627;
wire n_9803;
wire n_20572;
wire n_16698;
wire n_17041;
wire n_7601;
wire n_6346;
wire n_19833;
wire n_15729;
wire n_17519;
wire n_14737;
wire n_11676;
wire n_12266;
wire n_16949;
wire n_12287;
wire n_19713;
wire n_13485;
wire n_12991;
wire n_11134;
wire n_13735;
wire n_8886;
wire n_7211;
wire n_10933;
wire n_8506;
wire n_6494;
wire n_16365;
wire n_11548;
wire n_13041;
wire n_17037;
wire n_13154;
wire n_7822;
wire n_6453;
wire n_9307;
wire n_10762;
wire n_11342;
wire n_7785;
wire n_11266;
wire n_19706;
wire n_12479;
wire n_8352;
wire n_18941;
wire n_10360;
wire n_9450;
wire n_16777;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_12537;
wire n_17183;
wire n_9693;
wire n_17582;
wire n_12921;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_13686;
wire n_13645;
wire n_16753;
wire n_12215;
wire n_18473;
wire n_9880;
wire n_12467;
wire n_6329;
wire n_11607;
wire n_11546;
wire n_15259;
wire n_16946;
wire n_15460;
wire n_7158;
wire n_20546;
wire n_13400;
wire n_9905;
wire n_18717;
wire n_13331;
wire n_9456;
wire n_20285;
wire n_7044;
wire n_9710;
wire n_8623;
wire n_11113;
wire n_18593;
wire n_17769;
wire n_19193;
wire n_13812;
wire n_14970;
wire n_7838;
wire n_16969;
wire n_12731;
wire n_7518;
wire n_6147;
wire n_9199;
wire n_13544;
wire n_7791;
wire n_18172;
wire n_12616;
wire n_18333;
wire n_14375;
wire n_12653;
wire n_7146;
wire n_18081;
wire n_16580;
wire n_18498;
wire n_9363;
wire n_12047;
wire n_12587;
wire n_10747;
wire n_13110;
wire n_16628;
wire n_9422;
wire n_18344;
wire n_12348;
wire n_16929;
wire n_16099;
wire n_15590;
wire n_10843;
wire n_7888;
wire n_11823;
wire n_6397;
wire n_16869;
wire n_10997;
wire n_19855;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_19640;
wire n_19157;
wire n_6331;
wire n_13498;
wire n_9341;
wire n_7848;
wire n_6939;
wire n_18289;
wire n_11408;
wire n_13183;
wire n_12519;
wire n_17184;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_13007;
wire n_10112;
wire n_7304;
wire n_20065;
wire n_7223;
wire n_7833;
wire n_14868;
wire n_9297;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_9808;
wire n_18534;
wire n_7445;
wire n_11086;
wire n_6529;
wire n_11710;
wire n_6290;
wire n_10253;
wire n_6455;
wire n_15277;
wire n_18435;
wire n_13804;
wire n_12455;
wire n_13099;
wire n_19524;
wire n_18516;
wire n_7695;
wire n_7179;
wire n_7122;
wire n_12157;
wire n_19676;
wire n_6203;
wire n_15806;
wire n_20604;
wire n_13064;
wire n_7630;
wire n_16246;
wire n_20013;
wire n_8643;
wire n_15660;
wire n_15357;
wire n_8565;
wire n_10821;
wire n_19784;
wire n_13648;
wire n_6892;
wire n_15722;
wire n_14181;
wire n_15278;
wire n_18054;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_14213;
wire n_17320;
wire n_17885;
wire n_7051;
wire n_8477;
wire n_19766;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_14842;
wire n_13115;
wire n_11759;
wire n_20195;
wire n_8230;
wire n_12549;
wire n_20388;
wire n_11601;
wire n_11971;
wire n_12314;
wire n_11116;
wire n_12604;
wire n_13305;
wire n_8876;
wire n_19017;
wire n_9359;
wire n_14189;
wire n_15761;
wire n_8060;
wire n_11124;
wire n_6392;
wire n_17470;
wire n_15301;
wire n_7351;
wire n_9352;
wire n_7608;
wire n_17053;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_13202;
wire n_15350;
wire n_13638;
wire n_17948;
wire n_14392;
wire n_19953;
wire n_19347;
wire n_7027;
wire n_7992;
wire n_6912;
wire n_10330;
wire n_8276;
wire n_11465;
wire n_8027;
wire n_17808;
wire n_11265;
wire n_11125;
wire n_17244;
wire n_20348;
wire n_7783;
wire n_13220;
wire n_10276;
wire n_8978;
wire n_10594;
wire n_8245;
wire n_15072;
wire n_12910;
wire n_18725;
wire n_18215;
wire n_8454;
wire n_8891;
wire n_11690;
wire n_18719;
wire n_19142;
wire n_16194;
wire n_11373;
wire n_6403;
wire n_7947;
wire n_16826;
wire n_20370;
wire n_6491;
wire n_19519;
wire n_16321;
wire n_14072;
wire n_17120;
wire n_11412;
wire n_13039;
wire n_13130;
wire n_10441;
wire n_19500;
wire n_17237;
wire n_15671;
wire n_9124;
wire n_6661;
wire n_13719;
wire n_8847;
wire n_14548;
wire n_19099;
wire n_10841;
wire n_16076;
wire n_12313;
wire n_18071;
wire n_20266;
wire n_14661;
wire n_8356;
wire n_6136;
wire n_16384;
wire n_16416;
wire n_15305;
wire n_15588;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_13062;
wire n_7857;
wire n_7481;
wire n_14130;
wire n_14930;
wire n_10576;
wire n_16596;
wire n_6668;
wire n_15548;
wire n_16714;
wire n_19168;
wire n_6859;
wire n_18752;
wire n_13752;
wire n_10237;
wire n_19484;
wire n_13596;
wire n_12889;
wire n_18092;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_9515;
wire n_6971;
wire n_17957;
wire n_9642;
wire n_20470;
wire n_14231;
wire n_12385;
wire n_13219;
wire n_17449;
wire n_6351;
wire n_9382;
wire n_16392;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_19207;
wire n_13295;
wire n_16906;
wire n_18194;
wire n_17693;
wire n_6829;
wire n_17981;
wire n_13160;
wire n_15249;
wire n_11071;
wire n_10072;
wire n_17337;
wire n_10708;
wire n_13818;
wire n_15024;
wire n_8803;
wire n_18478;
wire n_19898;
wire n_9706;
wire n_15174;
wire n_17904;
wire n_10387;
wire n_13764;
wire n_20258;
wire n_19408;
wire n_11224;
wire n_8790;
wire n_15569;
wire n_10219;
wire n_11924;
wire n_15193;
wire n_9591;
wire n_6137;
wire n_14833;
wire n_10364;
wire n_11422;
wire n_8338;
wire n_14480;
wire n_12489;
wire n_8491;
wire n_16610;
wire n_9283;
wire n_19299;
wire n_12030;
wire n_20330;
wire n_12565;
wire n_15236;
wire n_14098;
wire n_9468;
wire n_14482;
wire n_17174;
wire n_14223;
wire n_15962;
wire n_12415;
wire n_17332;
wire n_10559;
wire n_13173;
wire n_15355;
wire n_15945;
wire n_14848;
wire n_18548;
wire n_7154;
wire n_16232;
wire n_8304;
wire n_19644;
wire n_19012;
wire n_11418;
wire n_6655;
wire n_19694;
wire n_19187;
wire n_9958;
wire n_14544;
wire n_7320;
wire n_16122;
wire n_18852;
wire n_14604;
wire n_14735;
wire n_19572;
wire n_19688;
wire n_13101;
wire n_6786;
wire n_8315;
wire n_16446;
wire n_15885;
wire n_17528;
wire n_18964;
wire n_11040;
wire n_11754;
wire n_14916;
wire n_9756;
wire n_13748;
wire n_11672;
wire n_10353;
wire n_10847;
wire n_10451;
wire n_15801;
wire n_17778;
wire n_12240;
wire n_12003;
wire n_7496;
wire n_12165;
wire n_19894;
wire n_10866;
wire n_18127;
wire n_9940;
wire n_6200;
wire n_14600;
wire n_11763;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_18730;
wire n_8535;
wire n_10653;
wire n_11587;
wire n_6373;
wire n_12280;
wire n_13461;
wire n_20253;
wire n_12492;
wire n_19535;
wire n_16282;
wire n_17011;
wire n_13188;
wire n_17639;
wire n_7131;
wire n_20271;
wire n_20416;
wire n_9586;
wire n_8909;
wire n_18977;
wire n_16356;
wire n_11843;
wire n_14614;
wire n_11629;
wire n_15147;
wire n_9554;
wire n_18246;
wire n_17180;
wire n_6546;
wire n_15927;
wire n_7060;
wire n_19439;
wire n_13217;
wire n_16332;
wire n_20489;
wire n_14397;
wire n_17971;
wire n_10853;
wire n_13802;
wire n_18559;
wire n_7761;
wire n_20055;
wire n_10338;
wire n_12978;
wire n_15668;
wire n_15137;
wire n_8496;
wire n_12476;
wire n_8568;
wire n_8852;
wire n_18423;
wire n_12023;
wire n_20560;
wire n_17655;
wire n_8637;
wire n_6168;
wire n_16225;
wire n_16677;
wire n_13413;
wire n_6450;
wire n_15153;
wire n_13203;
wire n_19128;
wire n_14462;
wire n_8456;
wire n_7137;
wire n_14933;
wire n_9920;
wire n_12598;
wire n_9039;
wire n_11854;
wire n_8573;
wire n_19070;
wire n_18623;
wire n_17389;
wire n_7743;
wire n_13230;
wire n_6179;
wire n_19230;
wire n_9125;
wire n_20244;
wire n_9139;
wire n_20080;
wire n_17941;
wire n_12733;
wire n_13750;
wire n_8775;
wire n_14104;
wire n_20228;
wire n_18695;
wire n_14684;
wire n_12245;
wire n_15713;
wire n_18124;
wire n_14572;
wire n_9972;
wire n_6083;
wire n_12909;
wire n_6434;
wire n_9157;
wire n_16417;
wire n_17880;
wire n_9324;
wire n_8807;
wire n_6933;
wire n_8521;
wire n_6547;
wire n_9442;
wire n_20145;
wire n_19374;
wire n_6984;
wire n_18394;
wire n_17392;
wire n_10763;
wire n_9957;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_17586;
wire n_18757;
wire n_6507;
wire n_9313;
wire n_6687;
wire n_9173;
wire n_6690;
wire n_7412;
wire n_12144;
wire n_9160;
wire n_9974;
wire n_19365;
wire n_12129;
wire n_14753;
wire n_13658;
wire n_20222;
wire n_14671;
wire n_16454;
wire n_17977;
wire n_18441;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_14674;
wire n_19496;
wire n_6524;
wire n_12835;
wire n_10129;
wire n_16089;
wire n_7523;
wire n_8654;
wire n_14229;
wire n_15060;
wire n_11241;
wire n_15520;
wire n_14188;
wire n_11508;
wire n_7141;
wire n_16139;
wire n_6505;
wire n_12636;
wire n_11227;
wire n_20221;
wire n_11218;
wire n_10195;
wire n_13722;
wire n_7327;
wire n_12938;
wire n_13057;
wire n_8367;
wire n_7367;
wire n_16439;
wire n_14897;
wire n_19251;
wire n_12173;
wire n_6905;
wire n_17520;
wire n_15925;
wire n_18255;
wire n_19275;
wire n_7368;
wire n_8011;
wire n_10263;
wire n_15141;
wire n_12411;
wire n_10280;
wire n_20484;
wire n_18634;
wire n_8570;
wire n_6163;
wire n_7628;
wire n_9074;
wire n_9408;
wire n_6553;
wire n_19190;
wire n_12568;
wire n_16163;
wire n_13478;
wire n_18256;
wire n_12970;
wire n_8902;
wire n_14295;
wire n_7557;
wire n_20022;
wire n_7128;
wire n_14367;
wire n_13915;
wire n_7594;
wire n_15057;
wire n_19479;
wire n_16300;
wire n_19236;
wire n_18288;
wire n_10504;
wire n_7788;
wire n_13783;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_20618;
wire n_7586;
wire n_7767;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_16402;
wire n_13705;
wire n_17986;
wire n_17771;
wire n_9277;
wire n_9257;
wire n_17773;
wire n_17070;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_18515;
wire n_7744;
wire n_10595;
wire n_7748;
wire n_6827;
wire n_20167;
wire n_19958;
wire n_18914;
wire n_11073;
wire n_20308;
wire n_7485;
wire n_18867;
wire n_11974;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_14920;
wire n_8671;
wire n_19196;
wire n_15313;
wire n_9671;
wire n_14994;
wire n_10080;
wire n_16505;
wire n_12228;
wire n_10570;
wire n_16120;
wire n_20119;
wire n_12929;
wire n_16065;
wire n_15075;
wire n_12261;
wire n_18007;
wire n_12106;
wire n_12291;
wire n_14510;
wire n_12124;
wire n_11755;
wire n_9510;
wire n_18055;
wire n_13497;
wire n_15406;
wire n_19529;
wire n_14396;
wire n_11918;
wire n_11748;
wire n_12433;
wire n_8701;
wire n_16810;
wire n_6499;
wire n_19678;
wire n_18158;
wire n_12217;
wire n_15922;
wire n_12097;
wire n_8097;
wire n_13851;
wire n_9679;
wire n_8645;
wire n_13272;
wire n_18954;
wire n_16411;
wire n_19507;
wire n_16717;
wire n_8824;
wire n_11673;
wire n_7712;
wire n_6276;
wire n_10499;
wire n_8340;
wire n_11387;
wire n_19975;
wire n_11333;
wire n_18425;
wire n_8455;
wire n_7208;
wire n_13613;
wire n_12185;
wire n_9770;
wire n_8681;
wire n_7406;
wire n_11417;
wire n_16044;
wire n_18656;
wire n_9592;
wire n_17507;
wire n_9180;
wire n_10922;
wire n_19013;
wire n_10718;
wire n_13821;
wire n_19198;
wire n_13712;
wire n_9625;
wire n_15041;
wire n_15393;
wire n_14144;
wire n_6851;
wire n_6460;
wire n_19429;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_20583;
wire n_15595;
wire n_8255;
wire n_15081;
wire n_8461;
wire n_6368;
wire n_16474;
wire n_20184;
wire n_6583;
wire n_16940;
wire n_17419;
wire n_20295;
wire n_12520;
wire n_17134;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_8792;
wire n_12436;
wire n_16344;
wire n_12808;
wire n_18275;
wire n_13801;
wire n_19286;
wire n_19920;
wire n_8523;
wire n_12143;
wire n_13879;
wire n_18064;
wire n_20084;
wire n_11806;
wire n_19682;
wire n_11050;
wire n_17714;
wire n_11484;
wire n_19483;
wire n_19183;
wire n_10295;
wire n_20418;
wire n_10336;
wire n_7716;
wire n_17903;
wire n_20256;
wire n_8954;
wire n_12212;
wire n_20277;
wire n_7540;
wire n_13231;
wire n_12624;
wire n_8552;
wire n_17412;
wire n_7558;
wire n_8373;
wire n_13165;
wire n_12151;
wire n_17407;
wire n_15204;
wire n_18284;
wire n_20188;
wire n_9970;
wire n_11365;
wire n_18138;
wire n_17016;
wire n_16081;
wire n_15341;
wire n_15477;
wire n_6233;
wire n_6377;
wire n_12402;
wire n_17959;
wire n_18782;
wire n_19942;
wire n_10361;
wire n_7143;
wire n_10424;
wire n_8965;
wire n_18454;
wire n_13476;
wire n_18399;
wire n_12162;
wire n_17087;
wire n_7497;
wire n_11829;
wire n_11517;
wire n_7793;
wire n_16102;
wire n_16274;
wire n_6991;
wire n_10556;
wire n_13776;
wire n_7248;
wire n_7204;
wire n_15835;
wire n_12852;
wire n_10567;
wire n_7578;
wire n_13343;
wire n_7654;
wire n_17339;
wire n_10230;
wire n_12675;
wire n_13907;
wire n_12821;
wire n_14782;
wire n_18756;
wire n_7120;
wire n_8728;
wire n_6335;
wire n_12837;
wire n_8386;
wire n_14070;
wire n_14330;
wire n_13491;
wire n_18654;
wire n_15748;
wire n_17995;
wire n_14235;
wire n_6173;
wire n_14851;
wire n_18012;
wire n_10058;
wire n_16471;
wire n_20619;
wire n_19434;
wire n_7757;
wire n_17539;
wire n_6630;
wire n_8396;
wire n_16560;
wire n_6612;
wire n_6606;
wire n_13450;
wire n_19533;
wire n_14178;
wire n_20314;
wire n_12907;
wire n_15500;
wire n_14891;
wire n_17051;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_9028;
wire n_17217;
wire n_8020;
wire n_9374;
wire n_20386;
wire n_13634;
wire n_18027;
wire n_10413;
wire n_19268;
wire n_19948;
wire n_17786;
wire n_12708;
wire n_10369;
wire n_6821;
wire n_9983;
wire n_6688;
wire n_8580;
wire n_9993;
wire n_13622;
wire n_11207;
wire n_16951;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_14794;
wire n_17684;
wire n_9237;
wire n_13931;
wire n_14404;
wire n_6557;
wire n_18302;
wire n_6753;
wire n_18164;
wire n_17151;
wire n_7341;
wire n_12088;
wire n_15423;
wire n_14377;
wire n_6639;
wire n_12508;
wire n_12096;
wire n_8832;
wire n_20059;
wire n_19412;
wire n_19399;
wire n_11098;
wire n_15815;
wire n_20537;
wire n_7957;
wire n_10938;
wire n_6627;
wire n_17147;
wire n_18019;
wire n_10927;
wire n_8592;
wire n_11204;
wire n_6190;
wire n_16920;
wire n_12701;
wire n_20187;
wire n_10578;
wire n_16199;
wire n_19113;
wire n_6615;
wire n_17331;
wire n_7294;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_8622;
wire n_15367;
wire n_19095;
wire n_8104;
wire n_18511;
wire n_17428;
wire n_10746;
wire n_9188;
wire n_16407;
wire n_18009;
wire n_19002;
wire n_8779;
wire n_10697;
wire n_11714;
wire n_16179;
wire n_15070;
wire n_20040;
wire n_7250;
wire n_8762;
wire n_17503;
wire n_18365;
wire n_17358;
wire n_13419;
wire n_9207;
wire n_11860;
wire n_17057;
wire n_10926;
wire n_8897;
wire n_11503;
wire n_17104;
wire n_8376;
wire n_18271;
wire n_18998;
wire n_15640;
wire n_6271;
wire n_15683;
wire n_16202;
wire n_8599;
wire n_13460;
wire n_15451;
wire n_15233;
wire n_9637;
wire n_6716;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_13105;
wire n_14467;
wire n_20154;
wire n_14789;
wire n_13076;
wire n_15526;
wire n_12950;
wire n_8628;
wire n_19867;
wire n_15150;
wire n_13028;
wire n_8547;
wire n_7113;
wire n_20510;
wire n_10433;
wire n_9116;
wire n_14096;
wire n_11983;
wire n_10839;
wire n_11813;
wire n_14583;
wire n_14893;
wire n_20148;
wire n_20504;
wire n_8275;
wire n_6198;
wire n_18270;
wire n_6762;
wire n_19826;
wire n_9035;
wire n_16960;
wire n_14915;
wire n_17780;
wire n_17075;
wire n_9678;
wire n_8247;
wire n_6577;
wire n_12956;
wire n_17373;
wire n_14856;
wire n_15235;
wire n_20634;
wire n_9284;
wire n_20039;
wire n_15711;
wire n_7604;
wire n_9606;
wire n_17018;
wire n_13459;
wire n_14268;
wire n_10297;
wire n_12553;
wire n_19928;
wire n_14127;
wire n_8827;
wire n_19884;
wire n_17937;
wire n_9549;
wire n_14894;
wire n_12866;
wire n_17801;
wire n_6845;
wire n_9482;
wire n_8877;
wire n_9412;
wire n_15561;
wire n_6321;
wire n_6819;
wire n_10136;
wire n_15148;
wire n_16457;
wire n_19560;
wire n_11356;
wire n_20615;
wire n_15955;
wire n_8688;
wire n_20250;
wire n_10692;
wire n_14826;
wire n_16421;
wire n_15776;
wire n_11280;
wire n_14987;
wire n_8686;
wire n_12239;
wire n_17641;
wire n_19823;
wire n_8403;
wire n_11493;
wire n_17742;
wire n_8588;
wire n_15229;
wire n_11339;
wire n_15804;
wire n_15269;
wire n_20394;
wire n_10471;
wire n_14946;
wire n_18727;
wire n_15674;
wire n_17933;
wire n_8780;
wire n_17384;
wire n_7958;
wire n_18037;
wire n_11885;
wire n_15855;
wire n_10777;
wire n_16490;
wire n_7760;
wire n_13306;
wire n_9753;
wire n_8722;
wire n_16489;
wire n_19580;
wire n_8589;
wire n_20130;
wire n_7573;
wire n_6281;
wire n_7364;
wire n_13133;
wire n_8608;
wire n_12874;
wire n_10469;
wire n_11194;
wire n_11480;
wire n_18650;
wire n_9342;
wire n_18062;
wire n_9329;
wire n_19257;
wire n_17119;
wire n_9868;
wire n_7048;
wire n_16491;
wire n_8145;
wire n_8928;
wire n_17638;
wire n_7682;
wire n_18584;
wire n_20643;
wire n_6231;
wire n_12509;
wire n_14902;
wire n_6932;
wire n_13527;
wire n_7901;
wire n_7658;
wire n_10055;
wire n_10979;
wire n_19753;
wire n_19765;
wire n_6996;
wire n_15935;
wire n_17674;
wire n_10408;
wire n_16180;
wire n_8572;
wire n_17182;
wire n_6337;
wire n_18212;
wire n_8227;
wire n_12936;
wire n_18424;
wire n_19947;
wire n_10482;
wire n_7405;
wire n_14151;
wire n_20538;
wire n_8314;
wire n_9386;
wire n_15120;
wire n_11121;
wire n_11270;
wire n_6310;
wire n_11689;
wire n_10003;
wire n_15601;
wire n_15936;
wire n_20426;
wire n_10321;
wire n_9661;
wire n_20452;
wire n_14284;
wire n_13232;
wire n_13001;
wire n_17377;
wire n_9901;
wire n_17334;
wire n_8934;
wire n_13059;
wire n_6365;
wire n_8407;
wire n_8567;
wire n_15455;
wire n_11288;
wire n_12772;
wire n_11042;
wire n_10726;
wire n_16534;
wire n_19304;
wire n_14681;
wire n_11272;
wire n_14230;
wire n_8283;
wire n_14546;
wire n_20361;
wire n_9882;
wire n_16484;
wire n_10637;
wire n_9205;
wire n_17464;
wire n_7972;
wire n_13512;
wire n_7916;
wire n_9368;
wire n_13069;
wire n_12362;
wire n_19038;
wire n_6167;
wire n_13233;
wire n_18495;
wire n_8008;
wire n_18833;
wire n_13297;
wire n_20551;
wire n_6307;
wire n_7483;
wire n_14873;
wire n_19891;
wire n_9504;
wire n_14840;
wire n_16556;
wire n_6267;
wire n_17861;
wire n_6568;
wire n_19083;
wire n_7507;
wire n_7159;
wire n_18038;
wire n_16072;
wire n_14083;
wire n_10189;
wire n_8697;
wire n_6813;
wire n_6669;
wire n_8420;
wire n_8297;
wire n_10881;
wire n_13519;
wire n_16583;
wire n_20425;
wire n_15641;
wire n_16007;
wire n_17129;
wire n_19869;
wire n_8639;
wire n_16796;
wire n_16510;
wire n_15892;
wire n_14049;
wire n_7562;
wire n_12019;
wire n_8176;
wire n_14529;
wire n_17624;
wire n_16106;
wire n_10891;
wire n_9026;
wire n_10803;
wire n_13190;
wire n_6188;
wire n_11695;
wire n_17595;
wire n_8113;
wire n_18922;
wire n_15877;
wire n_11453;
wire n_19233;
wire n_17896;
wire n_19088;
wire n_16445;
wire n_6318;
wire n_16997;
wire n_14690;
wire n_19252;
wire n_17356;
wire n_10290;
wire n_19705;
wire n_11862;
wire n_14839;
wire n_15409;
wire n_16207;
wire n_9433;
wire n_18568;
wire n_11660;
wire n_14249;
wire n_14241;
wire n_6604;
wire n_16101;
wire n_6391;
wire n_10284;
wire n_14446;
wire n_14719;
wire n_15575;
wire n_19896;
wire n_8522;
wire n_12971;
wire n_7942;
wire n_16599;
wire n_6473;
wire n_18620;
wire n_15696;
wire n_14558;
wire n_19695;
wire n_11318;
wire n_17198;
wire n_7725;
wire n_16950;
wire n_20517;
wire n_20131;
wire n_8626;
wire n_19277;
wire n_19475;
wire n_15095;
wire n_11487;
wire n_8441;
wire n_7778;
wire n_8397;
wire n_17916;
wire n_8726;
wire n_17250;
wire n_6958;
wire n_15417;
wire n_16615;
wire n_14667;
wire n_6523;
wire n_14713;
wire n_7531;
wire n_18686;
wire n_13214;
wire n_8615;
wire n_15975;
wire n_11062;
wire n_14202;
wire n_15859;
wire n_11933;
wire n_14554;
wire n_9887;
wire n_20380;
wire n_13211;
wire n_8316;
wire n_19654;
wire n_8057;
wire n_14874;
wire n_20566;
wire n_18198;
wire n_18550;
wire n_16824;
wire n_15098;
wire n_16832;
wire n_13336;
wire n_16074;
wire n_19487;
wire n_18664;
wire n_13102;
wire n_12894;
wire n_10492;
wire n_15769;
wire n_9247;
wire n_17340;
wire n_8378;
wire n_10526;
wire n_8725;
wire n_9570;
wire n_12356;
wire n_19454;
wire n_11077;
wire n_9846;
wire n_13262;
wire n_10764;
wire n_18005;
wire n_18429;
wire n_9677;
wire n_6804;
wire n_6603;
wire n_17812;
wire n_7534;
wire n_8201;
wire n_16485;
wire n_9348;
wire n_14262;
wire n_8696;
wire n_6396;
wire n_20072;
wire n_12630;
wire n_6890;
wire n_12022;
wire n_19929;
wire n_10741;
wire n_6109;
wire n_14727;
wire n_12425;
wire n_14762;
wire n_13507;
wire n_10915;
wire n_18290;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_17133;
wire n_17729;
wire n_15410;
wire n_9707;
wire n_16002;
wire n_16258;
wire n_13594;
wire n_20096;
wire n_10680;
wire n_14228;
wire n_16131;
wire n_11473;
wire n_19856;
wire n_11726;
wire n_15944;
wire n_12574;
wire n_20407;
wire n_8833;
wire n_10142;
wire n_7828;
wire n_9918;
wire n_18643;
wire n_15932;
wire n_16345;
wire n_9390;
wire n_19997;
wire n_10069;
wire n_17325;
wire n_8541;
wire n_18233;
wire n_13678;
wire n_12458;
wire n_19291;
wire n_14582;
wire n_6897;
wire n_13523;
wire n_9619;
wire n_11171;
wire n_15117;
wire n_20621;
wire n_19868;
wire n_9187;
wire n_16621;
wire n_13819;
wire n_15777;
wire n_14424;
wire n_18398;
wire n_14523;
wire n_11063;
wire n_18846;
wire n_20435;
wire n_9989;
wire n_8319;
wire n_12853;
wire n_12942;
wire n_9259;
wire n_12397;
wire n_16555;
wire n_15336;
wire n_14161;
wire n_6573;
wire n_16760;
wire n_7634;
wire n_13290;
wire n_13500;
wire n_11440;
wire n_16844;
wire n_10483;
wire n_17758;
wire n_20158;
wire n_7285;
wire n_11337;
wire n_12005;
wire n_11243;
wire n_8929;
wire n_9360;
wire n_18610;
wire n_20610;
wire n_9824;
wire n_15089;
wire n_20088;
wire n_8233;
wire n_6130;
wire n_7273;
wire n_14750;
wire n_17939;
wire n_14074;
wire n_20325;
wire n_12800;
wire n_16574;
wire n_15145;
wire n_17516;
wire n_8187;
wire n_9399;
wire n_15838;
wire n_15297;
wire n_13979;
wire n_9740;
wire n_12947;
wire n_20297;
wire n_20327;
wire n_17178;
wire n_20576;
wire n_9764;
wire n_20349;
wire n_15160;
wire n_12666;
wire n_7597;
wire n_12354;
wire n_14297;
wire n_17388;
wire n_16368;
wire n_12631;
wire n_19154;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_18426;
wire n_18073;
wire n_19995;
wire n_6921;
wire n_14675;
wire n_18905;
wire n_9826;
wire n_11942;
wire n_15998;
wire n_19138;
wire n_6624;
wire n_6956;
wire n_12966;
wire n_15851;
wire n_15884;
wire n_7329;
wire n_14502;
wire n_14533;
wire n_17935;
wire n_10752;
wire n_18630;
wire n_10067;
wire n_18021;
wire n_19841;
wire n_10399;
wire n_12498;
wire n_11010;
wire n_9590;
wire n_16017;
wire n_11588;
wire n_16346;
wire n_13956;
wire n_6880;
wire n_7418;
wire n_19305;
wire n_12387;
wire n_19783;
wire n_9497;
wire n_13255;
wire n_15911;
wire n_9219;
wire n_17376;
wire n_8028;
wire n_8914;
wire n_15276;
wire n_8391;
wire n_16343;
wire n_13749;
wire n_15552;
wire n_17722;
wire n_19370;
wire n_16228;
wire n_12862;
wire n_13621;
wire n_8216;
wire n_16953;
wire n_9982;
wire n_7804;
wire n_18948;
wire n_12656;
wire n_8313;
wire n_14828;
wire n_7656;
wire n_19150;
wire n_19971;
wire n_8263;
wire n_6438;
wire n_11936;
wire n_19132;
wire n_10374;
wire n_7332;
wire n_10382;
wire n_18247;
wire n_8374;
wire n_13223;
wire n_13451;
wire n_13939;
wire n_18909;
wire n_13728;
wire n_7386;
wire n_17824;
wire n_11018;
wire n_10981;
wire n_16014;
wire n_13379;
wire n_13781;
wire n_19311;
wire n_17513;
wire n_10344;
wire n_14613;
wire n_19451;
wire n_11515;
wire n_17466;
wire n_15881;
wire n_7637;
wire n_16577;
wire n_10318;
wire n_18422;
wire n_18091;
wire n_12890;
wire n_20067;
wire n_13994;
wire n_17060;
wire n_11972;
wire n_13484;
wire n_17298;
wire n_8460;
wire n_20462;
wire n_17468;
wire n_14593;
wire n_16013;
wire n_7409;
wire n_19266;
wire n_10735;
wire n_17153;
wire n_13807;
wire n_9825;
wire n_7444;
wire n_16942;
wire n_17569;
wire n_18661;
wire n_14033;
wire n_10393;
wire n_15221;
wire n_16090;
wire n_18467;
wire n_9045;
wire n_12281;
wire n_9373;
wire n_14337;
wire n_11809;
wire n_17994;
wire n_9967;
wire n_13553;
wire n_20291;
wire n_7187;
wire n_19039;
wire n_17063;
wire n_19692;
wire n_9182;
wire n_9365;
wire n_18960;
wire n_10909;
wire n_6336;
wire n_10083;
wire n_18891;
wire n_9224;
wire n_10347;
wire n_6541;
wire n_12410;
wire n_16327;
wire n_19238;
wire n_14707;
wire n_16043;
wire n_19677;
wire n_14612;
wire n_12294;
wire n_7603;
wire n_10667;
wire n_17688;
wire n_18794;
wire n_7979;
wire n_13382;
wire n_11675;
wire n_20094;
wire n_15543;
wire n_15906;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_11083;
wire n_17418;
wire n_7866;
wire n_7205;
wire n_18283;
wire n_11728;
wire n_11698;
wire n_9556;
wire n_8590;
wire n_16682;
wire n_17038;
wire n_15798;
wire n_11326;
wire n_6421;
wire n_19743;
wire n_11870;
wire n_7407;
wire n_20193;
wire n_6328;
wire n_11283;
wire n_6236;
wire n_11834;
wire n_13361;
wire n_17286;
wire n_15061;
wire n_6144;
wire n_11506;
wire n_10135;
wire n_13161;
wire n_14010;
wire n_16413;
wire n_19796;
wire n_15030;
wire n_18205;
wire n_9152;
wire n_16451;
wire n_19965;
wire n_19590;
wire n_8364;
wire n_15228;
wire n_15832;
wire n_10720;
wire n_10535;
wire n_17629;
wire n_19349;
wire n_17536;
wire n_6708;
wire n_11236;
wire n_18793;
wire n_19987;
wire n_18529;
wire n_6242;
wire n_12379;
wire n_18222;
wire n_12932;
wire n_14078;
wire n_18985;
wire n_8548;
wire n_19793;
wire n_10672;
wire n_7645;
wire n_14222;
wire n_16990;
wire n_20155;
wire n_12114;
wire n_10308;
wire n_11608;
wire n_14430;
wire n_10623;
wire n_6285;
wire n_16545;
wire n_19339;
wire n_13709;
wire n_17713;
wire n_9454;
wire n_10586;
wire n_8742;
wire n_12626;
wire n_11967;
wire n_9253;
wire n_15084;
wire n_13559;
wire n_20332;
wire n_20596;
wire n_8874;
wire n_15071;
wire n_11996;
wire n_9566;
wire n_11338;
wire n_13426;
wire n_18826;
wire n_7666;
wire n_11250;
wire n_15328;
wire n_7963;
wire n_6398;
wire n_8329;
wire n_9503;
wire n_8270;
wire n_16051;
wire n_11738;
wire n_18196;
wire n_11522;
wire n_7737;
wire n_16569;
wire n_8614;
wire n_18459;
wire n_9568;
wire n_15621;
wire n_18411;
wire n_20170;
wire n_8816;
wire n_9119;
wire n_19337;
wire n_13529;
wire n_6224;
wire n_18293;
wire n_20455;
wire n_19616;
wire n_6614;
wire n_18395;
wire n_20379;
wire n_12554;
wire n_8035;
wire n_12722;
wire n_6735;
wire n_17445;
wire n_20581;
wire n_10491;
wire n_12037;
wire n_15371;
wire n_17572;
wire n_13453;
wire n_15080;
wire n_20178;
wire n_9943;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_7152;
wire n_9575;
wire n_10409;
wire n_11822;
wire n_10521;
wire n_9610;
wire n_16483;
wire n_14016;
wire n_12323;
wire n_15566;
wire n_20298;
wire n_10527;
wire n_7570;
wire n_7817;
wire n_11394;
wire n_9928;
wire n_11820;
wire n_13897;
wire n_14792;
wire n_16290;
wire n_14248;
wire n_8370;
wire n_13300;
wire n_16296;
wire n_20521;
wire n_7566;
wire n_11940;
wire n_9217;
wire n_12901;
wire n_10518;
wire n_20480;
wire n_7617;
wire n_15170;
wire n_16936;
wire n_19262;
wire n_9771;
wire n_15774;
wire n_7718;
wire n_13844;
wire n_19246;
wire n_7396;
wire n_18543;
wire n_18930;
wire n_7998;
wire n_12432;
wire n_7561;
wire n_18349;
wire n_6810;
wire n_17010;
wire n_17040;
wire n_16130;
wire n_12879;
wire n_13746;
wire n_12559;
wire n_13508;
wire n_14660;
wire n_9899;
wire n_19930;
wire n_13004;
wire n_13479;
wire n_8277;
wire n_18014;
wire n_14437;
wire n_13759;
wire n_10486;
wire n_16613;
wire n_8724;
wire n_15938;
wire n_17216;
wire n_15146;
wire n_9995;
wire n_9076;
wire n_12351;
wire n_16360;
wire n_19146;
wire n_19878;
wire n_13359;
wire n_10372;
wire n_14867;
wire n_8867;
wire n_9491;
wire n_12702;
wire n_17811;
wire n_15188;
wire n_12439;
wire n_19478;
wire n_11008;
wire n_6125;
wire n_7314;
wire n_14186;
wire n_7526;
wire n_17816;
wire n_14023;
wire n_19758;
wire n_17890;
wire n_10736;
wire n_19550;
wire n_11575;
wire n_7004;
wire n_14418;
wire n_8308;
wire n_18897;
wire n_8165;
wire n_14283;
wire n_8400;
wire n_18177;
wire n_10446;
wire n_7879;
wire n_16372;
wire n_15958;
wire n_18853;
wire n_7696;
wire n_11570;
wire n_16567;
wire n_12952;
wire n_19096;
wire n_14795;
wire n_19318;
wire n_19886;
wire n_16425;
wire n_16769;
wire n_8217;
wire n_10603;
wire n_6962;
wire n_12004;
wire n_12830;
wire n_8858;
wire n_7246;
wire n_10255;
wire n_20172;
wire n_20420;
wire n_11490;
wire n_8689;
wire n_10113;
wire n_15086;
wire n_6853;
wire n_10188;
wire n_10686;
wire n_9841;
wire n_19916;
wire n_8743;
wire n_7087;
wire n_8753;
wire n_6191;
wire n_16838;
wire n_10974;
wire n_11067;
wire n_8627;
wire n_20294;
wire n_13659;
wire n_12034;
wire n_16586;
wire n_16056;
wire n_13303;
wire n_6894;
wire n_13346;
wire n_13702;
wire n_9179;
wire n_15894;
wire n_8752;
wire n_18237;
wire n_18367;
wire n_10937;
wire n_12134;
wire n_12449;
wire n_16399;
wire n_6284;
wire n_10167;
wire n_12524;
wire n_18113;
wire n_6883;
wire n_12963;
wire n_10428;
wire n_16860;
wire n_17869;
wire n_20140;
wire n_19199;
wire n_18682;
wire n_12366;
wire n_14951;
wire n_11068;
wire n_11035;
wire n_19148;
wire n_12729;
wire n_13292;
wire n_12198;
wire n_9420;
wire n_16995;
wire n_14336;
wire n_7825;
wire n_10079;
wire n_7212;
wire n_19436;
wire n_6966;
wire n_15435;
wire n_8634;
wire n_9531;
wire n_12605;
wire n_20202;
wire n_6253;
wire n_12828;
wire n_10258;
wire n_14960;
wire n_8532;
wire n_19109;
wire n_12661;
wire n_10588;
wire n_8991;
wire n_8065;
wire n_11140;
wire n_17882;
wire n_17677;
wire n_8518;
wire n_19845;
wire n_18226;
wire n_13017;
wire n_16884;
wire n_15199;
wire n_18153;
wire n_9812;
wire n_15419;
wire n_7361;
wire n_9949;
wire n_20200;
wire n_14889;
wire n_7228;
wire n_9576;
wire n_6338;
wire n_15267;
wire n_19366;
wire n_6266;
wire n_14796;
wire n_19125;
wire n_11364;
wire n_12790;
wire n_8632;
wire n_19069;
wire n_17397;
wire n_7018;
wire n_19952;
wire n_7975;
wire n_10009;
wire n_9279;
wire n_11902;
wire n_16782;
wire n_11993;
wire n_10443;
wire n_17317;
wire n_12813;
wire n_13534;
wire n_10384;
wire n_7978;
wire n_10293;
wire n_17422;
wire n_20036;
wire n_12312;
wire n_10074;
wire n_13097;
wire n_17850;
wire n_15786;
wire n_9632;
wire n_20542;
wire n_12256;
wire n_11812;
wire n_9711;
wire n_9431;
wire n_14650;
wire n_18068;
wire n_14610;
wire n_11505;
wire n_7316;
wire n_17938;
wire n_18955;
wire n_7103;
wire n_14601;
wire n_11363;
wire n_15794;
wire n_20164;
wire n_17066;
wire n_14645;
wire n_11151;
wire n_15825;
wire n_10716;
wire n_10664;
wire n_19819;
wire n_20392;
wire n_11434;
wire n_6873;
wire n_8494;
wire n_20056;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_19536;
wire n_10749;
wire n_8788;
wire n_10992;
wire n_19380;
wire n_10560;
wire n_10160;
wire n_7404;
wire n_13171;
wire n_12857;
wire n_18615;
wire n_9854;
wire n_14854;
wire n_15266;
wire n_7271;
wire n_9713;
wire n_16501;
wire n_19264;
wire n_10300;
wire n_9588;
wire n_14218;
wire n_15107;
wire n_6842;
wire n_13876;
wire n_18935;
wire n_14487;
wire n_9127;
wire n_20019;
wire n_16767;
wire n_9869;
wire n_14449;
wire n_17094;
wire n_12885;
wire n_15539;
wire n_9715;
wire n_17112;
wire n_8618;
wire n_18916;
wire n_12108;
wire n_7535;
wire n_20469;
wire n_11531;
wire n_19450;
wire n_9407;
wire n_14476;
wire n_15244;
wire n_19574;
wire n_11824;
wire n_20201;
wire n_6957;
wire n_9361;
wire n_13976;
wire n_16578;
wire n_18949;
wire n_13579;
wire n_11566;
wire n_17452;
wire n_16650;
wire n_14639;
wire n_8990;
wire n_17067;
wire n_6444;
wire n_19170;
wire n_7944;
wire n_19235;
wire n_11374;
wire n_8647;
wire n_15857;
wire n_7016;
wire n_10782;
wire n_13557;
wire n_20162;
wire n_16709;
wire n_6379;
wire n_15589;
wire n_17491;
wire n_17757;
wire n_12754;
wire n_13583;
wire n_17333;
wire n_19043;
wire n_17749;
wire n_16658;
wire n_13455;
wire n_19136;
wire n_6232;
wire n_9132;
wire n_20339;
wire n_10861;
wire n_17035;
wire n_8879;
wire n_19639;
wire n_11203;
wire n_16157;
wire n_11159;
wire n_8052;
wire n_6362;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_9332;
wire n_17097;
wire n_16765;
wire n_11030;
wire n_6326;
wire n_10073;
wire n_14619;
wire n_7241;
wire n_10419;
wire n_7172;
wire n_15427;
wire n_17364;
wire n_10333;
wire n_12430;
wire n_18330;
wire n_7235;
wire n_6239;
wire n_13407;
wire n_13676;
wire n_18391;
wire n_16694;
wire n_12557;
wire n_13788;
wire n_6974;
wire n_16537;
wire n_18227;
wire n_18666;
wire n_8939;
wire n_13584;
wire n_15471;
wire n_12139;
wire n_9030;
wire n_7657;
wire n_20075;
wire n_19433;
wire n_9665;
wire n_7096;
wire n_13327;
wire n_19098;
wire n_11197;
wire n_7442;
wire n_10093;
wire n_20351;
wire n_15428;
wire n_15014;
wire n_6174;
wire n_7999;
wire n_10675;
wire n_6087;
wire n_16311;
wire n_10107;
wire n_15536;
wire n_20061;
wire n_13224;
wire n_11469;
wire n_14046;
wire n_7041;
wire n_10742;
wire n_10829;
wire n_19115;
wire n_12389;
wire n_9309;
wire n_19632;
wire n_10620;
wire n_13971;
wire n_16750;
wire n_7672;
wire n_7318;
wire n_20368;
wire n_19325;
wire n_12995;
wire n_18261;
wire n_14406;
wire n_13209;
wire n_11883;
wire n_14959;
wire n_19979;
wire n_15387;
wire n_11901;
wire n_6352;
wire n_15973;
wire n_8542;
wire n_19747;
wire n_10859;
wire n_18446;
wire n_8576;
wire n_14807;
wire n_8038;
wire n_11572;
wire n_14493;
wire n_18306;
wire n_13113;
wire n_13387;
wire n_8716;
wire n_19411;
wire n_16807;
wire n_18538;
wire n_17576;
wire n_18665;
wire n_15538;
wire n_11399;
wire n_17578;
wire n_8768;
wire n_10884;
wire n_15870;
wire n_12035;
wire n_13006;
wire n_12791;
wire n_7600;
wire n_14742;
wire n_6644;
wire n_17878;
wire n_19528;
wire n_12810;
wire n_16930;
wire n_13947;
wire n_11322;
wire n_17562;
wire n_12241;
wire n_9343;
wire n_15895;
wire n_16554;
wire n_17779;
wire n_7347;
wire n_11057;
wire n_10969;
wire n_14474;
wire n_7383;
wire n_6805;
wire n_8863;
wire n_18501;
wire n_7759;
wire n_11551;
wire n_18049;
wire n_7479;
wire n_10598;
wire n_8947;
wire n_15494;
wire n_10717;
wire n_11118;
wire n_18579;
wire n_20592;
wire n_12674;
wire n_17727;
wire n_17839;
wire n_8510;
wire n_11410;
wire n_12230;
wire n_19282;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_17122;
wire n_16778;
wire n_12220;
wire n_6868;
wire n_16133;
wire n_12283;
wire n_7174;
wire n_9421;
wire n_19055;
wire n_13383;
wire n_18787;
wire n_17079;
wire n_8021;
wire n_7803;
wire n_15124;
wire n_12595;
wire n_11429;
wire n_15802;
wire n_15163;
wire n_13983;
wire n_9416;
wire n_6225;
wire n_6218;
wire n_17489;
wire n_9929;
wire n_12920;
wire n_13317;
wire n_9953;
wire n_6648;
wire n_15578;
wire n_10955;
wire n_7927;
wire n_11011;
wire n_9998;
wire n_11795;
wire n_9850;
wire n_12141;
wire n_20553;
wire n_9346;
wire n_7920;
wire n_12774;
wire n_14687;
wire n_20283;
wire n_11904;
wire n_8480;
wire n_17399;
wire n_7025;
wire n_15886;
wire n_17022;
wire n_15856;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_14357;
wire n_13044;
wire n_13228;
wire n_13518;
wire n_19763;
wire n_14008;
wire n_17069;
wire n_12746;
wire n_16162;
wire n_10970;
wire n_16285;
wire n_14927;
wire n_13881;
wire n_17205;
wire n_13747;
wire n_12532;
wire n_10238;
wire n_8931;
wire n_8334;
wire n_11681;
wire n_10890;
wire n_11202;
wire n_19513;
wire n_10552;
wire n_15254;
wire n_6595;
wire n_8539;
wire n_10205;
wire n_16947;
wire n_15747;
wire n_13899;
wire n_6306;
wire n_19386;
wire n_16235;
wire n_11663;
wire n_11331;
wire n_19472;
wire n_9528;
wire n_14348;
wire n_7583;
wire n_12201;
wire n_19334;
wire n_14086;
wire n_12499;
wire n_19173;
wire n_12448;
wire n_10610;
wire n_11187;
wire n_12761;
wire n_16455;
wire n_15004;
wire n_16625;
wire n_16025;
wire n_14552;
wire n_7353;
wire n_9490;
wire n_19767;
wire n_14575;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_7571;
wire n_16249;
wire n_20605;
wire n_16435;
wire n_16723;
wire n_11446;
wire n_10910;
wire n_8242;
wire n_20132;
wire n_11540;
wire n_13248;
wire n_17296;
wire n_19237;
wire n_9819;
wire n_15338;
wire n_8184;
wire n_20254;
wire n_6525;
wire n_13119;
wire n_12642;
wire n_12484;
wire n_6128;
wire n_13549;
wire n_17361;
wire n_16080;
wire n_9992;
wire n_15180;
wire n_15692;
wire n_19976;
wire n_12669;
wire n_14296;
wire n_6702;
wire n_19490;
wire n_11179;
wire n_17074;
wire n_7749;
wire n_10078;
wire n_11321;
wire n_14313;
wire n_9500;
wire n_18496;
wire n_8705;
wire n_19107;
wire n_11779;
wire n_7508;
wire n_14211;
wire n_7574;
wire n_13516;
wire n_14273;
wire n_20063;
wire n_12462;
wire n_16462;
wire n_18648;
wire n_6169;
wire n_18775;
wire n_15230;
wire n_12735;
wire n_10709;
wire n_12646;
wire n_19849;
wire n_15875;
wire n_7352;
wire n_10244;
wire n_20128;
wire n_18512;
wire n_12999;
wire n_12682;
wire n_14802;
wire n_6848;
wire n_17415;
wire n_10043;
wire n_14834;
wire n_8159;
wire n_14346;
wire n_16955;
wire n_7439;
wire n_17653;
wire n_14506;
wire n_18822;
wire n_16018;
wire n_14615;
wire n_15222;
wire n_6850;
wire n_18991;
wire n_15285;
wire n_13294;
wire n_6098;
wire n_20446;
wire n_7112;
wire n_11307;
wire n_19021;
wire n_17860;
wire n_18274;
wire n_9545;
wire n_9603;
wire n_9629;
wire n_18003;
wire n_12719;
wire n_10342;
wire n_15361;
wire n_19037;
wire n_16244;
wire n_17862;
wire n_13438;
wire n_15850;
wire n_9930;
wire n_14371;
wire n_12925;
wire n_14988;
wire n_9659;
wire n_16293;
wire n_9897;
wire n_9241;
wire n_14590;
wire n_14603;
wire n_8185;
wire n_11466;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_9291;
wire n_11982;
wire n_11873;
wire n_15821;
wire n_10185;
wire n_11182;
wire n_20037;
wire n_16250;
wire n_15768;
wire n_8220;
wire n_18807;
wire n_14145;
wire n_11991;
wire n_12875;
wire n_15064;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_13918;
wire n_13775;
wire n_9851;
wire n_11799;
wire n_8009;
wire n_7852;
wire n_10983;
wire n_9987;
wire n_7984;
wire n_18307;
wire n_19860;
wire n_18110;
wire n_14973;
wire n_16751;
wire n_7220;
wire n_18015;
wire n_20300;
wire n_18242;
wire n_6550;
wire n_8841;
wire n_12196;
wire n_15136;
wire n_10354;
wire n_7465;
wire n_13177;
wire n_12724;
wire n_14958;
wire n_6672;
wire n_16744;
wire n_17876;
wire n_15992;
wire n_7738;
wire n_17406;
wire n_19079;
wire n_8395;
wire n_6634;
wire n_14758;
wire n_18392;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_16802;
wire n_17909;
wire n_18439;
wire n_19022;
wire n_13311;
wire n_19700;
wire n_20587;
wire n_16020;
wire n_11513;
wire n_7464;
wire n_8937;
wire n_7115;
wire n_12087;
wire n_13675;
wire n_15022;
wire n_18693;
wire n_6104;
wire n_10537;
wire n_6082;
wire n_18305;
wire n_10426;
wire n_9167;
wire n_12082;
wire n_9655;
wire n_20448;
wire n_11436;
wire n_11729;
wire n_19276;
wire n_12989;
wire n_8845;
wire n_15198;
wire n_17902;
wire n_13620;
wire n_7702;
wire n_6676;
wire n_9976;
wire n_8042;
wire n_17144;
wire n_12464;
wire n_9560;
wire n_18362;
wire n_18886;
wire n_20264;
wire n_15007;
wire n_15197;
wire n_8519;
wire n_18982;
wire n_9319;
wire n_12450;
wire n_19776;
wire n_14648;
wire n_11767;
wire n_10985;
wire n_9401;
wire n_11586;
wire n_12149;
wire n_12002;
wire n_12836;
wire n_19506;
wire n_17084;
wire n_13548;
wire n_15710;
wire n_11195;
wire n_16240;
wire n_9747;
wire n_14526;
wire n_13487;
wire n_17190;
wire n_17973;
wire n_8586;
wire n_9058;
wire n_18707;
wire n_18547;
wire n_16700;
wire n_10780;
wire n_17940;
wire n_8756;
wire n_13406;
wire n_16371;
wire n_7923;
wire n_14040;
wire n_8602;
wire n_14054;
wire n_13469;
wire n_10411;
wire n_13249;
wire n_12984;
wire n_18840;
wire n_13587;
wire n_10090;
wire n_14872;
wire n_8112;
wire n_18959;
wire n_11567;
wire n_19428;
wire n_9292;
wire n_18771;
wire n_12197;
wire n_17753;
wire n_19134;
wire n_11580;
wire n_13326;
wire n_6474;
wire n_13082;
wire n_6226;
wire n_18518;
wire n_10856;
wire n_12403;
wire n_9584;
wire n_13692;
wire n_8194;
wire n_8055;
wire n_8579;
wire n_10914;
wire n_8360;
wire n_20340;
wire n_6425;
wire n_6493;
wire n_14382;
wire n_13396;
wire n_10071;
wire n_8755;
wire n_11565;
wire n_14911;
wire n_15405;
wire n_15643;
wire n_15420;
wire n_13052;
wire n_11013;
wire n_20486;
wire n_16762;
wire n_16634;
wire n_10035;
wire n_18094;
wire n_20247;
wire n_18673;
wire n_18980;
wire n_14962;
wire n_17435;
wire n_8108;
wire n_17065;
wire n_12068;
wire n_17285;
wire n_10041;
wire n_15499;
wire n_14514;
wire n_17612;
wire n_8498;
wire n_14256;
wire n_17073;
wire n_16773;
wire n_19320;
wire n_14082;
wire n_20160;
wire n_7280;
wire n_7886;
wire n_15728;
wire n_6884;
wire n_7664;
wire n_18292;
wire n_7012;
wire n_17354;
wire n_12486;
wire n_7376;
wire n_15347;
wire n_10137;
wire n_12084;
wire n_16517;
wire n_20032;
wire n_11863;
wire n_17868;
wire n_17033;
wire n_17234;
wire n_16174;
wire n_18059;
wire n_19015;
wire n_10794;
wire n_14703;
wire n_13533;
wire n_6274;
wire n_8838;
wire n_12109;
wire n_16283;
wire n_9562;
wire n_7007;
wire n_16088;
wire n_12320;
wire n_19245;
wire n_9759;
wire n_6992;
wire n_15226;
wire n_19742;
wire n_19859;
wire n_10206;
wire n_17736;
wire n_6322;
wire n_15425;
wire n_16878;
wire n_7616;
wire n_18294;
wire n_9733;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_13011;
wire n_9981;
wire n_18514;
wire n_16513;
wire n_6378;
wire n_14495;
wire n_16879;
wire n_12269;
wire n_13486;
wire n_11463;
wire n_17541;
wire n_17394;
wire n_7587;
wire n_17496;
wire n_6930;
wire n_17472;
wire n_19121;
wire n_12802;
wire n_11569;
wire n_10064;
wire n_7197;
wire n_9676;
wire n_7393;
wire n_11332;
wire n_13629;
wire n_13207;
wire n_18025;
wire n_7358;
wire n_9950;
wire n_18088;
wire n_13589;
wire n_15730;
wire n_18089;
wire n_20591;
wire n_17967;
wire n_19731;
wire n_6929;
wire n_16706;
wire n_11309;
wire n_8045;
wire n_16032;
wire n_19740;
wire n_19741;
wire n_18910;
wire n_16959;
wire n_8209;
wire n_14477;
wire n_9213;
wire n_7291;
wire n_14522;
wire n_16971;
wire n_19998;
wire n_20526;
wire n_13561;
wire n_14720;
wire n_7437;
wire n_16873;
wire n_7618;
wire n_8575;
wire n_6620;
wire n_6597;
wire n_11105;
wire n_13698;
wire n_13894;
wire n_6586;
wire n_10474;
wire n_12689;
wire n_18939;
wire n_8789;
wire n_20616;
wire n_7953;
wire n_19775;
wire n_13540;
wire n_20642;
wire n_6428;
wire n_14642;
wire n_12042;
wire n_14827;
wire n_15481;
wire n_13465;
wire n_11130;
wire n_16149;
wire n_11664;
wire n_18705;
wire n_17430;
wire n_15388;
wire n_19242;
wire n_10652;
wire n_13733;
wire n_13098;
wire n_20029;
wire n_9388;
wire n_12654;
wire n_10869;
wire n_18708;
wire n_19112;
wire n_11783;
wire n_17837;
wire n_9911;
wire n_19603;
wire n_16317;
wire n_15187;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_17897;
wire n_10473;
wire n_15712;
wire n_16985;
wire n_19941;
wire n_8493;
wire n_10957;
wire n_13517;
wire n_20049;
wire n_11188;
wire n_10442;
wire n_13973;
wire n_7150;
wire n_8252;
wire n_11774;
wire n_7015;
wire n_13206;
wire n_7249;
wire n_15939;
wire n_7985;
wire n_13637;
wire n_16705;
wire n_18163;
wire n_8893;
wire n_6372;
wire n_15904;
wire n_12768;
wire n_18369;
wire n_16047;
wire n_10165;
wire n_8156;
wire n_19674;
wire n_14923;
wire n_13031;
wire n_19029;
wire n_19316;
wire n_17912;
wire n_13155;
wire n_13410;
wire n_19581;
wire n_7814;
wire n_8660;
wire n_13124;
wire n_11095;
wire n_19546;
wire n_8606;
wire n_9663;
wire n_16584;
wire n_18340;
wire n_9743;
wire n_19048;
wire n_11584;
wire n_14169;
wire n_7700;
wire n_10158;
wire n_10582;
wire n_16151;
wire n_10427;
wire n_11816;
wire n_18808;
wire n_16420;
wire n_11693;
wire n_15429;
wire n_9248;
wire n_6138;
wire n_10835;
wire n_11411;
wire n_19681;
wire n_13823;
wire n_11386;
wire n_20159;
wire n_11604;
wire n_13323;
wire n_12164;
wire n_16919;
wire n_12824;
wire n_13434;
wire n_16680;
wire n_16938;
wire n_10844;
wire n_17793;
wire n_14153;
wire n_6802;
wire n_10654;
wire n_6909;
wire n_13445;
wire n_17177;
wire n_19074;
wire n_18182;
wire n_15760;
wire n_16712;
wire n_14746;
wire n_11097;
wire n_14606;
wire n_12052;
wire n_9746;
wire n_8073;
wire n_8821;
wire n_19922;
wire n_9440;
wire n_17253;
wire n_20457;
wire n_20212;
wire n_20142;
wire n_17264;
wire n_15475;
wire n_8663;
wire n_20114;
wire n_10553;
wire n_19770;
wire n_8309;
wire n_8945;
wire n_15121;
wire n_10988;
wire n_19209;
wire n_20175;
wire n_6112;
wire n_16192;
wire n_18030;
wire n_9041;
wire n_8166;
wire n_10108;
wire n_13865;
wire n_10307;
wire n_8215;
wire n_19538;
wire n_17497;
wire n_6180;
wire n_8809;
wire n_12382;
wire n_6476;
wire n_14428;
wire n_6566;
wire n_11173;
wire n_16218;
wire n_6872;
wire n_13998;
wire n_17825;
wire n_10587;
wire n_8713;
wire n_15450;
wire n_7111;
wire n_20607;
wire n_7967;
wire n_13522;
wire n_15609;
wire n_16423;
wire n_9002;
wire n_14670;
wire n_9130;
wire n_19016;
wire n_7180;
wire n_13530;
wire n_8604;
wire n_16362;
wire n_7263;
wire n_14318;
wire n_17673;
wire n_17004;
wire n_11802;
wire n_20215;
wire n_8005;
wire n_13942;
wire n_18230;
wire n_12570;
wire n_11905;
wire n_19326;
wire n_20007;
wire n_10202;
wire n_15295;
wire n_9104;
wire n_17050;
wire n_17408;
wire n_15445;
wire n_8272;
wire n_13997;
wire n_14402;
wire n_14882;
wire n_11051;
wire n_11214;
wire n_7000;
wire n_7398;
wire n_18335;
wire n_14232;
wire n_12882;
wire n_19300;
wire n_18057;
wire n_12617;
wire n_8236;
wire n_13137;
wire n_19612;
wire n_15933;
wire n_17188;
wire n_6325;
wire n_9840;
wire n_10348;
wire n_12495;
wire n_9581;
wire n_8070;
wire n_18468;
wire n_16786;
wire n_7802;
wire n_17118;
wire n_15353;
wire n_19623;
wire n_6629;
wire n_15993;
wire n_17699;
wire n_19605;
wire n_8175;
wire n_8953;
wire n_17546;
wire n_17279;
wire n_19111;
wire n_10373;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_19511;
wire n_6914;
wire n_14121;
wire n_10381;
wire n_20163;
wire n_10947;
wire n_16984;
wire n_11261;
wire n_16012;
wire n_13929;
wire n_17739;
wire n_10767;
wire n_19684;
wire n_14646;
wire n_14095;
wire n_15069;
wire n_14520;
wire n_14780;
wire n_19828;
wire n_19966;
wire n_11447;
wire n_12652;
wire n_15507;
wire n_8142;
wire n_11627;
wire n_6404;
wire n_12209;
wire n_6674;
wire n_17883;
wire n_13606;
wire n_11659;
wire n_13501;
wire n_9106;
wire n_8869;
wire n_8381;
wire n_17149;
wire n_9520;
wire n_14931;
wire n_18774;
wire n_7770;
wire n_6968;
wire n_16268;
wire n_12371;
wire n_20027;
wire n_11497;
wire n_14900;
wire n_15846;
wire n_13454;
wire n_16662;
wire n_9042;
wire n_17329;
wire n_8987;
wire n_11805;
wire n_14935;
wire n_6282;
wire n_12770;
wire n_19551;
wire n_11635;
wire n_15434;
wire n_16530;
wire n_12951;
wire n_9453;
wire n_8118;
wire n_12393;
wire n_16442;
wire n_9718;
wire n_10281;
wire n_12831;
wire n_6431;
wire n_19620;
wire n_19839;
wire n_15767;
wire n_12427;
wire n_7533;
wire n_7221;
wire n_16026;
wire n_15159;
wire n_10656;
wire n_6575;
wire n_8246;
wire n_8952;
wire n_15154;
wire n_9680;
wire n_12172;
wire n_12923;
wire n_12147;
wire n_19624;
wire n_20204;
wire n_13227;
wire n_19683;
wire n_8848;
wire n_12825;
wire n_8259;
wire n_15182;
wire n_8349;
wire n_6836;
wire n_11998;
wire n_19900;
wire n_8776;
wire n_19391;
wire n_7753;
wire n_6771;
wire n_14732;
wire n_9947;
wire n_16659;
wire n_10138;
wire n_12117;
wire n_10375;
wire n_14535;
wire n_6795;
wire n_12960;
wire n_18972;
wire n_14094;
wire n_13033;
wire n_15703;
wire n_19353;
wire n_7648;
wire n_12131;
wire n_12851;
wire n_19854;
wire n_7452;
wire n_10320;
wire n_9269;
wire n_15518;
wire n_14217;
wire n_10903;
wire n_17596;
wire n_15574;
wire n_14062;
wire n_8453;
wire n_12740;
wire n_8949;
wire n_10831;
wire n_9131;
wire n_17580;
wire n_10517;
wire n_16889;
wire n_10323;
wire n_10842;
wire n_17620;
wire n_16465;
wire n_20519;
wire n_11146;
wire n_10883;
wire n_17785;
wire n_19249;
wire n_20493;
wire n_20106;
wire n_12278;
wire n_18918;
wire n_19018;
wire n_17672;
wire n_18036;
wire n_17414;
wire n_10123;
wire n_10651;
wire n_17483;
wire n_17689;
wire n_18975;
wire n_14785;
wire n_8500;
wire n_17857;
wire n_12804;
wire n_20458;
wire n_12116;
wire n_17438;
wire n_13755;
wire n_10468;
wire n_14126;
wire n_14105;
wire n_8285;
wire n_8483;
wire n_19145;
wire n_17696;
wire n_11370;
wire n_16731;
wire n_9020;
wire n_9895;
wire n_16452;
wire n_11585;
wire n_13140;
wire n_13962;
wire n_13753;
wire n_15365;
wire n_17141;
wire n_12560;
wire n_19295;
wire n_18171;
wire n_13610;
wire n_8851;
wire n_13332;
wire n_15293;
wire n_19405;
wire n_6097;
wire n_19214;
wire n_19779;
wire n_7093;
wire n_7840;
wire n_18797;
wire n_10024;
wire n_16386;
wire n_17101;
wire n_15695;
wire n_7080;
wire n_17984;
wire n_14156;
wire n_10711;
wire n_7624;
wire n_19915;
wire n_16185;
wire n_9186;
wire n_10818;
wire n_18851;
wire n_15178;
wire n_12222;
wire n_11951;
wire n_7003;
wire n_13604;
wire n_10788;
wire n_17163;
wire n_10563;
wire n_8810;
wire n_20427;
wire n_14518;
wire n_16310;
wire n_16477;
wire n_13397;
wire n_10178;
wire n_17731;
wire n_15360;
wire n_13132;
wire n_6609;
wire n_10115;
wire n_17157;
wire n_16927;
wire n_12793;
wire n_11778;
wire n_12406;
wire n_7484;
wire n_16639;
wire n_6414;
wire n_9470;
wire n_15516;
wire n_13792;
wire n_18229;
wire n_9405;
wire n_6264;
wire n_17426;
wire n_13480;
wire n_20233;
wire n_19583;
wire n_13571;
wire n_10984;
wire n_19723;
wire n_20249;
wire n_18742;
wire n_20255;
wire n_12001;
wire n_7883;
wire n_13715;
wire n_16675;
wire n_7458;
wire n_15186;
wire n_16935;
wire n_18576;
wire n_13810;
wire n_14403;
wire n_7435;
wire n_6997;
wire n_10509;
wire n_19292;
wire n_13473;
wire n_18267;
wire n_15963;
wire n_14353;
wire n_16589;
wire n_19213;
wire n_11742;
wire n_6891;
wire n_10031;
wire n_19163;
wire n_12235;
wire n_7663;
wire n_12204;
wire n_10898;
wire n_14386;
wire n_18784;
wire n_16472;
wire n_17830;
wire n_12098;
wire n_7917;
wire n_12579;
wire n_9203;
wire n_15073;
wire n_7532;
wire n_9613;
wire n_13982;
wire n_19921;
wire n_18703;
wire n_12611;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_7968;
wire n_6382;
wire n_18542;
wire n_9141;
wire n_15867;
wire n_11027;
wire n_11852;
wire n_8377;
wire n_9913;
wire n_19911;
wire n_9286;
wire n_19646;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_10819;
wire n_14521;
wire n_20024;
wire n_9704;
wire n_19468;
wire n_19025;
wire n_9046;
wire n_16576;
wire n_6339;
wire n_8814;
wire n_8530;
wire n_9193;
wire n_16882;
wire n_20353;
wire n_7711;
wire n_16181;
wire n_15948;
wire n_8984;
wire n_17123;
wire n_9290;
wire n_14580;
wire n_14028;
wire n_19131;
wire n_14772;
wire n_13827;
wire n_14542;
wire n_18632;
wire n_7230;
wire n_17552;
wire n_7989;
wire n_9778;
wire n_20511;
wire n_18986;
wire n_20109;
wire n_18280;
wire n_15003;
wire n_13200;
wire n_16783;
wire n_12848;
wire n_18963;
wire n_10315;
wire n_18321;
wire n_19104;
wire n_17187;
wire n_17031;
wire n_11455;
wire n_12368;
wire n_17240;
wire n_19795;
wire n_13193;
wire n_19798;
wire n_8462;
wire n_18953;
wire n_9380;
wire n_19881;
wire n_10062;
wire n_18235;
wire n_20115;
wire n_19476;
wire n_8429;
wire n_10514;
wire n_12785;
wire n_15312;
wire n_14155;
wire n_7620;
wire n_20034;
wire n_15818;
wire n_6079;
wire n_16481;
wire n_16430;
wire n_19313;
wire n_16715;
wire n_8492;
wire n_16565;
wire n_8135;
wire n_16620;
wire n_8445;
wire n_6427;
wire n_14978;
wire n_18353;
wire n_12639;
wire n_8895;
wire n_7811;
wire n_14649;
wire n_15940;
wire n_19955;
wire n_12175;
wire n_13536;
wire n_10512;
wire n_14714;
wire n_11384;
wire n_8273;
wire n_12353;
wire n_14129;
wire n_9761;
wire n_16962;
wire n_9087;
wire n_17832;
wire n_17316;
wire n_15333;
wire n_10434;
wire n_12869;
wire n_8312;
wire n_6781;
wire n_18585;
wire n_13830;
wire n_6133;
wire n_14184;
wire n_11889;
wire n_14183;
wire n_6127;
wire n_19172;
wire n_17751;
wire n_11362;
wire n_19256;
wire n_8078;
wire n_14200;
wire n_16558;
wire n_7926;
wire n_19118;
wire n_6598;
wire n_20359;
wire n_15568;
wire n_12502;
wire n_16859;
wire n_18800;
wire n_16703;
wire n_19666;
wire n_13191;
wire n_10131;
wire n_15464;
wire n_17741;
wire n_6867;
wire n_12600;
wire n_14536;
wire n_16338;
wire n_6139;
wire n_12133;
wire n_19939;
wire n_7965;
wire n_12919;
wire n_10273;
wire n_11416;
wire n_17485;
wire n_14321;
wire n_7474;
wire n_11169;
wire n_8650;
wire n_17843;
wire n_14654;
wire n_10503;
wire n_14664;
wire n_13215;
wire n_16834;
wire n_10465;
wire n_16073;
wire n_10590;
wire n_19890;
wire n_13782;
wire n_15476;
wire n_8526;
wire n_13751;
wire n_19988;
wire n_17150;
wire n_14019;
wire n_19140;
wire n_19418;
wire n_20385;
wire n_6759;
wire n_10786;
wire n_19806;
wire n_7028;
wire n_9890;
wire n_11492;
wire n_19653;
wire n_18904;
wire n_6535;
wire n_18801;
wire n_16644;
wire n_9817;
wire n_11160;
wire n_18899;
wire n_9782;
wire n_12319;
wire n_10805;
wire n_17214;
wire n_20356;
wire n_6643;
wire n_17982;
wire n_9471;
wire n_17012;
wire n_14896;
wire n_17440;
wire n_12930;
wire n_17181;
wire n_8351;
wire n_9069;
wire n_17371;
wire n_14030;
wire n_8603;
wire n_17274;
wire n_16660;
wire n_11343;
wire n_19143;
wire n_12575;
wire n_11451;
wire n_16853;
wire n_20050;
wire n_13384;
wire n_16048;
wire n_16262;
wire n_17127;
wire n_15422;
wire n_9003;
wire n_18874;
wire n_12418;
wire n_14837;
wire n_7312;
wire n_11269;
wire n_16849;
wire n_14103;
wire n_6689;
wire n_7632;
wire n_9172;
wire n_14653;
wire n_19464;
wire n_17275;
wire n_8980;
wire n_17573;
wire n_11311;
wire n_6698;
wire n_18553;
wire n_17345;
wire n_17770;
wire n_13242;
wire n_7707;
wire n_13282;
wire n_14436;
wire n_12113;
wire n_14599;
wire n_16087;
wire n_13352;
wire n_17648;
wire n_18116;
wire n_17853;
wire n_14812;
wire n_17871;
wire n_11293;
wire n_14728;
wire n_19184;
wire n_6363;
wire n_8619;
wire n_19224;
wire n_18217;
wire n_18812;
wire n_15122;
wire n_10134;
wire n_11603;
wire n_7277;
wire n_11271;
wire n_14778;
wire n_15714;
wire n_17270;
wire n_12015;
wire n_8146;
wire n_13690;
wire n_11562;
wire n_10194;
wire n_17085;
wire n_8910;
wire n_6408;
wire n_6150;
wire n_10077;
wire n_13619;
wire n_18508;
wire n_12031;
wire n_9278;
wire n_10889;
wire n_10010;
wire n_20472;
wire n_14996;
wire n_12126;
wire n_14543;
wire n_8550;
wire n_11094;
wire n_20046;
wire n_14747;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_9739;
wire n_14358;
wire n_9480;
wire n_17886;
wire n_12195;
wire n_19369;
wire n_6679;
wire n_19294;
wire n_13289;
wire n_13182;
wire n_16265;
wire n_16466;
wire n_13324;
wire n_9541;
wire n_11286;
wire n_15215;
wire n_18947;
wire n_17748;
wire n_16379;
wire n_16728;
wire n_7097;
wire n_8140;
wire n_15111;
wire n_18563;
wire n_8527;
wire n_12899;
wire n_18917;
wire n_17621;
wire n_19570;
wire n_7909;
wire n_6303;
wire n_8935;
wire n_15759;
wire n_20556;
wire n_10734;
wire n_16441;
wire n_15383;
wire n_11560;
wire n_10395;
wire n_14966;
wire n_11435;
wire n_15255;
wire n_6214;
wire n_9370;
wire n_13136;
wire n_6692;
wire n_14322;
wire n_12331;
wire n_8093;
wire n_13349;
wire n_9956;
wire n_17007;
wire n_6552;
wire n_17096;
wire n_8327;
wire n_13096;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_17005;
wire n_9487;
wire n_16791;
wire n_14608;
wire n_7306;
wire n_16153;
wire n_10118;
wire n_18791;
wire n_7470;
wire n_13800;
wire n_19593;
wire n_7693;
wire n_20568;
wire n_20498;
wire n_15662;
wire n_20077;
wire n_10002;
wire n_11242;
wire n_17974;
wire n_15923;
wire n_20052;
wire n_13694;
wire n_17494;
wire n_9660;
wire n_16233;
wire n_20371;
wire n_17344;
wire n_13093;
wire n_9328;
wire n_16511;
wire n_15274;
wire n_16410;
wire n_7653;
wire n_8354;
wire n_14276;
wire n_6959;
wire n_8353;
wire n_6388;
wire n_13185;
wire n_11053;
wire n_18635;
wire n_12159;
wire n_9434;
wire n_18450;
wire n_13855;
wire n_10902;
wire n_19596;
wire n_8348;
wire n_7032;
wire n_19086;
wire n_18806;
wire n_8211;
wire n_11304;
wire n_9681;
wire n_10485;
wire n_7475;
wire n_18448;
wire n_6435;
wire n_10536;
wire n_9079;
wire n_15544;
wire n_18738;
wire n_19564;
wire n_16145;
wire n_19424;
wire n_17512;
wire n_18931;
wire n_18988;
wire n_8653;
wire n_8920;
wire n_17521;
wire n_10950;
wire n_17477;
wire n_6682;
wire n_6823;
wire n_14550;
wire n_9089;
wire n_15346;
wire n_13477;
wire n_18200;
wire n_8942;
wire n_10978;
wire n_8222;
wire n_13808;
wire n_6822;
wire n_8553;
wire n_19608;
wire n_17068;
wire n_10187;
wire n_11014;
wire n_17508;
wire n_15033;
wire n_17789;
wire n_9564;
wire n_7391;
wire n_9230;
wire n_19301;
wire n_19297;
wire n_10768;
wire n_14067;
wire n_6389;
wire n_15903;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_13970;
wire n_19866;
wire n_15247;
wire n_16656;
wire n_10065;
wire n_8700;
wire n_13408;
wire n_17585;
wire n_15248;
wire n_13727;
wire n_17500;
wire n_13025;
wire n_10268;
wire n_18728;
wire n_14801;
wire n_12601;
wire n_15399;
wire n_17549;
wire n_13641;
wire n_20520;
wire n_19588;
wire n_19493;
wire n_8750;
wire n_17473;
wire n_17746;
wire n_10305;
wire n_16862;
wire n_12807;
wire n_15669;
wire n_18018;
wire n_7321;
wire n_8200;
wire n_16055;
wire n_19053;
wire n_18179;
wire n_18564;
wire n_12981;
wire n_19950;
wire n_6254;
wire n_13542;
wire n_8212;
wire n_20293;
wire n_20047;
wire n_9016;
wire n_14426;
wire n_15456;
wire n_11545;
wire n_8846;
wire n_12665;
wire n_19469;
wire n_16526;
wire n_16397;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_12592;
wire n_17467;
wire n_9029;
wire n_6837;
wire n_18860;
wire n_11043;
wire n_9414;
wire n_18539;
wire n_7023;
wire n_9615;
wire n_14205;
wire n_18532;
wire n_10779;
wire n_11061;
wire n_16495;
wire n_17922;
wire n_15742;
wire n_16686;
wire n_16347;
wire n_9811;
wire n_7899;
wire n_8631;
wire n_16385;
wire n_19141;
wire n_14723;
wire n_19205;
wire n_10520;
wire n_17437;
wire n_13531;
wire n_7797;
wire n_18641;
wire n_13880;
wire n_7687;
wire n_19992;
wire n_18251;
wire n_7582;
wire n_10541;
wire n_14587;
wire n_8959;
wire n_17326;
wire n_10614;
wire n_18834;
wire n_7809;
wire n_16877;
wire n_18169;
wire n_8425;
wire n_11257;
wire n_15176;
wire n_9910;
wire n_16790;
wire n_10217;
wire n_17255;
wire n_10743;
wire n_13424;
wire n_14658;
wire n_15066;
wire n_20481;
wire n_9651;
wire n_15474;
wire n_15316;
wire n_10270;
wire n_11115;
wire n_8001;
wire n_17417;
wire n_20260;
wire n_7529;
wire n_14233;
wire n_6881;
wire n_19269;
wire n_9544;
wire n_17324;
wire n_7520;
wire n_9831;
wire n_18245;
wire n_9697;
wire n_18878;
wire n_18414;
wire n_8362;
wire n_6300;
wire n_8256;
wire n_9310;
wire n_10132;
wire n_12091;
wire n_8704;
wire n_17589;
wire n_6132;
wire n_17493;
wire n_9294;
wire n_11747;
wire n_6395;
wire n_7054;
wire n_11858;
wire n_14027;
wire n_7433;
wire n_16316;
wire n_10075;
wire n_10423;
wire n_17762;
wire n_6171;
wire n_17291;
wire n_17895;
wire n_11895;
wire n_13458;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_10886;
wire n_18720;
wire n_13091;
wire n_13003;
wire n_6387;
wire n_10192;
wire n_9465;
wire n_13811;
wire n_19459;
wire n_14011;
wire n_10436;
wire n_19026;
wire n_12794;
wire n_15496;
wire n_6342;
wire n_17744;
wire n_15260;
wire n_15104;
wire n_12483;
wire n_20086;
wire n_16374;
wire n_18173;
wire n_17251;
wire n_18945;
wire n_17381;
wire n_9959;
wire n_15055;
wire n_11015;
wire n_18712;
wire n_9631;
wire n_14751;
wire n_6194;
wire n_20226;
wire n_18313;
wire n_12815;
wire n_15913;
wire n_10431;
wire n_9945;
wire n_17694;
wire n_16314;
wire n_15115;
wire n_8746;
wire n_20319;
wire n_11183;
wire n_10019;
wire n_8531;
wire n_12093;
wire n_19296;
wire n_11581;
wire n_6459;
wire n_8379;
wire n_13100;
wire n_16154;
wire n_12334;
wire n_18397;
wire n_9209;
wire n_7311;
wire n_18234;
wire n_7669;
wire n_8793;
wire n_12355;
wire n_19340;
wire n_15052;
wire n_9767;
wire n_9838;
wire n_9300;
wire n_11500;
wire n_12943;
wire n_20632;
wire n_17598;
wire n_17956;
wire n_20622;
wire n_11021;
wire n_8543;
wire n_16502;
wire n_7189;
wire n_13067;
wire n_6258;
wire n_16688;
wire n_10243;
wire n_9700;
wire n_18114;
wire n_18802;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_10596;
wire n_20512;
wire n_19671;
wire n_12140;
wire n_8063;
wire n_12599;
wire n_19419;
wire n_8032;
wire n_7427;
wire n_13250;
wire n_11190;
wire n_11794;
wire n_10519;
wire n_17630;
wire n_10163;
wire n_17409;
wire n_20186;
wire n_16544;
wire n_17529;
wire n_18979;
wire n_12330;
wire n_8129;
wire n_14819;
wire n_14890;
wire n_15871;
wire n_13906;
wire n_6760;
wire n_14265;
wire n_13664;
wire n_13566;
wire n_12591;
wire n_12466;
wire n_9509;
wire n_20089;
wire n_10874;
wire n_6825;
wire n_19558;
wire n_11831;
wire n_16213;
wire n_14399;
wire n_9628;
wire n_18940;
wire n_19348;
wire n_18279;
wire n_19655;
wire n_10250;
wire n_18658;
wire n_14063;
wire n_16657;
wire n_17584;
wire n_12041;
wire n_16734;
wire n_17783;
wire n_15157;
wire n_13074;
wire n_14716;
wire n_12876;
wire n_15286;
wire n_14698;
wire n_19152;
wire n_18633;
wire n_6468;
wire n_14323;
wire n_18565;
wire n_13071;
wire n_6857;
wire n_12536;
wire n_10795;
wire n_16333;
wire n_15116;
wire n_8049;
wire n_7762;
wire n_9467;
wire n_7186;
wire n_13739;
wire n_11157;
wire n_19809;
wire n_9097;
wire n_14364;
wire n_15472;
wire n_13234;
wire n_9314;
wire n_7017;
wire n_16718;
wire n_7830;
wire n_19217;
wire n_17380;
wire n_8084;
wire n_14113;
wire n_8289;
wire n_11178;
wire n_20492;
wire n_16428;
wire n_19010;
wire n_14938;
wire n_14784;
wire n_11432;
wire n_14179;
wire n_17755;
wire n_7191;
wire n_14979;
wire n_10412;
wire n_12650;
wire n_19935;
wire n_14324;
wire n_12859;
wire n_17763;
wire n_7961;
wire n_17176;
wire n_10617;
wire n_16524;
wire n_10544;
wire n_13030;
wire n_17819;
wire n_18475;
wire n_15094;
wire n_16880;
wire n_20287;
wire n_20153;
wire n_11952;
wire n_6422;
wire n_13896;
wire n_16473;
wire n_9873;
wire n_13299;
wire n_13042;
wire n_15658;
wire n_10095;
wire n_15873;
wire n_8268;
wire n_6160;
wire n_19749;
wire n_7066;
wire n_18128;
wire n_7789;
wire n_6192;
wire n_10056;
wire n_16597;
wire n_17627;
wire n_18815;
wire n_20296;
wire n_11919;
wire n_11414;
wire n_17705;
wire n_17728;
wire n_19457;
wire n_17618;
wire n_7344;
wire n_9888;
wire n_10037;
wire n_18029;
wire n_6707;
wire n_12744;
wire n_19601;
wire n_11136;
wire n_19790;
wire n_19527;
wire n_19672;
wire n_6787;
wire n_11620;
wire n_15480;
wire n_10179;
wire n_14038;
wire n_18726;
wire n_11215;
wire n_11890;
wire n_9366;
wire n_14253;
wire n_7915;
wire n_9077;
wire n_8406;
wire n_15919;
wire n_16652;
wire n_12443;
wire n_6463;
wire n_11683;
wire n_20135;
wire n_8554;
wire n_7538;
wire n_12934;
wire n_19547;
wire n_18981;
wire n_6799;
wire n_19368;
wire n_6487;
wire n_8818;
wire n_16648;
wire n_16724;
wire n_10466;
wire n_11953;
wire n_6563;
wire n_20415;
wire n_7554;
wire n_19005;
wire n_18881;
wire n_15926;
wire n_20210;
wire n_16943;
wire n_11089;
wire n_6341;
wire n_13422;
wire n_7421;
wire n_10166;
wire n_7489;
wire n_14702;
wire n_13179;
wire n_15844;
wire n_11839;
wire n_18039;
wire n_19874;
wire n_13834;
wire n_18277;
wire n_8341;
wire n_11193;
wire n_17800;
wire n_17613;
wire n_7188;
wire n_11217;
wire n_15651;
wire n_17759;
wire n_20014;
wire n_6923;
wire n_9287;
wire n_7991;
wire n_10877;
wire n_16737;
wire n_14686;
wire n_12214;
wire n_16259;
wire n_8926;
wire n_10766;
wire n_10086;
wire n_13924;
wire n_9608;
wire n_19539;
wire n_20313;
wire n_20251;
wire n_8817;
wire n_8190;
wire n_11488;
wire n_13671;
wire n_18571;
wire n_14876;
wire n_6987;
wire n_18265;
wire n_11037;
wire n_16925;
wire n_18740;
wire n_14319;
wire n_16763;
wire n_17462;
wire n_15287;
wire n_7671;
wire n_13150;
wire n_15103;
wire n_12541;
wire n_8649;
wire n_19757;
wire n_14818;
wire n_19508;
wire n_20422;
wire n_8303;
wire n_6153;
wire n_16512;
wire n_13809;
wire n_8059;
wire n_18364;
wire n_11665;
wire n_6579;
wire n_13590;
wire n_16747;
wire n_11138;
wire n_11731;
wire n_16257;
wire n_16200;
wire n_16023;
wire n_16041;
wire n_6789;
wire n_12100;
wire n_15327;
wire n_17718;
wire n_13471;
wire n_17615;
wire n_19063;
wire n_8862;
wire n_16161;
wire n_10580;
wire n_17287;
wire n_6164;
wire n_13261;
wire n_9675;
wire n_7786;
wire n_16923;
wire n_11454;
wire n_7609;
wire n_8900;
wire n_12523;
wire n_6934;
wire n_6737;
wire n_18388;
wire n_8478;
wire n_16988;
wire n_6695;
wire n_12395;
wire n_17475;
wire n_17363;
wire n_8497;
wire n_10770;
wire n_6410;
wire n_17873;
wire n_15592;
wire n_16064;
wire n_18524;
wire n_15319;
wire n_14452;
wire n_17894;
wire n_13464;
wire n_12670;
wire n_16817;
wire n_18336;
wire n_7667;
wire n_10203;
wire n_10980;
wire n_9174;
wire n_17835;
wire n_17459;
wire n_10082;
wire n_7182;
wire n_7365;
wire n_10467;
wire n_9849;
wire n_17476;
wire n_9856;
wire n_18449;
wire n_17591;
wire n_18672;
wire n_18848;
wire n_11668;
wire n_7885;
wire n_15684;
wire n_16720;
wire n_9349;
wire n_17423;
wire n_11091;
wire n_10940;
wire n_16463;
wire n_15976;
wire n_18100;
wire n_17723;
wire n_8839;
wire n_12891;
wire n_11615;
wire n_11059;
wire n_16403;
wire n_14616;
wire n_16799;
wire n_17965;
wire n_7745;
wire n_12941;
wire n_20219;
wire n_14258;
wire n_12200;
wire n_14024;
wire n_17212;
wire n_8684;
wire n_13682;
wire n_6249;
wire n_11060;
wire n_18943;
wire n_11461;
wire n_10714;
wire n_6969;
wire n_7459;
wire n_6161;
wire n_8206;
wire n_18070;
wire n_18338;
wire n_19908;
wire n_6607;
wire n_9335;
wire n_9452;
wire n_11427;
wire n_19293;
wire n_12673;
wire n_14694;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_19818;
wire n_19208;
wire n_9427;
wire n_17817;
wire n_6294;
wire n_9611;
wire n_18371;
wire n_9021;
wire n_16269;
wire n_9250;
wire n_11212;
wire n_13145;
wire n_9550;
wire n_16591;
wire n_11263;
wire n_10641;
wire n_18805;
wire n_16566;
wire n_13195;
wire n_8694;
wire n_13965;
wire n_11994;
wire n_13358;
wire n_18759;
wire n_16693;
wire n_14519;
wire n_6123;
wire n_11000;
wire n_16125;
wire n_20430;
wire n_19403;
wire n_8191;
wire n_10325;
wire n_16354;
wire n_10298;
wire n_6922;
wire n_16701;
wire n_7698;
wire n_12854;
wire n_16427;
wire n_16336;
wire n_8431;
wire n_19631;
wire n_16248;
wire n_10400;
wire n_19081;
wire n_9177;
wire n_9060;
wire n_11947;
wire n_14496;
wire n_9096;
wire n_13952;
wire n_11697;
wire n_16963;
wire n_18074;
wire n_7891;
wire n_14413;
wire n_8517;
wire n_10901;
wire n_11034;
wire n_10549;
wire n_12115;
wire n_11499;
wire n_10825;
wire n_17292;
wire n_18023;
wire n_14777;
wire n_14057;
wire n_17788;
wire n_16406;
wire n_12558;
wire n_11984;
wire n_11948;
wire n_7477;
wire n_17028;
wire n_15654;
wire n_17289;
wire n_11402;
wire n_11401;
wire n_17828;
wire n_19679;
wire n_17820;
wire n_10581;
wire n_14949;
wire n_17487;
wire n_18372;
wire n_12086;
wire n_16952;
wire n_16449;
wire n_11589;
wire n_11246;
wire n_18266;
wire n_16606;
wire n_14460;
wire n_13216;
wire n_12849;
wire n_11312;
wire n_13786;
wire n_9344;
wire n_19719;
wire n_10865;
wire n_7378;
wire n_10738;
wire n_9798;
wire n_15491;
wire n_14925;
wire n_11612;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_13414;
wire n_7498;
wire n_11916;
wire n_7501;
wire n_10421;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_12764;
wire n_15325;
wire n_18987;
wire n_20268;
wire n_19091;
wire n_14238;
wire n_16918;
wire n_12409;
wire n_11625;
wire n_17054;
wire n_20053;
wire n_6592;
wire n_9712;
wire n_8585;
wire n_6626;
wire n_19877;
wire n_14042;
wire n_9220;
wire n_17312;
wire n_12763;
wire n_18460;
wire n_17272;
wire n_20599;
wire n_16394;
wire n_18869;
wire n_20136;
wire n_15310;
wire n_17989;
wire n_8698;
wire n_12584;
wire n_14435;
wire n_10376;
wire n_15510;
wire n_7515;
wire n_17567;
wire n_9994;
wire n_14226;
wire n_7309;
wire n_15811;
wire n_8559;
wire n_20123;
wire n_17670;
wire n_15618;
wire n_10224;
wire n_15849;
wire n_18758;
wire n_20545;
wire n_19951;
wire n_9391;
wire n_16105;
wire n_8514;
wire n_9134;
wire n_14159;
wire n_14515;
wire n_12268;
wire n_18990;
wire n_12077;
wire n_15321;
wire n_14757;
wire n_12534;
wire n_6846;
wire n_13271;
wire n_11481;
wire n_10175;
wire n_15812;
wire n_16292;
wire n_18458;
wire n_6886;
wire n_17019;
wire n_8405;
wire n_15223;
wire n_11350;
wire n_11925;
wire n_16033;
wire n_8672;
wire n_6446;
wire n_9430;
wire n_19279;
wire n_7218;
wire n_11407;
wire n_19548;
wire n_12710;
wire n_19331;
wire n_8440;
wire n_7005;
wire n_9776;
wire n_16736;
wire n_6777;
wire n_18156;
wire n_11987;
wire n_18208;
wire n_19206;
wire n_8475;
wire n_8029;
wire n_18845;
wire n_18527;
wire n_13089;
wire n_15459;
wire n_15192;
wire n_18360;
wire n_16836;
wire n_13167;
wire n_20602;
wire n_12329;
wire n_15013;
wire n_6953;
wire n_16710;
wire n_14945;
wire n_18660;
wire n_18348;
wire n_19658;
wire n_18487;
wire n_9834;
wire n_16353;
wire n_12318;
wire n_13278;
wire n_13597;
wire n_7089;
wire n_18232;
wire n_20317;
wire n_6332;
wire n_20206;
wire n_7403;
wire n_7338;
wire n_7129;
wire n_13938;
wire n_13251;
wire n_8566;
wire n_7343;
wire n_12766;
wire n_18913;
wire n_8317;
wire n_12229;
wire n_6116;
wire n_7492;
wire n_13319;
wire n_9071;
wire n_10415;
wire n_7694;
wire n_11711;
wire n_18637;
wire n_15666;
wire n_20509;
wire n_11931;
wire n_8109;
wire n_18971;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_7987;
wire n_9133;
wire n_16054;
wire n_12664;
wire n_14942;
wire n_7434;
wire n_9009;
wire n_6155;
wire n_20449;
wire n_7269;
wire n_9777;
wire n_15359;
wire n_9063;
wire n_7787;
wire n_15035;
wire n_18500;
wire n_19085;
wire n_18536;
wire n_6261;
wire n_19893;
wire n_10096;
wire n_13617;
wire n_10025;
wire n_18779;
wire n_6299;
wire n_20573;
wire n_11753;
wire n_7425;
wire n_19061;
wire n_11150;
wire n_18199;
wire n_16111;
wire n_6316;
wire n_6292;
wire n_9726;
wire n_13884;
wire n_17125;
wire n_7719;
wire n_6220;
wire n_12783;
wire n_17671;
wire n_14195;
wire n_18363;
wire n_20479;
wire n_7938;
wire n_7935;
wire n_8458;
wire n_6772;
wire n_16902;
wire n_16646;
wire n_14300;
wire n_6077;
wire n_11512;
wire n_17090;
wire n_14678;
wire n_13599;
wire n_17282;
wire n_15008;
wire n_13647;
wire n_13683;
wire n_19094;
wire n_10147;
wire n_17921;
wire n_17197;
wire n_18503;
wire n_20474;
wire n_9298;
wire n_18058;
wire n_16939;
wire n_14497;
wire n_14280;
wire n_13724;
wire n_9301;
wire n_12054;
wire n_15827;
wire n_8099;
wire n_17256;
wire n_11595;
wire n_17806;
wire n_13768;
wire n_16707;
wire n_8578;
wire n_7222;
wire n_13838;
wire n_10046;
wire n_10397;
wire n_19379;
wire n_10936;
wire n_12442;
wire n_8611;
wire n_8819;
wire n_17927;
wire n_15123;
wire n_9835;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_7875;
wire n_13153;
wire n_7643;
wire n_13441;
wire n_16082;
wire n_10207;
wire n_13857;
wire n_18872;
wire n_10401;
wire n_19352;
wire n_7242;
wire n_17737;
wire n_19240;
wire n_13816;
wire n_18355;
wire n_17215;
wire n_19737;
wire n_14736;
wire n_10139;
wire n_13246;
wire n_14061;
wire n_12986;
wire n_11381;
wire n_16378;
wire n_16109;
wire n_7224;
wire n_12441;
wire n_15789;
wire n_16611;
wire n_16172;
wire n_7746;
wire n_18108;
wire n_16277;
wire n_16598;
wire n_17588;
wire n_12516;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_6653;
wire n_16806;
wire n_15512;
wire n_18836;
wire n_12377;
wire n_18486;
wire n_9965;
wire n_13650;
wire n_16789;
wire n_15636;
wire n_15946;
wire n_6501;
wire n_18063;
wire n_9990;
wire n_10005;
wire n_12905;
wire n_11426;
wire n_15311;
wire n_8505;
wire n_19827;
wire n_17667;
wire n_7884;
wire n_11258;
wire n_19879;
wire n_15498;
wire n_20477;
wire n_7417;
wire n_18097;
wire n_12513;
wire n_13395;
wire n_20016;
wire n_7388;
wire n_11657;
wire n_8717;
wire n_9064;
wire n_17420;
wire n_14135;
wire n_8571;
wire n_16482;
wire n_12514;
wire n_10048;
wire n_16809;
wire n_14194;
wire n_13825;
wire n_19945;
wire n_18942;
wire n_8243;
wire n_6347;
wire n_9593;
wire n_20630;
wire n_13398;
wire n_8449;
wire n_17605;
wire n_13204;
wire n_14331;
wire n_18994;
wire n_9406;
wire n_8967;
wire n_9322;
wire n_15017;
wire n_8031;
wire n_15591;
wire n_12188;
wire n_16609;
wire n_9232;
wire n_15167;
wire n_12299;
wire n_16739;
wire n_15706;
wire n_11327;
wire n_15900;
wire n_12000;
wire n_17281;
wire n_19004;
wire n_14182;
wire n_10279;
wire n_15853;
wire n_14352;
wire n_13889;
wire n_17864;
wire n_7081;
wire n_13015;
wire n_20112;
wire n_7319;
wire n_15831;
wire n_7644;
wire n_11176;
wire n_9883;
wire n_11135;
wire n_11275;
wire n_18850;
wire n_12700;
wire n_12904;
wire n_14623;
wire n_7910;
wire n_9034;
wire n_7084;
wire n_14073;
wire n_8074;
wire n_13639;
wire n_15989;
wire n_8860;
wire n_15514;
wire n_9266;
wire n_16210;
wire n_10027;
wire n_12784;
wire n_18639;
wire n_12877;
wire n_14677;
wire n_14261;
wire n_18020;
wire n_10616;
wire n_8587;
wire n_16016;
wire n_15550;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_9078;
wire n_16297;
wire n_16896;
wire n_13198;
wire n_15914;
wire n_13741;
wire n_12610;
wire n_14416;
wire n_11251;
wire n_12293;
wire n_6470;
wire n_11598;
wire n_8368;
wire n_15691;
wire n_17560;
wire n_8322;
wire n_16127;
wire n_6187;
wire n_8300;
wire n_9378;
wire n_12206;
wire n_18112;
wire n_17488;
wire n_17427;
wire n_11400;
wire n_19532;
wire n_19870;
wire n_6693;
wire n_15848;
wire n_11563;
wire n_12444;
wire n_18586;
wire n_16409;
wire n_14513;
wire n_12778;
wire n_12485;
wire n_15995;
wire n_14602;
wire n_11468;
wire n_16150;
wire n_9683;
wire n_17403;
wire n_15132;
wire n_11878;
wire n_15843;
wire n_16666;
wire n_15749;
wire n_7449;
wire n_15638;
wire n_16547;
wire n_14289;
wire n_16479;
wire n_10751;
wire n_16967;
wire n_10240;
wire n_10691;
wire n_9561;
wire n_19351;
wire n_16104;
wire n_20445;
wire n_9773;
wire n_9745;
wire n_15413;
wire n_10216;
wire n_15628;
wire n_17733;
wire n_10150;
wire n_12581;
wire n_17395;
wire n_6652;
wire n_10971;
wire n_20116;
wire n_18506;
wire n_7674;
wire n_14516;
wire n_18484;
wire n_12305;
wire n_12170;
wire n_9630;
wire n_13927;
wire n_13313;
wire n_15308;
wire n_17025;
wire n_9255;
wire n_10231;
wire n_8310;
wire n_16500;
wire n_9758;
wire n_15175;
wire n_8936;
wire n_7126;
wire n_18413;
wire n_15206;
wire n_9691;
wire n_12997;
wire n_14005;
wire n_14293;
wire n_14334;
wire n_7690;
wire n_15245;
wire n_15225;
wire n_11223;
wire n_13562;
wire n_14537;
wire n_6950;
wire n_10038;
wire n_17794;
wire n_15614;
wire n_20234;
wire n_18101;
wire n_19087;
wire n_11221;
wire n_15772;
wire n_14245;
wire n_20322;
wire n_17659;
wire n_11448;
wire n_17321;
wire n_18272;
wire n_8328;
wire n_15502;
wire n_15076;
wire n_12576;
wire n_7258;
wire n_10579;
wire n_13345;
wire n_8336;
wire n_20376;
wire n_17492;
wire n_19324;
wire n_20008;
wire n_11445;
wire n_13151;
wire n_11552;
wire n_15102;
wire n_14733;
wire n_14317;
wire n_19807;
wire n_16220;
wire n_9852;
wire n_11623;
wire n_18599;
wire n_14131;
wire n_8041;
wire n_10676;
wire n_10540;
wire n_10299;
wire n_17931;
wire n_16993;
wire n_12845;
wire n_11645;
wire n_10200;
wire n_13164;
wire n_13662;
wire n_16275;
wire n_17062;
wire n_13340;
wire n_17887;
wire n_17192;
wire n_9939;
wire n_7766;
wire n_19397;
wire n_12797;
wire n_20561;
wire n_6758;
wire n_19709;
wire n_9481;
wire n_7955;
wire n_17081;
wire n_12012;
wire n_7287;
wire n_10076;
wire n_6464;
wire n_18675;
wire n_20508;
wire n_11554;
wire n_9635;
wire n_19619;
wire n_14308;
wire n_8181;
wire n_8254;
wire n_13452;
wire n_8071;
wire n_20606;
wire n_17480;
wire n_11628;
wire n_20218;
wire n_11549;
wire n_20177;
wire n_17162;
wire n_12286;
wire n_9001;
wire n_19517;
wire n_16107;
wire n_14545;
wire n_18031;
wire n_8013;
wire n_19670;
wire n_16683;
wire n_17804;
wire n_12347;
wire n_19346;
wire n_17424;
wire n_20262;
wire n_19394;
wire n_17818;
wire n_20378;
wire n_12698;
wire n_6540;
wire n_16086;
wire n_17383;
wire n_11871;
wire n_16857;
wire n_15326;
wire n_17555;
wire n_18957;
wire n_7722;
wire n_20329;
wire n_9240;
wire n_8293;
wire n_14726;
wire n_14180;
wire n_18697;
wire n_10548;
wire n_12957;
wire n_11616;
wire n_8791;
wire n_8288;
wire n_12786;
wire n_10678;
wire n_6757;
wire n_17752;
wire n_18045;
wire n_8323;
wire n_10391;
wire n_13176;
wire n_9784;
wire n_19647;
wire n_7990;
wire n_18368;
wire n_10036;
wire n_17631;
wire n_14905;
wire n_15128;
wire n_8720;
wire n_12205;
wire n_11989;
wire n_16912;
wire n_16215;
wire n_14009;
wire n_15787;
wire n_19943;
wire n_7148;
wire n_9417;
wire n_12020;
wire n_18875;
wire n_6835;
wire n_11624;
wire n_20275;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_19290;
wire n_6247;
wire n_11234;
wire n_10919;
wire n_12099;
wire n_12858;
wire n_15351;
wire n_18170;
wire n_19159;
wire n_7544;
wire n_9336;
wire n_19750;
wire n_8854;
wire n_6645;
wire n_16177;
wire n_10727;
wire n_10885;
wire n_13201;
wire n_14759;
wire n_13274;
wire n_18621;
wire n_9312;
wire n_7469;
wire n_10895;
wire n_11977;
wire n_15576;
wire n_11696;
wire n_11734;
wire n_9533;
wire n_9494;
wire n_11507;
wire n_17290;
wire n_15337;
wire n_17276;
wire n_7082;
wire n_14749;
wire n_18731;
wire n_20000;
wire n_19306;
wire n_11320;
wire n_11837;
wire n_19458;
wire n_8260;
wire n_13898;
wire n_16507;
wire n_16543;
wire n_11938;
wire n_6418;
wire n_17003;
wire n_18814;
wire n_10571;
wire n_19202;
wire n_19664;
wire n_9807;
wire n_9057;
wire n_8706;
wire n_7945;
wire n_8894;
wire n_19244;
wire n_12053;
wire n_15947;
wire n_17738;
wire n_12619;
wire n_20488;
wire n_11289;
wire n_13555;
wire n_12582;
wire n_18919;
wire n_12423;
wire n_15426;
wire n_14137;
wire n_16905;
wire n_17765;
wire n_14163;
wire n_15523;
wire n_7328;
wire n_19298;
wire n_10958;
wire n_15682;
wire n_9479;
wire n_15556;
wire n_14041;
wire n_18622;
wire n_9181;
wire n_19338;
wire n_19385;
wire n_6578;
wire n_14763;
wire n_19319;
wire n_17686;
wire n_18381;
wire n_10879;
wire n_19481;
wire n_6589;
wire n_10639;
wire n_16359;
wire n_17448;
wire n_18657;
wire n_16037;
wire n_9276;
wire n_13351;
wire n_16805;
wire n_15937;
wire n_20453;
wire n_16141;
wire n_9821;
wire n_11112;
wire n_11723;
wire n_16647;
wire n_14393;
wire n_12364;
wire n_12420;
wire n_6567;
wire n_20574;
wire n_9508;
wire n_16231;
wire n_20423;
wire n_17805;
wire n_20181;
wire n_17318;
wire n_11906;
wire n_20586;
wire n_14298;
wire n_9741;
wire n_10180;
wire n_14112;
wire n_10650;
wire n_12120;
wire n_12021;
wire n_10157;
wire n_7423;
wire n_10402;
wire n_12515;
wire n_17283;
wire n_9166;
wire n_12895;
wire n_12045;
wire n_6940;
wire n_12726;
wire n_12668;
wire n_7835;
wire n_15437;
wire n_20536;
wire n_6320;
wire n_20570;
wire n_9969;
wire n_11437;
wire n_14068;
wire n_14853;
wire n_16735;
wire n_11869;
wire n_20214;
wire n_10836;
wire n_16375;
wire n_8072;
wire n_13117;
wire n_7130;
wire n_11282;
wire n_17720;
wire n_14700;
wire n_16382;
wire n_7491;
wire n_18944;
wire n_18474;
wire n_20636;
wire n_20138;
wire n_9636;
wire n_7559;
wire n_13175;
wire n_9833;
wire n_9095;
wire n_15757;
wire n_18465;
wire n_15979;
wire n_19076;
wire n_6731;
wire n_6154;
wire n_6943;
wire n_12038;
wire n_8210;
wire n_12644;
wire n_11826;
wire n_18241;
wire n_10888;
wire n_10116;
wire n_16764;
wire n_14808;
wire n_18135;
wire n_11764;
wire n_6600;
wire n_14140;
wire n_10696;
wire n_7355;
wire n_18688;
wire n_9331;
wire n_10170;
wire n_14479;
wire n_20183;
wire n_8331;
wire n_19883;
wire n_18109;
wire n_14172;
wire n_7270;
wire n_18721;
wire n_6967;
wire n_19241;
wire n_6742;
wire n_18117;
wire n_13525;
wire n_14997;
wire n_15931;
wire n_6691;
wire n_14799;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_19062;
wire n_12634;
wire n_14774;
wire n_12680;
wire n_11613;
wire n_10233;
wire n_19721;
wire n_15492;
wire n_18443;
wire n_17343;
wire n_10810;
wire n_12176;
wire n_10311;
wire n_9140;
wire n_18533;
wire n_19427;
wire n_12094;
wire n_9736;
wire n_12517;
wire n_6517;
wire n_18431;
wire n_15441;
wire n_9225;
wire n_17353;
wire n_11923;
wire n_12071;
wire n_13832;
wire n_8105;
wire n_9031;
wire n_19406;
wire n_13087;
wire n_13972;
wire n_15436;
wire n_17920;
wire n_15633;
wire n_19937;
wire n_12339;
wire n_10602;
wire n_16630;
wire n_14632;
wire n_6393;
wire n_15969;
wire n_8154;
wire n_13849;
wire n_11131;
wire n_10778;
wire n_17961;
wire n_19912;
wire n_13258;
wire n_9014;
wire n_13166;
wire n_8509;
wire n_6364;
wire n_16754;
wire n_15482;
wire n_16217;
wire n_19467;
wire n_11003;
wire n_18132;
wire n_12723;
wire n_19762;
wire n_14097;
wire n_18741;
wire n_19973;
wire n_8372;
wire n_17042;
wire n_10088;
wire n_20552;
wire n_14887;
wire n_7225;
wire n_8077;
wire n_18530;
wire n_20341;
wire n_16948;
wire n_6755;
wire n_18934;
wire n_13762;
wire n_13037;
wire n_11573;
wire n_10145;
wire n_7509;
wire n_14225;
wire n_11005;
wire n_6255;
wire n_18611;
wire n_19903;
wire n_6840;
wire n_17675;
wire n_8423;
wire n_9577;
wire n_19149;
wire n_12589;
wire n_14143;
wire n_6488;
wire n_8337;
wire n_7164;
wire n_14044;
wire n_17431;
wire n_18249;
wire n_18561;
wire n_18134;
wire n_17000;
wire n_12699;
wire n_12927;
wire n_16588;
wire n_8199;
wire n_17456;
wire n_8656;
wire n_14909;
wire n_10918;
wire n_13122;
wire n_15553;
wire n_12663;
wire n_16349;
wire n_17165;
wire n_20125;
wire n_15841;
wire n_17623;
wire n_11127;
wire n_18083;
wire n_7134;
wire n_9547;
wire n_16350;
wire n_8346;
wire n_8761;
wire n_15458;
wire n_9085;
wire n_13734;
wire n_8226;
wire n_17532;
wire n_7079;
wire n_9084;
wire n_20365;
wire n_14051;
wire n_20078;
wire n_17680;
wire n_9889;
wire n_12375;
wire n_12556;
wire n_13723;
wire n_10168;
wire n_12156;
wire n_13128;
wire n_13490;
wire n_17663;
wire n_14913;
wire n_10621;
wire n_9731;
wire n_6572;
wire n_9604;
wire n_7962;
wire n_15382;
wire n_20466;
wire n_7755;
wire n_16031;
wire n_6080;
wire n_8387;
wire n_12076;
wire n_10613;
wire n_6717;
wire n_7473;
wire n_20464;
wire n_11359;
wire n_19404;
wire n_19064;
wire n_15997;
wire n_19562;
wire n_10561;
wire n_19335;
wire n_14695;
wire n_16251;
wire n_13212;
wire n_16978;
wire n_15166;
wire n_18304;
wire n_15138;
wire n_16516;
wire n_18517;
wire n_17533;
wire n_14405;
wire n_7038;
wire n_14081;
wire n_8177;
wire n_17616;
wire n_12025;
wire n_8962;
wire n_9538;
wire n_14254;
wire n_16137;
wire n_6145;
wire n_6539;
wire n_6926;
wire n_13421;
wire n_13495;
wire n_13474;
wire n_14903;
wire n_13949;
wire n_12383;
wire n_11912;
wire n_14967;
wire n_9423;
wire n_16619;
wire n_20550;
wire n_12962;
wire n_18823;
wire n_16263;
wire n_11666;
wire n_12459;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_16369;
wire n_17213;
wire n_6710;
wire n_19745;
wire n_18326;
wire n_19402;
wire n_17664;
wire n_9056;
wire n_12496;
wire n_12814;
wire n_15943;
wire n_18714;
wire n_11921;
wire n_8495;
wire n_14532;
wire n_8783;
wire n_14557;
wire n_19805;
wire n_12603;
wire n_15392;
wire n_14340;
wire n_18444;
wire n_14032;
wire n_16944;
wire n_15702;
wire n_7262;
wire n_12967;
wire n_14899;
wire n_12232;
wire n_18115;
wire n_18847;
wire n_11859;
wire n_15773;
wire n_19771;
wire n_15307;
wire n_14111;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9553;
wire n_11633;
wire n_7506;
wire n_8551;
wire n_14361;
wire n_12760;
wire n_18291;
wire n_19633;
wire n_14943;
wire n_12590;
wire n_15605;
wire n_17711;
wire n_7142;
wire n_12577;
wire n_18951;
wire n_10182;
wire n_16813;
wire n_13928;
wire n_19342;
wire n_7125;
wire n_11655;
wire n_12069;
wire n_16899;
wire n_15656;
wire n_18455;
wire n_16957;
wire n_10317;
wire n_12270;
wire n_16021;
wire n_9196;
wire n_19934;
wire n_14555;
wire n_10893;
wire n_9251;
wire n_9973;
wire n_11117;
wire n_8064;
wire n_8468;
wire n_10201;
wire n_12210;
wire n_8778;
wire n_17106;
wire n_14168;
wire n_15342;
wire n_15534;
wire n_10539;
wire n_14080;
wire n_11777;
wire n_17402;
wire n_13975;
wire n_10121;
wire n_8198;
wire n_19054;
wire n_6828;
wire n_7255;
wire n_12189;
wire n_9270;
wire n_14142;
wire n_9099;
wire n_7350;
wire n_10814;
wire n_16034;
wire n_9627;
wire n_17008;
wire n_16563;
wire n_6664;
wire n_17575;
wire n_13131;
wire n_14941;
wire n_11154;
wire n_11700;
wire n_20428;
wire n_16128;
wire n_10975;
wire n_9460;
wire n_17698;
wire n_11652;
wire n_14320;
wire n_11056;
wire n_19229;
wire n_6238;
wire n_13932;
wire n_16804;
wire n_15606;
wire n_10459;
wire n_20501;
wire n_6545;
wire n_11583;
wire n_15866;
wire n_9766;
wire n_20041;
wire n_10463;
wire n_14764;
wire n_19897;
wire n_8734;
wire n_7074;
wire n_12564;
wire n_19443;
wire n_13433;
wire n_15505;
wire n_10403;
wire n_7037;
wire n_13697;
wire n_11784;
wire n_20549;
wire n_9025;
wire n_14244;
wire n_7928;
wire n_12886;
wire n_6532;
wire n_7293;
wire n_18638;
wire n_13000;
wire n_14362;
wire n_15996;
wire n_6721;
wire n_18825;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_18537;
wire n_9597;
wire n_11892;
wire n_15731;
wire n_19909;
wire n_8299;
wire n_12473;
wire n_11421;
wire n_11966;
wire n_18704;
wire n_19530;
wire n_17450;
wire n_18011;
wire n_12748;
wire n_16829;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_17305;
wire n_18047;
wire n_8188;
wire n_7078;
wire n_13831;
wire n_16792;
wire n_18572;
wire n_11423;
wire n_18378;
wire n_20211;
wire n_9567;
wire n_9061;
wire n_17154;
wire n_16922;
wire n_8664;
wire n_16552;
wire n_16867;
wire n_16638;
wire n_14783;
wire n_13268;
wire n_10740;
wire n_10457;
wire n_19042;
wire n_17968;
wire n_14158;
wire n_9701;
wire n_19247;
wire n_14236;
wire n_18849;
wire n_13510;
wire n_14640;
wire n_6659;
wire n_9709;
wire n_9295;
wire n_16678;
wire n_10264;
wire n_15029;
wire n_14286;
wire n_12528;
wire n_17640;
wire n_6182;
wire n_12717;
wire n_6520;
wire n_12660;
wire n_17651;
wire n_17662;
wire n_11547;
wire n_19680;
wire n_20273;
wire n_13520;
wire n_19668;
wire n_20028;
wire n_8501;
wire n_10301;
wire n_13018;
wire n_18240;
wire n_15139;
wire n_8076;
wire n_6826;
wire n_11395;
wire n_9107;
wire n_19630;
wire n_11279;
wire n_18370;
wire n_11724;
wire n_20429;
wire n_11789;
wire n_14152;
wire n_14869;
wire n_19989;
wire n_19354;
wire n_8014;
wire n_19030;
wire n_7768;
wire n_8638;
wire n_16294;
wire n_14651;
wire n_7982;
wire n_8804;
wire n_11383;
wire n_20598;
wire n_15882;
wire n_17740;
wire n_6879;
wire n_17059;
wire n_7567;
wire n_8433;
wire n_10932;
wire n_10619;
wire n_17263;
wire n_9156;
wire n_16113;
wire n_16848;
wire n_18749;
wire n_20082;
wire n_10248;
wire n_9748;
wire n_13365;
wire n_7771;
wire n_11780;
wire n_16289;
wire n_7701;
wire n_16342;
wire n_17278;
wire n_6720;
wire n_11930;
wire n_6888;
wire n_12628;
wire n_8122;
wire n_17095;
wire n_13444;
wire n_16504;
wire n_8432;
wire n_7592;
wire n_14209;
wire n_20305;
wire n_19462;
wire n_18651;
wire n_6590;
wire n_18243;
wire n_11876;
wire n_19110;
wire n_7151;
wire n_8950;
wire n_18683;
wire n_10758;
wire n_13431;
wire n_12538;
wire n_14025;
wire n_7758;
wire n_13779;
wire n_12446;
wire n_15954;
wire n_9355;
wire n_15386;
wire n_14620;
wire n_15349;
wire n_9582;
wire n_11009;
wire n_9288;
wire n_6308;
wire n_7897;
wire n_17701;
wire n_7118;
wire n_8284;
wire n_9702;
wire n_18767;
wire n_15378;
wire n_7422;
wire n_17881;
wire n_6738;
wire n_12307;
wire n_8703;
wire n_15839;
wire n_16135;
wire n_17661;
wire n_14999;
wire n_19377;
wire n_13720;
wire n_7339;
wire n_13706;
wire n_13903;
wire n_9051;
wire n_8545;
wire n_10385;
wire n_10105;
wire n_15785;
wire n_20530;
wire n_19056;
wire n_17114;
wire n_10251;
wire n_15234;
wire n_18796;
wire n_17524;
wire n_9980;
wire n_14394;
wire n_20098;
wire n_18679;
wire n_17261;
wire n_9555;
wire n_14845;
wire n_19906;
wire n_7713;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_16182;
wire n_19239;
wire n_10304;
wire n_6936;
wire n_15934;
wire n_16827;
wire n_16121;
wire n_7487;
wire n_9986;
wire n_13794;
wire n_13537;
wire n_9397;
wire n_18616;
wire n_17574;
wire n_9855;
wire n_10568;
wire n_13463;
wire n_9496;
wire n_16241;
wire n_10796;
wire n_10016;
wire n_10030;
wire n_12864;
wire n_9653;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_13936;
wire n_13933;
wire n_7815;
wire n_7934;
wire n_11578;
wire n_6865;
wire n_7276;
wire n_18595;
wire n_8739;
wire n_17078;
wire n_6747;
wire n_13714;
wire n_12725;
wire n_6640;
wire n_16030;
wire n_16079;
wire n_11908;
wire n_18166;
wire n_6462;
wire n_17372;
wire n_9781;
wire n_13159;
wire n_14788;
wire n_13287;
wire n_11913;
wire n_7034;
wire n_13389;
wire n_17726;
wire n_9906;
wire n_12317;
wire n_13302;
wire n_10092;
wire n_6833;
wire n_6793;
wire n_16766;
wire n_17834;
wire n_11815;
wire n_6295;
wire n_11231;
wire n_13740;
wire n_17966;
wire n_19278;
wire n_19926;
wire n_8137;
wire n_12027;
wire n_15218;
wire n_17366;
wire n_19114;
wire n_17514;
wire n_7014;
wire n_17975;
wire n_10430;
wire n_16697;
wire n_8305;
wire n_18147;
wire n_18751;
wire n_6709;
wire n_17525;
wire n_6712;
wire n_7416;
wire n_14553;
wire n_9657;
wire n_16594;
wire n_16370;
wire n_6743;
wire n_16223;
wire n_12412;
wire n_11880;
wire n_14528;
wire n_20150;
wire n_9485;
wire n_13940;
wire n_11249;
wire n_15449;
wire n_10119;
wire n_11986;
wire n_14798;
wire n_17579;
wire n_12118;
wire n_14409;
wire n_14724;
wire n_18451;
wire n_14291;
wire n_8625;
wire n_6919;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_19957;
wire n_9192;
wire n_20635;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_8179;
wire n_19360;
wire n_11861;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_7453;
wire n_10684;
wire n_18095;
wire n_15039;
wire n_17929;
wire n_17027;
wire n_8806;
wire n_17400;
wire n_6619;
wire n_19234;
wire n_16434;
wire n_20405;
wire n_13930;
wire n_8149;
wire n_10390;
wire n_20073;
wire n_7210;
wire n_6718;
wire n_15400;
wire n_17411;
wire n_16866;
wire n_15485;
wire n_18499;
wire n_18789;
wire n_14841;
wire n_16726;
wire n_13624;
wire n_18603;
wire n_19480;
wire n_8269;
wire n_13805;
wire n_18786;
wire n_8968;
wire n_16243;
wire n_7855;
wire n_14029;
wire n_14056;
wire n_13695;
wire n_6981;
wire n_13288;
wire n_19465;
wire n_16917;
wire n_11519;
wire n_13065;
wire n_11229;
wire n_18655;
wire n_16159;
wire n_17570;
wire n_11397;
wire n_12840;
wire n_12846;
wire n_14705;
wire n_17660;
wire n_8401;
wire n_7854;
wire n_10577;
wire n_11324;
wire n_12945;
wire n_17385;
wire n_10151;
wire n_6439;
wire n_8240;
wire n_12850;
wire n_7714;
wire n_16193;
wire n_9305;
wire n_9999;
wire n_17495;
wire n_11361;
wire n_6945;
wire n_18617;
wire n_7029;
wire n_19009;
wire n_20180;
wire n_10186;
wire n_17236;
wire n_11841;
wire n_6618;
wire n_14453;
wire n_19824;
wire n_19882;
wire n_20389;
wire n_17545;
wire n_13094;
wire n_7317;
wire n_17558;
wire n_9461;
wire n_6816;
wire n_10928;
wire n_6502;
wire n_6250;
wire n_6288;
wire n_7522;
wire n_9618;
wire n_6118;
wire n_18961;
wire n_19772;
wire n_11808;
wire n_17970;
wire n_13257;
wire n_17160;
wire n_18778;
wire n_18509;
wire n_17636;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_13922;
wire n_13423;
wire n_18149;
wire n_10252;
wire n_16641;
wire n_11555;
wire n_6869;
wire n_14625;
wire n_10345;
wire n_10059;
wire n_8325;
wire n_7621;
wire n_7359;
wire n_12394;
wire n_13578;
wire n_19540;
wire n_14204;
wire n_9005;
wire n_8274;
wire n_12954;
wire n_19703;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_14688;
wire n_10644;
wire n_12801;
wire n_18594;
wire n_13708;
wire n_10365;
wire n_11781;
wire n_20312;
wire n_9648;
wire n_12965;
wire n_12788;
wire n_9498;
wire n_15707;
wire n_16328;
wire n_20127;
wire n_15396;
wire n_19804;
wire n_15909;
wire n_11884;
wire n_20146;
wire n_19516;
wire n_19734;
wire n_13371;
wire n_7971;
wire n_12264;
wire n_8232;
wire n_9649;
wire n_8904;
wire n_16977;
wire n_19287;
wire n_10629;
wire n_7070;
wire n_8382;
wire n_18950;
wire n_13856;
wire n_15607;
wire n_15879;
wire n_7259;
wire n_12274;
wire n_14588;
wire n_19985;
wire n_8128;
wire n_15746;
wire n_15921;
wire n_19545;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_12586;
wire n_8794;
wire n_11760;
wire n_19203;
wire n_17222;
wire n_20505;
wire n_8205;
wire n_9907;
wire n_19887;
wire n_13088;
wire n_6976;
wire n_13538;
wire n_11024;
wire n_18437;
wire n_6304;
wire n_7640;
wire n_13701;
wire n_10498;
wire n_11424;
wire n_12585;
wire n_14021;
wire n_10635;
wire n_13626;
wire n_20403;
wire n_19218;
wire n_12832;
wire n_8067;
wire n_12301;
wire n_9643;
wire n_18973;
wire n_18402;
wire n_15822;
wire n_11881;
wire n_14980;
wire n_7727;
wire n_18968;
wire n_11935;
wire n_17561;
wire n_18766;
wire n_18901;
wire n_8719;
wire n_16140;
wire n_19223;
wire n_18046;
wire n_15493;
wire n_12615;
wire n_13357;
wire n_10802;
wire n_17148;
wire n_7565;
wire n_16624;
wire n_20225;
wire n_7631;
wire n_20614;
wire n_13869;
wire n_16903;
wire n_7387;
wire n_9212;
wire n_12167;
wire n_9473;
wire n_13026;
wire n_10490;
wire n_15019;
wire n_13499;
wire n_17107;
wire n_14843;
wire n_10647;
wire n_9320;
wire n_10523;
wire n_16781;
wire n_19738;
wire n_12298;
wire n_10081;
wire n_12569;
wire n_14929;
wire n_18497;
wire n_20288;
wire n_12456;
wire n_8655;
wire n_17039;
wire n_10808;
wire n_6333;
wire n_8745;
wire n_18504;
wire n_8086;
wire n_15466;
wire n_13943;
wire n_17124;
wire n_7379;
wire n_17530;
wire n_8901;
wire n_11078;
wire n_8695;
wire n_8173;
wire n_12072;
wire n_10545;
wire n_17945;
wire n_16557;
wire n_20093;
wire n_14141;
wire n_9379;
wire n_11992;
wire n_15790;
wire n_17061;
wire n_14880;
wire n_13142;
wire n_13180;
wire n_10453;
wire n_16975;
wire n_16716;
wire n_13785;
wire n_7742;
wire n_9274;
wire n_20395;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_17230;
wire n_12863;
wire n_10352;
wire n_19876;
wire n_19449;
wire n_16830;
wire n_17851;
wire n_8507;
wire n_8415;
wire n_10713;
wire n_6680;
wire n_10954;
wire n_7432;
wire n_16036;
wire n_13978;
wire n_13941;
wire n_15339;
wire n_13439;
wire n_16152;
wire n_14133;
wire n_14433;
wire n_13187;
wire n_13162;
wire n_7505;
wire n_18521;
wire n_15059;
wire n_8244;
wire n_7494;
wire n_18380;
wire n_17071;
wire n_13661;
wire n_9546;
wire n_7589;
wire n_17764;
wire n_19969;
wire n_11296;
wire n_13770;
wire n_18636;
wire n_8723;
wire n_13511;
wire n_18016;
wire n_11019;
wire n_7843;
wire n_19544;
wire n_19258;
wire n_14569;
wire n_7902;
wire n_6496;
wire n_15744;
wire n_7756;
wire n_15557;
wire n_18244;
wire n_8342;
wire n_8940;
wire n_14154;
wire n_8472;
wire n_10000;
wire n_12812;
wire n_7988;
wire n_14174;
wire n_7500;
wire n_10246;
wire n_18236;
wire n_14269;
wire n_9822;
wire n_13991;
wire n_17523;
wire n_14821;
wire n_17330;
wire n_15096;
wire n_14992;
wire n_10125;
wire n_9065;
wire n_16637;
wire n_18627;
wire n_9086;
wire n_9153;
wire n_10505;
wire n_11064;
wire n_6908;
wire n_8237;
wire n_9093;
wire n_19046;
wire n_7266;
wire n_17928;
wire n_8046;
wire n_13284;
wire n_16521;
wire n_9198;
wire n_20580;
wire n_8335;
wire n_9142;
wire n_17697;
wire n_15820;
wire n_18239;
wire n_15486;
wire n_9493;
wire n_19371;
wire n_11330;
wire n_12720;
wire n_7794;
wire n_19139;
wire n_20431;
wire n_13318;
wire n_15917;
wire n_6605;
wire n_19748;
wire n_12687;
wire n_18278;
wire n_17510;
wire n_19106;
wire n_13208;
wire n_13867;
wire n_15594;
wire n_17807;
wire n_17841;
wire n_11796;
wire n_18339;
wire n_16881;
wire n_12789;
wire n_12127;
wire n_17232;
wire n_16976;
wire n_8037;
wire n_13673;
wire n_14119;
wire n_16775;
wire n_12573;
wire n_19400;
wire n_15214;
wire n_13045;
wire n_19913;
wire n_17347;
wire n_18684;
wire n_6806;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_6960;
wire n_8169;
wire n_12265;
wire n_17777;
wire n_7504;
wire n_15971;
wire n_11678;
wire n_19814;
wire n_8023;
wire n_12251;
wire n_16307;
wire n_8130;
wire n_16911;
wire n_15294;
wire n_18676;
wire n_16288;
wire n_7116;
wire n_17992;
wire n_6999;
wire n_14741;
wire n_20436;
wire n_11046;
wire n_11079;
wire n_15581;
wire n_11065;
wire n_8339;
wire n_19058;
wire n_14215;
wire n_20290;
wire n_17368;
wire n_18104;
wire n_8499;
wire n_15356;
wire n_18525;
wire n_6882;
wire n_10775;
wire n_9526;
wire n_17511;
wire n_18762;
wire n_15571;
wire n_7983;
wire n_10863;
wire n_17138;
wire n_17700;
wire n_13993;
wire n_10986;
wire n_8366;
wire n_8102;
wire n_19126;
wire n_18087;
wire n_8022;
wire n_17226;
wire n_19212;
wire n_10262;
wire n_10239;
wire n_14577;
wire n_14984;
wire n_20514;
wire n_18183;
wire n_8913;
wire n_16772;
wire n_14699;
wire n_20074;
wire n_10335;
wire n_15362;
wire n_11301;
wire n_15101;
wire n_18154;
wire n_11703;
wire n_6374;
wire n_17013;
wire n_6628;
wire n_13483;
wire n_18923;
wire n_16551;
wire n_17803;
wire n_6570;
wire n_20358;
wire n_8556;
wire n_8040;
wire n_11821;
wire n_13121;
wire n_13989;
wire n_10755;
wire n_16998;
wire n_15200;
wire n_17349;
wire n_10682;
wire n_6371;
wire n_8079;
wire n_8595;
wire n_15887;
wire n_10022;
wire n_13803;
wire n_14066;
wire n_7856;
wire n_6148;
wire n_7625;
wire n_12775;
wire n_7863;
wire n_6989;
wire n_8958;
wire n_12833;
wire n_12090;
wire n_6896;
wire n_13687;
wire n_19852;
wire n_7623;
wire n_7217;
wire n_14540;
wire n_16784;
wire n_8115;
wire n_9398;
wire n_15320;
wire n_12915;
wire n_6196;
wire n_13149;
wire n_18748;
wire n_14091;
wire n_15755;
wire n_8412;
wire n_6485;
wire n_14478;
wire n_17848;
wire n_10177;
wire n_6107;
wire n_16689;
wire n_11944;
wire n_7796;
wire n_6994;
wire n_15986;
wire n_14570;
wire n_16068;
wire n_13797;
wire n_13013;
wire n_13238;
wire n_9446;
wire n_11129;
wire n_7234;
wire n_10296;
wire n_8119;
wire n_8641;
wire n_12988;
wire n_17136;
wire n_20524;
wire n_13344;
wire n_11139;
wire n_17766;
wire n_8436;
wire n_12685;
wire n_14239;
wire n_8659;
wire n_14045;
wire n_19575;
wire n_7849;
wire n_12667;
wire n_18747;
wire n_15635;
wire n_10018;
wire n_7297;
wire n_15183;
wire n_7298;
wire n_15118;
wire n_9129;
wire n_10141;
wire n_14162;
wire n_8224;
wire n_20522;
wire n_15679;
wire n_13014;
wire n_19744;
wire n_10897;
wire n_10449;
wire n_7861;
wire n_14303;
wire n_7039;
wire n_11349;
wire n_7077;
wire n_12540;
wire n_19160;
wire n_13239;
wire n_15942;
wire n_17583;
wire n_18552;
wire n_9143;
wire n_8287;
wire n_19967;
wire n_7950;
wire n_8607;
wire n_17032;
wire n_6248;
wire n_16768;
wire n_16134;
wire n_20149;
wire n_10452;
wire n_7806;
wire n_15928;
wire n_16092;
wire n_7595;
wire n_8066;
wire n_12349;
wire n_14282;
wire n_6715;
wire n_6714;
wire n_11308;
wire n_16266;
wire n_8416;
wire n_20070;
wire n_14167;
wire n_9113;
wire n_7149;
wire n_10363;
wire n_13623;
wire n_11511;
wire n_15833;
wire n_16046;
wire n_9393;
wire n_15974;
wire n_13845;
wire n_12709;
wire n_13432;
wire n_12771;
wire n_17760;
wire n_20523;
wire n_14787;
wire n_19502;
wire n_7303;
wire n_6616;
wire n_17100;
wire n_10781;
wire n_7315;
wire n_9886;
wire n_13244;
wire n_18969;
wire n_6185;
wire n_10943;
wire n_12344;
wire n_13843;
wire n_17191;
wire n_13404;
wire n_18689;
wire n_7268;
wire n_10094;
wire n_16295;
wire n_10084;
wire n_19259;
wire n_13870;
wire n_13791;
wire n_6955;
wire n_9932;
wire n_16745;
wire n_13900;
wire n_16224;
wire n_14652;
wire n_8741;
wire n_7232;
wire n_7377;
wire n_19461;
wire n_16132;
wire n_19425;
wire n_6646;
wire n_19789;
wire n_15149;
wire n_14844;
wire n_16907;
wire n_14391;
wire n_11541;
wire n_15495;
wire n_9801;
wire n_19312;
wire n_8773;
wire n_6369;
wire n_19837;
wire n_8394;
wire n_11155;
wire n_7542;
wire n_13213;
wire n_12231;
wire n_17643;
wire n_8410;
wire n_14756;
wire n_18144;
wire n_7739;
wire n_19474;
wire n_14384;
wire n_15905;
wire n_12552;
wire n_11069;
wire n_16795;
wire n_9941;
wire n_20282;
wire n_17131;
wire n_11369;
wire n_14210;
wire n_20637;
wire n_15788;
wire n_13362;
wire n_7010;
wire n_9728;
wire n_16690;
wire n_20111;
wire n_7219;
wire n_9662;
wire n_12896;
wire n_15694;
wire n_8774;
wire n_18690;
wire n_19494;
wire n_7299;
wire n_9936;
wire n_6195;
wire n_9530;
wire n_14692;
wire n_7471;
wire n_10455;
wire n_15488;
wire n_11393;
wire n_7741;
wire n_9466;
wire n_16525;
wire n_7790;
wire n_16315;
wire n_19283;
wire n_6149;
wire n_17918;
wire n_7002;
wire n_12428;
wire n_15814;
wire n_10265;
wire n_16676;
wire n_18736;
wire n_15756;
wire n_19495;
wire n_11995;
wire n_14378;
wire n_18299;
wire n_11371;
wire n_14191;
wire n_19267;
wire n_16546;
wire n_18252;
wire n_17454;
wire n_16144;
wire n_16669;
wire n_6902;
wire n_10100;
wire n_18607;
wire n_15743;
wire n_7478;
wire n_19587;
wire n_19130;
wire n_7456;
wire n_13600;
wire n_8503;
wire n_8196;
wire n_16062;
wire n_17712;
wire n_9787;
wire n_10846;
wire n_13363;
wire n_19648;
wire n_9786;
wire n_18681;
wire n_14908;
wire n_12908;
wire n_18692;
wire n_17168;
wire n_14201;
wire n_8923;
wire n_13315;
wire n_18900;
wire n_6736;
wire n_19231;
wire n_14597;
wire n_15663;
wire n_9115;
wire n_11833;
wire n_11897;
wire n_19675;
wire n_7443;
wire n_11285;
wire n_9977;
wire n_8051;
wire n_16719;
wire n_9242;
wire n_11262;
wire n_12880;
wire n_8651;
wire n_13959;
wire n_10732;
wire n_6885;
wire n_10851;
wire n_10221;
wire n_9299;
wire n_11162;
wire n_13685;
wire n_14693;
wire n_8842;
wire n_19780;
wire n_16915;
wire n_14486;
wire n_7730;
wire n_11592;
wire n_15090;
wire n_8467;
wire n_17043;
wire n_15385;
wire n_16094;
wire n_6417;
wire n_13281;
wire n_15627;
wire n_10996;
wire n_8676;
wire n_9853;
wire n_13192;
wire n_7448;
wire n_17170;
wire n_19045;
wire n_17351;
wire n_18060;
wire n_15048;
wire n_16393;
wire n_17135;
wire n_20292;
wire n_6199;
wire n_9823;
wire n_15739;
wire n_12937;
wire n_10698;
wire n_16891;
wire n_18118;
wire n_14665;
wire n_6726;
wire n_7011;
wire n_10870;
wire n_11066;
wire n_17327;
wire n_13886;
wire n_16887;
wire n_6576;
wire n_8906;
wire n_17117;
wire n_8482;
wire n_7952;
wire n_16242;
wire n_14489;
wire n_13774;
wire n_13847;
wire n_6915;
wire n_19645;
wire n_12529;
wire n_20414;
wire n_12103;
wire n_7834;
wire n_17072;
wire n_8409;
wire n_17889;
wire n_14053;
wire n_19321;
wire n_8930;
wire n_16564;
wire n_14581;
wire n_18811;
wire n_7890;
wire n_11950;
wire n_12461;
wire n_11415;
wire n_7265;
wire n_7986;
wire n_17809;
wire n_17900;
wire n_9879;
wire n_18744;
wire n_11390;
wire n_20021;
wire n_17238;
wire n_11669;
wire n_14712;
wire n_15717;
wire n_8250;
wire n_10601;
wire n_9158;
wire n_18591;
wire n_16945;
wire n_7717;
wire n_9518;
wire n_18187;
wire n_18462;
wire n_18260;
wire n_11739;
wire n_10497;
wire n_14561;
wire n_18405;
wire n_13301;
wire n_8298;
wire n_7860;
wire n_14212;
wire n_7335;
wire n_9815;
wire n_13158;
wire n_11044;
wire n_15967;
wire n_15530;
wire n_11679;
wire n_8450;
wire n_17665;
wire n_17799;
wire n_7499;
wire n_19718;
wire n_7292;
wire n_12398;
wire n_17089;
wire n_9043;
wire n_7397;
wire n_10789;
wire n_17020;
wire n_12705;
wire n_7977;
wire n_12847;
wire n_13047;
wire n_6861;
wire n_14470;
wire n_15497;
wire n_7847;
wire n_15952;
wire n_13178;
wire n_19777;
wire n_18609;
wire n_12404;
wire n_11606;
wire n_19817;
wire n_11452;
wire n_15734;
wire n_6217;
wire n_20152;
wire n_10797;
wire n_7289;
wire n_17656;
wire n_14110;
wire n_14806;
wire n_7354;
wire n_18312;
wire n_13824;
wire n_7960;
wire n_15620;
wire n_18053;
wire n_12912;
wire n_12211;
wire n_6115;
wire n_13377;
wire n_16493;
wire n_6416;
wire n_6838;
wire n_10068;
wire n_11988;
wire n_19927;
wire n_19034;
wire n_6256;
wire n_15645;
wire n_6613;
wire n_11438;
wire n_15965;
wire n_18877;
wire n_6361;
wire n_14981;
wire n_11348;
wire n_9685;
wire n_11685;
wire n_6678;
wire n_8662;
wire n_15058;
wire n_16539;
wire n_14971;
wire n_19801;
wire n_12429;
wire n_14734;
wire n_20265;
wire n_14494;
wire n_14956;
wire n_7325;
wire n_14866;
wire n_19123;
wire n_6370;
wire n_9923;
wire n_13743;
wire n_7166;
wire n_7356;
wire n_13378;
wire n_11319;
wire n_16981;
wire n_7873;
wire n_16418;
wire n_20189;
wire n_19363;
wire n_17795;
wire n_12640;
wire n_10063;
wire n_13092;
wire n_14292;
wire n_20289;
wire n_8419;
wire n_19497;
wire n_9862;
wire n_11385;
wire n_11355;
wire n_18659;
wire n_11674;
wire n_12535;
wire n_19031;
wire n_12327;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_8430;
wire n_15719;
wire n_12058;
wire n_14879;
wire n_16143;
wire n_18387;
wire n_15164;
wire n_7052;
wire n_16755;
wire n_10496;
wire n_14149;
wire n_18225;
wire n_9960;
wire n_10998;
wire n_19180;
wire n_7502;
wire n_14216;
wire n_16380;
wire n_7919;
wire n_20554;
wire n_10800;
wire n_17962;
wire n_7085;
wire n_12065;
wire n_13950;
wire n_18952;
wire n_13732;
wire n_16422;
wire n_14968;
wire n_10993;
wire n_15542;
wire n_14985;
wire n_15910;
wire n_20267;
wire n_17734;
wire n_14443;
wire n_16136;
wire n_14285;
wire n_9734;
wire n_7288;
wire n_16325;
wire n_16842;
wire n_17355;
wire n_20281;
wire n_10495;
wire n_9004;
wire n_19981;
wire n_6610;
wire n_10612;
wire n_10260;
wire n_12285;
wire n_6750;
wire n_9150;
wire n_14508;
wire n_15092;
wire n_20259;
wire n_12683;
wire n_18535;
wire n_19691;
wire n_18457;
wire n_14566;
wire n_7869;
wire n_7165;
wire n_13386;
wire n_13846;
wire n_7683;
wire n_16437;
wire n_9587;
wire n_10671;
wire n_10193;
wire n_11718;
wire n_19333;
wire n_14383;
wire n_16695;
wire n_11680;
wire n_14683;
wire n_18685;
wire n_17052;
wire n_7322;
wire n_17378;
wire n_11658;
wire n_12226;
wire n_13492;
wire n_14001;
wire n_15397;
wire n_15840;
wire n_7880;
wire n_20567;
wire n_16855;
wire n_19120;
wire n_16937;
wire n_9919;
wire n_12135;
wire n_19485;
wire n_17092;
wire n_8829;
wire n_19308;
wire n_13381;
wire n_8971;
wire n_18076;
wire n_16667;
wire n_16897;
wire n_10558;
wire n_9579;
wire n_9475;
wire n_17603;
wire n_20366;
wire n_15273;
wire n_9049;
wire n_13718;
wire n_18701;
wire n_14775;
wire n_18809;
wire n_11045;
wire n_16756;
wire n_11340;
wire n_16965;
wire n_7675;
wire n_11903;
wire n_13279;
wire n_20410;
wire n_19704;
wire n_13644;
wire n_20242;
wire n_13291;
wire n_10174;
wire n_20324;
wire n_7524;
wire n_15897;
wire n_11564;
wire n_14015;
wire n_8925;
wire n_12946;
wire n_16729;
wire n_18406;
wire n_13513;
wire n_12916;
wire n_8471;
wire n_12521;
wire n_18925;
wire n_9800;
wire n_11382;
wire n_19578;
wire n_10098;
wire n_11745;
wire n_15240;
wire n_15564;
wire n_17002;
wire n_14350;
wire n_7733;
wire n_17405;
wire n_18711;
wire n_19090;
wire n_13773;
wire n_14109;
wire n_6982;
wire n_20117;
wire n_7345;
wire n_17526;
wire n_14136;
wire n_7385;
wire n_10923;
wire n_20528;
wire n_14176;
wire n_11149;
wire n_19889;
wire n_12635;
wire n_8488;
wire n_9543;
wire n_11443;
wire n_15765;
wire n_6855;
wire n_18176;
wire n_10665;
wire n_12906;
wire n_13467;
wire n_18374;
wire n_18700;
wire n_7907;
wire n_6312;
wire n_11532;
wire n_9415;
wire n_14343;
wire n_18619;
wire n_9147;
wire n_11209;
wire n_15918;
wire n_16212;
wire n_11790;
wire n_19189;
wire n_19444;
wire n_18148;
wire n_16313;
wire n_10420;
wire n_17058;
wire n_18309;
wire n_16363;
wire n_6131;
wire n_15232;
wire n_20491;
wire n_12105;
wire n_14329;
wire n_19392;
wire n_15721;
wire n_10444;
wire n_11377;
wire n_8018;
wire n_18557;
wire n_7937;
wire n_9176;
wire n_20103;
wire n_7819;
wire n_10631;
wire n_7305;
wire n_6334;
wire n_16780;
wire n_8884;
wire n_19222;
wire n_20171;
wire n_8751;
wire n_11864;
wire n_11006;
wire n_15018;
wire n_6617;
wire n_7511;
wire n_6533;
wire n_14108;
wire n_19829;
wire n_15439;
wire n_16049;
wire n_19875;
wire n_8178;
wire n_14000;
wire n_14372;
wire n_17911;
wire n_12046;
wire n_10212;
wire n_18566;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_11172;
wire n_10089;
wire n_14947;
wire n_8560;
wire n_14748;
wire n_18895;
wire n_20068;
wire n_19722;
wire n_18466;
wire n_10004;
wire n_12488;
wire n_11110;
wire n_17338;
wire n_16211;
wire n_15001;
wire n_8674;
wire n_12977;
wire n_7584;
wire n_13328;
wire n_10892;
wire n_18556;
wire n_10493;
wire n_19195;
wire n_10405;
wire n_15037;
wire n_17386;
wire n_7964;
wire n_17091;
wire n_14349;
wire n_6278;
wire n_7022;
wire n_12691;
wire n_11033;
wire n_19760;
wire n_19072;
wire n_18203;
wire n_14356;
wire n_19028;
wire n_16926;
wire n_16006;
wire n_12651;
wire n_19194;
wire n_16476;
wire n_7486;
wire n_6756;
wire n_16373;
wire n_18792;
wire n_14190;
wire n_8563;
wire n_17223;
wire n_15546;
wire n_11534;
wire n_14157;
wire n_14344;
wire n_9221;
wire n_7906;
wire n_6411;
wire n_10285;
wire n_14488;
wire n_11032;
wire n_13582;
wire n_17950;
wire n_7302;
wire n_18162;
wire n_20633;
wire n_19725;
wire n_11174;
wire n_18574;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_18544;
wire n_10294;
wire n_10106;
wire n_17865;
wire n_9934;
wire n_9234;
wire n_10674;
wire n_6534;
wire n_16011;
wire n_6265;
wire n_18185;
wire n_8087;
wire n_7607;
wire n_14458;
wire n_17540;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_20543;
wire n_13565;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_18965;
wire n_13784;
wire n_13468;
wire n_12363;
wire n_18201;
wire n_7553;
wire n_6824;
wire n_19625;
wire n_11788;
wire n_12544;
wire n_20240;
wire n_13036;
wire n_20496;
wire n_14146;
wire n_13199;
wire n_20248;
wire n_6903;
wire n_13009;
wire n_10908;
wire n_10339;
wire n_9908;
wire n_9486;
wire n_13002;
wire n_13868;
wire n_7903;
wire n_18596;
wire n_11877;
wire n_8864;
wire n_7384;
wire n_18674;
wire n_13285;
wire n_20476;
wire n_8610;
wire n_19075;
wire n_7894;
wire n_11750;
wire n_7055;
wire n_18722;
wire n_8520;
wire n_16458;
wire n_13374;
wire n_12055;
wire n_7639;
wire n_16520;
wire n_20231;
wire n_12811;
wire n_12186;
wire n_13032;
wire n_11001;
wire n_9512;
wire n_14199;
wire n_17858;
wire n_13684;
wire n_9170;
wire n_15108;
wire n_9616;
wire n_16898;
wire n_9073;
wire n_12897;
wire n_18325;
wire n_12272;
wire n_9302;
wire n_19068;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_9171;
wire n_8279;
wire n_12191;
wire n_17432;
wire n_9580;
wire n_8019;
wire n_13963;
wire n_17707;
wire n_18842;
wire n_7832;
wire n_9540;
wire n_17242;
wire n_11137;
wire n_8390;
wire n_8898;
wire n_14316;
wire n_8613;
wire n_18300;
wire n_8464;
wire n_15701;
wire n_6423;
wire n_15612;
wire n_18804;
wire n_7441;
wire n_12112;
wire n_13060;
wire n_16187;
wire n_9449;
wire n_19787;
wire n_14817;
wire n_9050;
wire n_6121;
wire n_14087;
wire n_15980;
wire n_20066;
wire n_14438;
wire n_16253;
wire n_7133;
wire n_12202;
wire n_13836;
wire n_8661;
wire n_7424;
wire n_19774;
wire n_16671;
wire n_12870;
wire n_11156;
wire n_10611;
wire n_10715;
wire n_12333;
wire n_8609;
wire n_17666;
wire n_17219;
wire n_7626;
wire n_13576;
wire n_7310;
wire n_17451;
wire n_12119;
wire n_12618;
wire n_16093;
wire n_17266;
wire n_20213;
wire n_15129;
wire n_17146;
wire n_16209;
wire n_14306;
wire n_8873;
wire n_11891;
wire n_16276;
wire n_18427;
wire n_12401;
wire n_13055;
wire n_7323;
wire n_7301;
wire n_18600;
wire n_17633;
wire n_13829;
wire n_16533;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_20577;
wire n_17815;
wire n_7244;
wire n_10745;
wire n_7633;
wire n_18760;
wire n_13937;
wire n_9437;
wire n_18724;
wire n_8640;
wire n_14359;
wire n_6186;
wire n_16933;
wire n_6803;
wire n_8437;
wire n_8427;
wire n_10605;
wire n_14013;
wire n_14419;
wire n_9933;
wire n_11449;
wire n_15251;
wire n_9892;
wire n_18976;
wire n_16727;
wire n_9462;
wire n_19447;
wire n_15854;
wire n_19438;
wire n_12501;
wire n_17518;
wire n_8843;
wire n_9891;
wire n_15810;
wire n_10643;
wire n_16974;
wire n_10872;
wire n_13987;
wire n_15626;
wire n_13416;
wire n_12798;
wire n_14885;
wire n_9925;
wire n_16066;
wire n_9757;
wire n_10008;
wire n_13726;
wire n_14412;
wire n_17587;
wire n_12243;
wire n_8562;
wire n_19714;
wire n_12614;
wire n_11378;
wire n_14631;
wire n_10032;
wire n_13425;
wire n_9806;
wire n_17105;
wire n_17233;
wire n_7021;
wire n_13591;
wire n_18296;
wire n_11713;
wire n_16972;
wire n_15586;
wire n_6355;
wire n_17821;
wire n_12931;
wire n_15525;
wire n_7215;
wire n_17790;
wire n_17566;
wire n_14332;
wire n_18379;
wire n_8016;
wire n_10645;
wire n_11096;
wire n_10604;
wire n_17398;
wire n_6564;
wire n_11161;
wire n_8709;
wire n_12491;
wire n_11216;
wire n_14368;
wire n_18390;
wire n_10966;
wire n_19310;
wire n_19871;
wire n_20110;
wire n_19650;
wire n_6442;
wire n_18359;
wire n_7925;
wire n_15126;
wire n_19289;
wire n_20097;
wire n_6871;
wire n_16846;
wire n_9389;
wire n_12074;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_19665;
wire n_12745;
wire n_9752;
wire n_14473;
wire n_12887;
wire n_18997;
wire n_10341;
wire n_19521;
wire n_15816;
wire n_18314;
wire n_7138;
wire n_17341;
wire n_8712;
wire n_19254;
wire n_20363;
wire n_8837;
wire n_17652;
wire n_14641;
wire n_16506;
wire n_17543;
wire n_15433;
wire n_15953;
wire n_9721;
wire n_11344;
wire n_12658;
wire n_9197;
wire n_19167;
wire n_14740;
wire n_9210;
wire n_6893;
wire n_8905;
wire n_13008;
wire n_18832;
wire n_18691;
wire n_7807;
wire n_18126;
wire n_14198;
wire n_14846;
wire n_9917;
wire n_12056;
wire n_14539;
wire n_8106;
wire n_20381;
wire n_12238;
wire n_19226;
wire n_12976;
wire n_14420;
wire n_18562;
wire n_11888;
wire n_13243;
wire n_14314;
wire n_16642;
wire n_14227;
wire n_10309;
wire n_11099;
wire n_8974;
wire n_14164;
wire n_10050;
wire n_9871;
wire n_19652;
wire n_19996;
wire n_10306;
wire n_7606;
wire n_7193;
wire n_18180;
wire n_18142;
wire n_13632;
wire n_13020;
wire n_13148;
wire n_10429;
wire n_11470;
wire n_13871;
wire n_20387;
wire n_9903;
wire n_17208;
wire n_11102;
wire n_9228;
wire n_11539;
wire n_7710;
wire n_17792;
wire n_16166;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_9522;
wire n_15617;
wire n_15463;
wire n_11076;
wire n_14339;
wire n_16005;
wire n_6769;
wire n_9148;
wire n_11054;
wire n_10754;
wire n_9275;
wire n_10223;
wire n_8896;
wire n_19727;
wire n_7206;
wire n_6895;
wire n_13598;
wire n_17979;
wire n_10228;
wire n_8758;
wire n_8617;
wire n_17953;
wire n_13966;
wire n_12530;
wire n_9463;
wire n_13077;
wire n_16309;
wire n_10425;
wire n_8069;
wire n_6481;
wire n_19144;
wire n_15201;
wire n_9997;
wire n_6384;
wire n_13828;
wire n_7541;
wire n_6906;
wire n_14562;
wire n_9844;
wire n_12826;
wire n_8318;
wire n_10366;
wire n_15015;
wire n_19122;
wire n_7334;
wire n_20280;
wire n_16376;
wire n_14991;
wire n_10225;
wire n_6257;
wire n_20490;
wire n_20360;
wire n_8383;
wire n_12621;
wire n_11290;
wire n_17080;
wire n_12518;
wire n_19033;
wire n_14047;
wire n_9052;
wire n_17447;
wire n_17678;
wire n_6587;
wire n_7781;
wire n_7360;
wire n_14568;
wire n_11702;
wire n_19395;
wire n_16970;
wire n_11372;
wire n_20424;
wire n_10817;
wire n_15324;
wire n_8355;
wire n_19501;
wire n_17098;
wire n_12741;
wire n_18041;
wire n_7101;
wire n_7530;
wire n_15006;
wire n_20113;
wire n_15619;
wire n_19914;
wire n_20460;
wire n_18911;
wire n_9860;
wire n_12510;
wire n_11756;
wire n_8369;
wire n_9022;
wire n_9103;
wire n_17142;
wire n_8831;
wire n_12233;
wire n_8853;
wire n_6252;
wire n_18403;
wire n_6211;
wire n_15716;
wire n_17499;
wire n_17898;
wire n_17172;
wire n_8081;
wire n_16608;
wire n_17310;
wire n_13442;
wire n_14444;
wire n_18531;
wire n_10484;
wire n_11744;
wire n_17247;
wire n_10288;
wire n_18838;
wire n_10388;
wire n_6189;
wire n_20209;
wire n_15299;
wire n_11072;
wire n_19836;
wire n_13944;
wire n_9492;
wire n_6413;
wire n_7419;
wire n_6506;
wire n_18476;
wire n_17086;
wire n_9727;
wire n_6935;
wire n_13019;
wire n_12703;
wire n_13079;
wire n_18343;
wire n_15369;
wire n_15134;
wire n_16110;
wire n_19420;
wire n_9375;
wire n_17715;
wire n_8770;
wire n_15453;
wire n_6105;
wire n_10964;
wire n_19739;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_7841;
wire n_9458;
wire n_20335;
wire n_8466;
wire n_6527;
wire n_15275;
wire n_19092;
wire n_8094;
wire n_6430;
wire n_18268;
wire n_10987;
wire n_12684;
wire n_20473;
wire n_11965;
wire n_14696;
wire n_15093;
wire n_12324;
wire n_14006;
wire n_6666;
wire n_8321;
wire n_20126;
wire n_19116;
wire n_9954;
wire n_8735;
wire n_11722;
wire n_12310;
wire n_6594;
wire n_19471;
wire n_20197;
wire n_7095;
wire n_16672;
wire n_11701;
wire n_18010;
wire n_13917;
wire n_7184;
wire n_9617;
wire n_13546;
wire n_14595;
wire n_17001;
wire n_7908;
wire n_7974;
wire n_7551;
wire n_11980;
wire n_11255;
wire n_13592;
wire n_17224;
wire n_11720;
wire n_20269;
wire n_13874;
wire n_6482;
wire n_15506;
wire n_9810;
wire n_14469;
wire n_16201;
wire n_17690;
wire n_8043;
wire n_16377;
wire n_14492;
wire n_14134;
wire n_11990;
wire n_10103;
wire n_15457;
wire n_14345;
wire n_16847;
wire n_6841;
wire n_10153;
wire n_17622;
wire n_17952;
wire n_8171;
wire n_20437;
wire n_9006;
wire n_19641;
wire n_6774;
wire n_16964;
wire n_8600;
wire n_14816;
wire n_8710;
wire n_12806;
wire n_14302;
wire n_8549;
wire n_10172;
wire n_8054;
wire n_13904;
wire n_16614;
wire n_18694;
wire n_17045;
wire n_15784;
wire n_18613;
wire n_11969;
wire n_7914;
wire n_16388;
wire n_6521;
wire n_8857;
wire n_14243;
wire n_9040;
wire n_6162;
wire n_8010;
wire n_6432;
wire n_13574;
wire n_12762;
wire n_16740;
wire n_9830;
wire n_18870;
wire n_10761;
wire n_18781;
wire n_11579;
wire n_15303;
wire n_8291;
wire n_18017;
wire n_20143;
wire n_11535;
wire n_18400;
wire n_12975;
wire n_16291;
wire n_13850;
wire n_6740;
wire n_11510;
wire n_6315;
wire n_17866;
wire n_12736;
wire n_9111;
wire n_7156;
wire n_9163;
wire n_15461;
wire n_6910;
wire n_6262;
wire n_14800;
wire n_7703;
wire n_6319;
wire n_17352;
wire n_14888;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_6536;
wire n_6175;
wire n_7040;
wire n_8280;
wire n_12390;
wire n_18898;
wire n_10235;
wire n_6978;
wire n_12805;
wire n_6093;
wire n_11649;
wire n_16306;
wire n_18485;
wire n_9190;
wire n_6947;
wire n_14918;
wire n_8203;
wire n_6099;
wire n_20478;
wire n_6140;
wire n_15489;
wire n_19980;
wire n_12914;
wire n_17159;
wire n_17721;
wire n_9506;
wire n_18440;
wire n_6415;
wire n_18883;
wire n_20311;
wire n_16542;
wire n_15158;
wire n_10828;
wire n_18866;
wire n_12300;
wire n_15389;
wire n_7549;
wire n_17308;
wire n_17425;
wire n_11281;
wire n_13056;
wire n_16019;
wire n_17732;
wire n_12337;
wire n_18520;
wire n_13466;
wire n_15082;
wire n_8871;
wire n_11114;
wire n_19442;
wire n_8418;
wire n_7740;
wire n_20417;
wire n_13050;
wire n_10860;
wire n_18259;
wire n_17517;
wire n_16208;
wire n_20627;
wire n_19327;
wire n_15209;
wire n_12273;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_12712;
wire n_15078;
wire n_13012;
wire n_19895;
wire n_8924;
wire n_20134;
wire n_20500;
wire n_12752;
wire n_6928;
wire n_10880;
wire n_15511;
wire n_19600;
wire n_18204;
wire n_20081;
wire n_14278;
wire n_8214;
wire n_12777;
wire n_14706;
wire n_20278;
wire n_20302;
wire n_7043;
wire n_11462;
wire n_11732;
wire n_18137;
wire n_12819;
wire n_10214;
wire n_8241;
wire n_8442;
wire n_9572;
wire n_15282;
wire n_9229;
wire n_19505;
wire n_16812;
wire n_16038;
wire n_12237;
wire n_18350;
wire n_6134;
wire n_13372;
wire n_11375;
wire n_11267;
wire n_9602;
wire n_9311;
wire n_19482;
wire n_6593;
wire n_8630;
wire n_19432;
wire n_9884;
wire n_9876;
wire n_9260;
wire n_14534;
wire n_19832;
wire n_13630;
wire n_16535;
wire n_13700;
wire n_10406;
wire n_17859;
wire n_6746;
wire n_11985;
wire n_8447;
wire n_6443;
wire n_14290;
wire n_7980;
wire n_8828;
wire n_18631;
wire n_17687;
wire n_19820;
wire n_6749;
wire n_10965;
wire n_10798;
wire n_19657;
wire n_7732;
wire n_13325;
wire n_14850;
wire n_15135;
wire n_20338;
wire n_16196;
wire n_11911;
wire n_11442;
wire n_18862;
wire n_14064;
wire n_14524;
wire n_8859;
wire n_16883;
wire n_11388;
wire n_11651;
wire n_17946;
wire n_10154;
wire n_18663;
wire n_7922;
wire n_17469;
wire n_15826;
wire n_19101;
wire n_10033;
wire n_17877;
wire n_8311;
wire n_12253;
wire n_15005;
wire n_11147;
wire n_12928;
wire n_9877;
wire n_8764;
wire n_19361;
wire n_16167;
wire n_19452;
wire n_12990;
wire n_20239;
wire n_14246;
wire n_6920;
wire n_19902;
wire n_11817;
wire n_8729;
wire n_10359;
wire n_20384;
wire n_14957;
wire n_13447;
wire n_6907;
wire n_7144;
wire n_16579;
wire n_11479;
wire n_11737;
wire n_8048;
wire n_12028;
wire n_7072;
wire n_13095;
wire n_8253;
wire n_18592;
wire n_15032;
wire n_11600;
wire n_16607;
wire n_15085;
wire n_16390;
wire n_10722;
wire n_8088;
wire n_17855;
wire n_10666;
wire n_15440;
wire n_8516;
wire n_8302;
wire n_17717;
wire n_20042;
wire n_15610;
wire n_15329;
wire n_8167;
wire n_7859;
wire n_14315;
wire n_7872;
wire n_13858;
wire n_17913;
wire n_7480;
wire n_16255;
wire n_8944;
wire n_10023;
wire n_10999;
wire n_18716;
wire n_10410;
wire n_19732;
wire n_16983;
wire n_8975;
wire n_17009;
wire n_19888;
wire n_11305;
wire n_17668;
wire n_9101;
wire n_15631;
wire n_14755;
wire n_8825;
wire n_12969;
wire n_12260;
wire n_12016;
wire n_8266;
wire n_8981;
wire n_17082;
wire n_8771;
wire n_15750;
wire n_12939;
wire n_20533;
wire n_20419;
wire n_15038;
wire n_17925;
wire n_10404;
wire n_8138;
wire n_6638;
wire n_12779;
wire n_17505;
wire n_17199;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_9211;
wire n_8124;
wire n_7366;
wire n_9395;
wire n_17348;
wire n_8147;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_10700;
wire n_17743;
wire n_10968;
wire n_14247;
wire n_9716;
wire n_16155;
wire n_15418;
wire n_11970;
wire n_7918;
wire n_6651;
wire n_12308;
wire n_10783;
wire n_12163;
wire n_11523;
wire n_12944;
wire n_7472;
wire n_9737;
wire n_10812;
wire n_14709;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_19847;
wire n_10001;
wire n_13280;
wire n_12145;
wire n_11088;
wire n_8160;
wire n_20129;
wire n_11405;
wire n_19274;
wire n_13103;
wire n_18385;
wire n_15630;
wire n_10977;
wire n_11299;
wire n_10615;
wire n_11542;
wire n_7647;
wire n_12426;
wire n_16222;
wire n_15068;
wire n_15442;
wire n_9054;
wire n_10532;
wire n_17776;
wire n_13995;
wire n_13073;
wire n_6728;
wire n_19907;
wire n_20139;
wire n_16029;
wire n_13556;
wire n_13367;
wire n_10771;
wire n_11441;
wire n_14203;
wire n_17269;
wire n_19802;
wire n_12844;
wire n_7073;
wire n_9755;
wire n_10104;
wire n_9117;
wire n_19426;
wire n_9381;
wire n_12049;
wire n_14498;
wire n_6549;
wire n_19708;
wire n_20398;
wire n_6096;
wire n_7853;
wire n_12526;
wire n_8890;
wire n_16575;
wire n_7721;
wire n_7192;
wire n_19602;
wire n_20279;
wire n_11206;
wire n_11593;
wire n_15807;
wire n_11786;
wire n_12737;
wire n_17258;
wire n_15113;
wire n_9273;
wire n_8970;
wire n_16910;
wire n_10640;
wire n_10729;
wire n_14656;
wire n_20194;
wire n_16052;
wire n_20507;
wire n_14745;
wire n_20375;
wire n_19243;
wire n_7635;
wire n_19712;
wire n_11268;
wire n_17121;
wire n_14760;
wire n_20589;
wire n_11501;
wire n_7227;
wire n_13390;
wire n_8030;
wire n_8687;
wire n_13264;
wire n_12010;
wire n_9738;
wire n_12026;
wire n_17481;
wire n_8633;
wire n_17645;
wire n_19999;
wire n_7689;
wire n_6511;
wire n_18470;
wire n_7099;
wire n_14676;
wire n_6358;
wire n_18880;
wire n_11313;
wire n_10438;
wire n_6986;
wire n_8801;
wire n_16438;
wire n_8219;
wire n_15373;
wire n_18580;
wire n_10575;
wire n_11028;
wire n_12171;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_14906;
wire n_15211;
wire n_10760;
wire n_15334;
wire n_7731;
wire n_11527;
wire n_18404;
wire n_16486;
wire n_9535;
wire n_12490;
wire n_8486;
wire n_12829;
wire n_18662;
wire n_11610;
wire n_12739;
wire n_7132;
wire n_17021;
wire n_17710;
wire n_6663;
wire n_12609;
wire n_18248;
wire n_8155;
wire n_11360;
wire n_11868;
wire n_8098;
wire n_9191;
wire n_17791;
wire n_18202;
wire n_6376;
wire n_18141;
wire n_12888;
wire n_19407;
wire n_8485;
wire n_14852;
wire n_7001;
wire n_9650;
wire n_13070;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_14491;
wire n_15011;
wire n_17607;
wire n_9664;
wire n_20367;
wire n_14928;
wire n_13778;
wire n_9931;
wire n_16470;
wire n_16419;
wire n_16956;
wire n_14634;
wire n_10753;
wire n_13174;
wire n_7108;
wire n_14455;
wire n_17164;
wire n_11879;
wire n_7876;
wire n_17175;
wire n_20638;
wire n_9656;
wire n_8148;
wire n_8150;
wire n_20601;
wire n_12596;
wire n_15398;
wire n_15593;
wire n_18175;
wire n_16424;
wire n_13945;
wire n_8986;
wire n_19367;
wire n_20137;
wire n_12697;
wire n_7260;
wire n_6409;
wire n_11939;
wire n_14347;
wire n_7552;
wire n_19052;
wire n_17969;
wire n_12166;
wire n_10646;
wire n_15725;
wire n_11704;
wire n_20548;
wire n_17506;
wire n_18050;
wire n_8763;
wire n_8679;
wire n_7239;
wire n_15582;
wire n_16415;
wire n_9848;
wire n_14447;
wire n_11962;
wire n_9227;
wire n_7050;
wire n_17137;
wire n_6623;
wire n_13951;
wire n_13968;
wire n_10378;
wire n_16924;
wire n_13316;
wire n_10313;
wire n_13689;
wire n_8139;
wire n_17268;
wire n_18000;
wire n_19384;
wire n_19288;
wire n_19431;
wire n_10773;
wire n_18210;
wire n_8830;
wire n_14836;
wire n_12867;
wire n_15960;
wire n_7568;
wire n_15343;
wire n_6354;
wire n_6344;
wire n_12123;
wire n_9772;
wire n_18885;
wire n_15370;
wire n_7949;
wire n_7724;
wire n_18001;
wire n_6305;
wire n_12547;
wire n_16148;
wire n_20557;
wire n_15577;
wire n_16550;
wire n_19066;
wire n_8646;
wire n_13415;
wire n_10259;
wire n_7107;
wire n_17111;
wire n_6457;
wire n_8597;
wire n_17951;
wire n_17379;
wire n_7123;
wire n_8117;
wire n_15169;
wire n_10213;
wire n_13888;
wire n_16592;
wire n_8208;
wire n_19373;
wire n_20004;
wire n_8536;
wire n_17252;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_16475;
wire n_13892;
wire n_16361;
wire n_14559;
wire n_16831;
wire n_19696;
wire n_17110;
wire n_14052;
wire n_14311;
wire n_13765;
wire n_10332;
wire n_7709;
wire n_15290;
wire n_11874;
wire n_13926;
wire n_10171;
wire n_15184;
wire n_18131;
wire n_6386;
wire n_12803;
wire n_19518;
wire n_6208;
wire n_6739;
wire n_15779;
wire n_8202;
wire n_15366;
wire n_12734;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_10269;
wire n_19504;
wire n_12262;
wire n_14910;
wire n_14385;
wire n_14499;
wire n_8738;
wire n_9126;
wire n_15368;
wire n_19077;
wire n_11376;
wire n_9438;
wire n_18433;
wire n_7808;
wire n_6544;
wire n_9122;
wire n_14731;
wire n_20227;
wire n_20397;
wire n_16337;
wire n_17691;
wire n_8721;
wire n_12820;
wire n_9912;
wire n_6356;
wire n_13558;
wire n_10148;
wire n_19491;
wire n_16890;
wire n_13890;
wire n_9264;
wire n_14483;
wire n_8326;
wire n_8670;
wire n_15179;
wire n_7638;
wire n_15724;
wire n_19303;
wire n_20412;
wire n_10234;
wire n_8836;
wire n_7019;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_13521;
wire n_19788;
wire n_20611;
wire n_14926;
wire n_10731;
wire n_9878;
wire n_14591;
wire n_14363;
wire n_14576;
wire n_17797;
wire n_11498;
wire n_10513;
wire n_7296;
wire n_7575;
wire n_7083;
wire n_7720;
wire n_11643;
wire n_6268;
wire n_6456;
wire n_11103;
wire n_16823;
wire n_16966;
wire n_14088;
wire n_17926;
wire n_13817;
wire n_9971;
wire n_19579;
wire n_10894;
wire n_14118;
wire n_18082;
wire n_9524;
wire n_20534;
wire n_9243;
wire n_6467;
wire n_9282;
wire n_6796;
wire n_19821;
wire n_18821;
wire n_12417;
wire n_13225;
wire n_20045;
wire n_17006;
wire n_10208;
wire n_20107;
wire n_10804;
wire n_6486;
wire n_17246;
wire n_17167;
wire n_20513;
wire n_18357;
wire n_8438;
wire n_13355;
wire n_18160;
wire n_18614;
wire n_20475;
wire n_10793;
wire n_14672;
wire n_15127;
wire n_6732;
wire n_12711;
wire n_20454;
wire n_12219;
wire n_10440;
wire n_9695;
wire n_11306;
wire n_19169;
wire n_19813;
wire n_8757;
wire n_13035;
wire n_7020;
wire n_13021;
wire n_12893;
wire n_8596;
wire n_11292;
wire n_20238;
wire n_13502;
wire n_6298;
wire n_12289;
wire n_10813;
wire n_10757;
wire n_13046;
wire n_13935;
wire n_16670;
wire n_11431;
wire n_13646;
wire n_18186;
wire n_6197;
wire n_6658;
wire n_8834;
wire n_16429;
wire n_15262;
wire n_10822;
wire n_18773;
wire n_7104;
wire n_7467;
wire n_14609;
wire n_9534;
wire n_13380;
wire n_17369;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_11836;
wire n_6602;
wire n_10924;
wire n_17421;
wire n_11186;
wire n_9742;
wire n_6484;
wire n_19642;
wire n_12527;
wire n_19800;
wire n_9019;
wire n_13891;
wire n_8985;
wire n_7692;
wire n_19463;
wire n_12477;
wire n_14325;
wire n_15503;
wire n_10418;
wire n_19589;
wire n_10875;
wire n_11736;
wire n_7560;
wire n_16270;
wire n_14729;
wire n_11846;
wire n_12400;
wire n_16861;
wire n_9145;
wire n_12092;
wire n_12295;
wire n_9754;
wire n_19549;
wire n_9315;
wire n_18483;
wire n_7451;
wire n_6734;
wire n_7476;
wire n_18096;
wire n_7495;
wire n_7392;
wire n_9765;
wire n_6941;
wire n_7829;
wire n_8680;
wire n_20461;
wire n_16522;
wire n_20246;
wire n_10394;
wire n_11391;
wire n_15462;
wire n_20328;
wire n_12714;
wire n_16779;
wire n_19024;
wire n_9763;
wire n_11070;
wire n_13337;
wire n_15112;
wire n_18146;
wire n_9162;
wire n_19977;
wire n_14849;
wire n_16661;
wire n_11648;
wire n_19044;
wire n_10322;
wire n_7135;
wire n_8555;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_15912;
wire n_16206;
wire n_19812;
wire n_8508;
wire n_19509;
wire n_18827;
wire n_16529;
wire n_8207;
wire n_11653;
wire n_20033;
wire n_11717;
wire n_15246;
wire n_14940;
wire n_6165;
wire n_19153;
wire n_17553;
wire n_15395;
wire n_12838;
wire n_19918;
wire n_18813;
wire n_13505;
wire n_12776;
wire n_19962;
wire n_7033;
wire n_13156;
wire n_15529;
wire n_10710;
wire n_8850;
wire n_14647;
wire n_18384;
wire n_8002;
wire n_19610;
wire n_16722;
wire n_9090;
wire n_16412;
wire n_12008;
wire n_6119;
wire n_9261;
wire n_8301;
wire n_17453;
wire n_12223;
wire n_18706;
wire n_16758;
wire n_10942;
wire n_19983;
wire n_11430;
wire n_13010;
wire n_19073;
wire n_11239;
wire n_10953;
wire n_7842;
wire n_6202;
wire n_17831;
wire n_12898;
wire n_19523;
wire n_15540;
wire n_10343;
wire n_9258;
wire n_10286;
wire n_10371;
wire n_14990;
wire n_16691;
wire n_7236;
wire n_10257;
wire n_11219;
wire n_20232;
wire n_10047;
wire n_14541;
wire n_20609;
wire n_16186;
wire n_13766;
wire n_11226;
wire n_16989;
wire n_11413;
wire n_16617;
wire n_13710;
wire n_11232;
wire n_9105;
wire n_12080;
wire n_16261;
wire n_19512;
wire n_9668;
wire n_13335;
wire n_14022;
wire n_11276;
wire n_10744;
wire n_9870;
wire n_11334;
wire n_7678;
wire n_13075;
wire n_13736;
wire n_13129;
wire n_9178;
wire n_16118;
wire n_6504;
wire n_13586;
wire n_15813;
wire n_10597;
wire n_17382;
wire n_16281;
wire n_11827;
wire n_13049;
wire n_13961;
wire n_17413;
wire n_15745;
wire n_20400;
wire n_6684;
wire n_19084;
wire n_13063;
wire n_20057;
wire n_9323;
wire n_19728;
wire n_6961;
wire n_13252;
wire n_9922;
wire n_12024;
wire n_13084;
wire n_16622;
wire n_15374;
wire n_18123;
wire n_16440;
wire n_7929;
wire n_16821;
wire n_10572;
wire n_16431;
wire n_19272;
wire n_19455;
wire n_13985;
wire n_17594;
wire n_20411;
wire n_14124;
wire n_19119;
wire n_17658;
wire n_13552;
wire n_18086;
wire n_12681;
wire n_18419;
wire n_13022;
wire n_18583;
wire n_17047;
wire n_9513;
wire n_16447;
wire n_16124;
wire n_15446;
wire n_10555;
wire n_19179;
wire n_10314;
wire n_6988;
wire n_13656;
wire n_18967;
wire n_20585;
wire n_6834;
wire n_6817;
wire n_6927;
wire n_20017;
wire n_16841;
wire n_15470;
wire n_6215;
wire n_20316;
wire n_15754;
wire n_17375;
wire n_7862;
wire n_16708;
wire n_17439;
wire n_10630;
wire n_17955;
wire n_8808;
wire n_10061;
wire n_15599;
wire n_11865;
wire n_13024;
wire n_10694;
wire n_20499;
wire n_11041;
wire n_14490;
wire n_9708;
wire n_15479;
wire n_7119;
wire n_8889;
wire n_13986;
wire n_9790;
wire n_11973;
wire n_13329;
wire n_7874;
wire n_8490;
wire n_10329;
wire n_9979;
wire n_8767;
wire n_13946;
wire n_9505;
wire n_15028;
wire n_7102;
wire n_7420;
wire n_13618;
wire n_19838;
wire n_10662;
wire n_18653;
wire n_17534;
wire n_14993;
wire n_14327;
wire n_8624;
wire n_11022;
wire n_10247;
wire n_8796;
wire n_17829;
wire n_10733;
wire n_10472;
wire n_12597;
wire n_13744;
wire n_12834;
wire n_10066;
wire n_17239;
wire n_14335;
wire n_6419;
wire n_18989;
wire n_15087;
wire n_6244;
wire n_6900;
wire n_9337;
wire n_15219;
wire n_9432;
wire n_17295;
wire n_19563;
wire n_7705;
wire n_18331;
wire n_7932;
wire n_7058;
wire n_15009;
wire n_8262;
wire n_9874;
wire n_7981;
wire n_12588;
wire n_17203;
wire n_15648;
wire n_17548;
wire n_9231;
wire n_20230;
wire n_18612;
wire n_7973;
wire n_6815;
wire n_15634;
wire n_9569;
wire n_14823;
wire n_19938;
wire n_14691;
wire n_16908;
wire n_16508;
wire n_9719;
wire n_8358;
wire n_9552;
wire n_13822;
wire n_14948;
wire n_6317;
wire n_10756;
wire n_20333;
wire n_17099;
wire n_14387;
wire n_16572;
wire n_11797;
wire n_18889;
wire n_18933;
wire n_14106;
wire n_18788;
wire n_13616;
wire n_18667;
wire n_7820;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_15468;
wire n_9633;
wire n_13627;
wire n_19040;
wire n_13112;
wire n_10042;
wire n_10478;
wire n_16581;
wire n_18597;
wire n_13163;
wire n_8754;
wire n_9847;
wire n_16968;
wire n_18098;
wire n_10367;
wire n_10867;
wire n_7460;
wire n_9519;
wire n_19735;
wire n_14814;
wire n_6367;
wire n_13564;
wire n_12671;
wire n_8714;
wire n_13260;
wire n_17302;
wire n_10085;
wire n_20023;
wire n_8182;
wire n_16165;
wire n_14090;
wire n_7200;
wire n_15424;
wire n_17301;
wire n_15554;
wire n_15836;
wire n_15966;
wire n_16009;
wire n_15309;
wire n_14463;
wire n_13503;
wire n_11152;
wire n_16318;
wire n_20182;
wire n_14166;
wire n_10122;
wire n_9327;
wire n_16175;
wire n_14271;
wire n_7059;
wire n_14425;
wire n_6327;
wire n_11964;
wire n_7826;
wire n_19078;
wire n_7076;
wire n_11403;
wire n_6866;
wire n_17108;
wire n_9387;
wire n_14596;
wire n_6514;
wire n_9794;
wire n_20571;
wire n_16387;
wire n_11142;
wire n_20147;
wire n_17434;
wire n_17509;
wire n_20261;
wire n_10862;
wire n_8911;
wire n_8248;
wire n_11476;
wire n_13633;
wire n_14538;
wire n_19534;
wire n_17999;
wire n_11367;
wire n_15478;
wire n_16797;
wire n_12676;
wire n_20432;
wire n_18755;
wire n_13913;
wire n_19166;
wire n_8733;
wire n_7976;
wire n_13080;
wire n_13403;
wire n_17444;
wire n_14952;
wire n_10386;
wire n_12128;
wire n_14060;
wire n_14018;
wire n_15959;
wire n_11026;
wire n_13309;
wire n_15292;
wire n_11467;
wire n_12672;
wire n_12063;
wire n_8330;
wire n_15560;
wire n_15065;
wire n_9696;
wire n_20220;
wire n_15771;
wire n_15508;
wire n_20555;
wire n_17990;
wire n_14148;
wire n_12924;
wire n_16331;
wire n_12732;
wire n_17171;
wire n_12649;
wire n_17458;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_6649;
wire n_6283;
wire n_12843;
wire n_14279;
wire n_17856;
wire n_19573;
wire n_15687;
wire n_8540;
wire n_11248;
wire n_9915;
wire n_6089;
wire n_7588;
wire n_18480;
wire n_10017;
wire n_20540;
wire n_11141;
wire n_11093;
wire n_19556;
wire n_17716;
wire n_19873;
wire n_6713;
wire n_18750;
wire n_15968;
wire n_17893;
wire n_13181;
wire n_18303;
wire n_16487;
wire n_17592;
wire n_15047;
wire n_8343;
wire n_7593;
wire n_17156;
wire n_17908;
wire n_14085;
wire n_8068;
wire n_19599;
wire n_7764;
wire n_20357;
wire n_19634;
wire n_10196;
wire n_14573;
wire n_17433;
wire n_19453;
wire n_20085;
wire n_8693;
wire n_6454;
wire n_12625;
wire n_12177;
wire n_7307;
wire n_14512;
wire n_6918;
wire n_16214;
wire n_13761;
wire n_19576;
wire n_19065;
wire n_16219;
wire n_17017;
wire n_14456;
wire n_13364;
wire n_11494;
wire n_14743;
wire n_10218;
wire n_18492;
wire n_19127;
wire n_14859;
wire n_8062;
wire n_11832;
wire n_6375;
wire n_12974;
wire n_13078;
wire n_7047;
wire n_6632;
wire n_17241;
wire n_15795;
wire n_10542;
wire n_16814;
wire n_10681;
wire n_15162;
wire n_9732;
wire n_16494;
wire n_13370;
wire n_11894;
wire n_10222;
wire n_10524;
wire n_6705;
wire n_17988;
wire n_8629;
wire n_9517;
wire n_15237;
wire n_15862;
wire n_6591;
wire n_13643;
wire n_9780;
wire n_13607;
wire n_6289;
wire n_8524;
wire n_19355;
wire n_18907;
wire n_14114;
wire n_14904;
wire n_6512;
wire n_13820;
wire n_6703;
wire n_12122;
wire n_13428;
wire n_17958;
wire n_19667;
wire n_17194;
wire n_19686;
wire n_6086;
wire n_20483;
wire n_16668;
wire n_18139;
wire n_12184;
wire n_10210;
wire n_12571;
wire n_6219;
wire n_11853;
wire n_19626;
wire n_16770;
wire n_9609;
wire n_10029;
wire n_6761;
wire n_8972;
wire n_19919;
wire n_11725;
wire n_13635;
wire n_10801;
wire n_9206;
wire n_18488;
wire n_15698;
wire n_6811;
wire n_16865;
wire n_18642;
wire n_11622;
wire n_12336;
wire n_18345;
wire n_19754;
wire n_12543;
wire n_16129;
wire n_9705;
wire n_16585;
wire n_17490;
wire n_9624;
wire n_20306;
wire n_10389;
wire n_15688;
wire n_13677;
wire n_13757;
wire n_14036;
wire n_12463;
wire n_10990;
wire n_11640;
wire n_12263;
wire n_8982;
wire n_17899;
wire n_13910;
wire n_7086;
wire n_9532;
wire n_18195;
wire n_6601;
wire n_16247;
wire n_13196;
wire n_17482;
wire n_19261;
wire n_8034;
wire n_15824;
wire n_9836;
wire n_11525;
wire n_11999;
wire n_10837;
wire n_18921;
wire n_20299;
wire n_10554;
wire n_8994;
wire n_17827;
wire n_8413;
wire n_19986;
wire n_10149;
wire n_19473;
wire n_19393;
wire n_20020;
wire n_15791;
wire n_12190;
wire n_15484;
wire n_15152;
wire n_19961;
wire n_11847;
wire n_11976;
wire n_20346;
wire n_12511;
wire n_11167;
wire n_8765;
wire n_8213;
wire n_14472;
wire n_10534;
wire n_11049;
wire n_14974;
wire n_8451;
wire n_19410;
wire n_12743;
wire n_16523;
wire n_8731;
wire n_8385;
wire n_15587;
wire n_7370;
wire n_15322;
wire n_13539;
wire n_9350;
wire n_18324;
wire n_19383;
wire n_17917;
wire n_7026;
wire n_7053;
wire n_14618;
wire n_9226;
wire n_18810;
wire n_10608;
wire n_16355;
wire n_7173;
wire n_7042;
wire n_17314;
wire n_17915;
wire n_19225;
wire n_19011;
wire n_16774;
wire n_16436;
wire n_10638;
wire n_17923;
wire n_9112;
wire n_18582;
wire n_18970;
wire n_19284;
wire n_9235;
wire n_16570;
wire n_19124;
wire n_13852;
wire n_9333;
wire n_17813;
wire n_14089;
wire n_20641;
wire n_15758;
wire n_11804;
wire n_14234;
wire n_14125;
wire n_6562;
wire n_12809;
wire n_18770;
wire n_11052;
wire n_17350;
wire n_18598;
wire n_6671;
wire n_13470;
wire n_6812;
wire n_12361;
wire n_19151;
wire n_9488;
wire n_10748;
wire n_13068;
wire n_19158;
wire n_18795;
wire n_20459;
wire n_7792;
wire n_15985;
wire n_8161;
wire n_18798;
wire n_10014;
wire n_15723;
wire n_16840;
wire n_18698;
wire n_10677;
wire n_18269;
wire n_15852;
wire n_18857;
wire n_19216;
wire n_12321;
wire n_11247;
wire n_18581;
wire n_8384;
wire n_6445;
wire n_18079;
wire n_13106;
wire n_19863;
wire n_14294;
wire n_17609;
wire n_6701;
wire n_14862;
wire n_7380;
wire n_8736;
wire n_11514;
wire n_12470;
wire n_18604;
wire n_12994;
wire n_10215;
wire n_20005;
wire n_18768;
wire n_14059;
wire n_10834;
wire n_17632;
wire n_20257;
wire n_17611;
wire n_19341;
wire n_12064;
wire n_12696;
wire n_18024;
wire n_15735;
wire n_11133;
wire n_20054;
wire n_17143;
wire n_18341;
wire n_10871;
wire n_16405;
wire n_14624;
wire n_16600;
wire n_15036;
wire n_17695;
wire n_18193;
wire n_19489;
wire n_11571;
wire n_14120;
wire n_8844;
wire n_13147;
wire n_7641;
wire n_6106;
wire n_14407;
wire n_14260;
wire n_16845;
wire n_18924;
wire n_17307;
wire n_7169;
wire n_10407;
wire n_19330;
wire n_14175;
wire n_11941;
wire n_15780;
wire n_18085;
wire n_15189;
wire n_8110;
wire n_9008;
wire n_12079;
wire n_15335;
wire n_19147;
wire n_15227;
wire n_8805;
wire n_7209;
wire n_18908;
wire n_15026;
wire n_13895;
wire n_6979;
wire n_13222;
wire n_17284;
wire n_15987;
wire n_10462;
wire n_20440;
wire n_11769;
wire n_8856;
wire n_19362;
wire n_6142;
wire n_20582;
wire n_14901;
wire n_7769;
wire n_17034;
wire n_10291;
wire n_18575;
wire n_18764;
wire n_17502;
wire n_14333;
wire n_7233;
wire n_8732;
wire n_13506;
wire n_7602;
wire n_9296;
wire n_18587;
wire n_7390;
wire n_10669;
wire n_19515;
wire n_8231;
wire n_20161;
wire n_13717;
wire n_7598;
wire n_12440;
wire n_19032;
wire n_8908;
wire n_16085;
wire n_6767;
wire n_12782;
wire n_10111;
wire n_19186;
wire n_19629;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_20009;
wire n_17796;
wire n_7045;
wire n_8740;
wire n_11727;
wire n_6788;
wire n_12192;
wire n_17342;
wire n_14465;
wire n_13412;
wire n_11749;
wire n_11300;
wire n_6143;
wire n_20569;
wire n_13457;
wire n_12551;
wire n_18066;
wire n_12497;
wire n_15043;
wire n_16602;
wire n_16864;
wire n_16761;
wire n_7679;
wire n_20593;
wire n_18133;
wire n_20529;
wire n_7936;
wire n_8966;
wire n_10287;
wire n_8538;
wire n_12101;
wire n_11145;
wire n_16684;
wire n_19594;
wire n_10349;
wire n_16340;
wire n_7490;
wire n_7545;
wire n_7160;
wire n_9809;
wire n_10750;
wire n_7295;
wire n_14338;
wire n_7348;
wire n_19071;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_17554;
wire n_16071;
wire n_15394;
wire n_16875;
wire n_15941;
wire n_20439;
wire n_9558;
wire n_11594;
wire n_8715;
wire n_12474;
wire n_7162;
wire n_16655;
wire n_20272;
wire n_12346;
wire n_18167;
wire n_8371;
wire n_13916;
wire n_15195;
wire n_11458;
wire n_17056;
wire n_12244;
wire n_18753;
wire n_16188;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_7681;
wire n_11504;
wire n_19972;
wire n_16850;
wire n_13981;
wire n_11516;
wire n_8392;
wire n_14659;
wire n_8095;
wire n_10830;
wire n_16868;
wire n_17644;
wire n_7503;
wire n_6854;
wire n_17254;
wire n_18733;
wire n_12953;
wire n_15224;
wire n_9215;
wire n_11406;
wire n_19835;
wire n_11047;
wire n_14963;
wire n_8050;
wire n_12817;
wire n_8399;
wire n_16916;
wire n_13866;
wire n_12435;
wire n_10946;
wire n_18106;
wire n_7065;
wire n_9216;
wire n_11961;
wire n_6122;
wire n_7911;
wire n_17486;
wire n_17504;
wire n_7330;
wire n_14605;
wire n_9202;
wire n_13543;
wire n_10351;
wire n_13772;
wire n_7493;
wire n_12940;
wire n_10460;
wire n_15487;
wire n_19221;
wire n_10334;
wire n_11614;
wire n_15242;
wire n_8422;
wire n_12224;
wire n_7088;
wire n_9394;
wire n_8878;
wire n_7440;
wire n_17681;
wire n_17676;
wire n_14797;
wire n_9622;
wire n_14177;
wire n_14093;
wire n_14607;
wire n_10191;
wire n_17919;
wire n_12679;
wire n_11168;
wire n_14921;
wire n_20406;
wire n_10911;
wire n_12756;
wire n_16097;
wire n_9845;
wire n_16147;
wire n_7374;
wire n_14389;
wire n_19514;
wire n_11937;
wire n_17277;
wire n_8251;
wire n_14621;
wire n_18864;
wire n_20468;
wire n_17875;
wire n_11192;
wire n_6852;
wire n_8677;
wire n_9091;
wire n_17206;
wire n_13914;
wire n_14663;
wire n_16921;
wire n_17559;
wire n_9699;
wire n_13277;
wire n_12340;
wire n_18143;
wire n_16742;
wire n_18464;
wire n_13494;
wire n_9751;
wire n_20525;
wire n_10543;
wire n_7924;
wire n_17225;
wire n_20443;
wire n_7659;
wire n_20539;
wire n_16203;
wire n_8875;
wire n_20079;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_12662;
wire n_15697;
wire n_17879;
wire n_18140;
wire n_9293;
wire n_12503;
wire n_18510;
wire n_15202;
wire n_18218;
wire n_12871;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_18224;
wire n_16400;
wire n_20441;
wire n_10809;
wire n_16934;
wire n_10899;
wire n_9639;
wire n_11898;
wire n_15250;
wire n_17193;
wire n_6711;
wire n_11997;
wire n_8946;
wire n_13090;
wire n_18984;
wire n_13541;
wire n_20092;
wire n_16958;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_17396;
wire n_7275;
wire n_8795;
wire n_7195;
wire n_11199;
wire n_17642;
wire n_11264;
wire n_19791;
wire n_7610;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_16229;
wire n_10006;
wire n_11757;
wire n_18447;
wire n_12622;
wire n_6353;
wire n_12659;
wire n_6818;
wire n_7539;
wire n_12629;
wire n_12868;
wire n_19263;
wire n_10275;
wire n_7775;
wire n_11392;
wire n_7930;
wire n_7661;
wire n_16498;
wire n_19673;
wire n_14165;
wire n_17309;
wire n_19413;
wire n_13787;
wire n_13674;
wire n_18311;
wire n_13912;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_11278;
wire n_14445;
wire n_7548;
wire n_16732;
wire n_6156;
wire n_12913;
wire n_7064;
wire n_19285;
wire n_16839;
wire n_16798;
wire n_12154;
wire n_8000;
wire n_14427;
wire n_18327;
wire n_6917;
wire n_6937;
wire n_20527;
wire n_9963;
wire n_17211;
wire n_20337;
wire n_7324;
wire n_10152;
wire n_17568;
wire n_6301;
wire n_18061;
wire n_16815;
wire n_18022;
wire n_15570;
wire n_15562;
wire n_17207;
wire n_19000;
wire n_7729;
wire n_19622;
wire n_6436;
wire n_16987;
wire n_18337;
wire n_20320;
wire n_6699;
wire n_12926;
wire n_14809;
wire n_14725;
wire n_16892;
wire n_19717;
wire n_6874;
wire n_6259;
wire n_9340;
wire n_16527;
wire n_17963;
wire n_6677;
wire n_12161;
wire n_11735;
wire n_20450;
wire n_8769;
wire n_6764;
wire n_10324;
wire n_11189;
wire n_8815;
wire n_12044;
wire n_9303;
wire n_8261;
wire n_13104;
wire n_19730;
wire n_7139;
wire n_16819;
wire n_16612;
wire n_20309;
wire n_9722;
wire n_12155;
wire n_15664;
wire n_12373;
wire n_19376;
wire n_14579;
wire n_17930;
wire n_8665;
wire n_15847;
wire n_7751;
wire n_18763;
wire n_20352;
wire n_14718;
wire n_19253;
wire n_18298;
wire n_13116;
wire n_19781;
wire n_14589;
wire n_12386;
wire n_14257;
wire n_16492;
wire n_16811;
wire n_8835;
wire n_18645;
wire n_20354;
wire n_10688;
wire n_16771;
wire n_12964;
wire n_20069;
wire n_16404;
wire n_15099;
wire n_20144;
wire n_7579;
wire n_16874;
wire n_11687;
wire n_20157;
wire n_8870;
wire n_7155;
wire n_6475;
wire n_7699;
wire n_15951;
wire n_6103;
wire n_8781;
wire n_6394;
wire n_18618;
wire n_14102;
wire n_20438;
wire n_17196;
wire n_12267;
wire n_15803;
wire n_8365;
wire n_13780;
wire n_16699;
wire n_19844;
wire n_7194;
wire n_6752;
wire n_6426;
wire n_8025;
wire n_8502;
wire n_7612;
wire n_20628;
wire n_16999;
wire n_18843;
wire n_11120;
wire n_6350;
wire n_19702;
wire n_7736;
wire n_16040;
wire n_14259;
wire n_20030;
wire n_6159;
wire n_13360;
wire n_8479;
wire n_14214;
wire n_15558;
wire n_17306;
wire n_6235;
wire n_17996;
wire n_12647;
wire n_7662;
wire n_15340;
wire n_16061;
wire n_7773;
wire n_16776;
wire n_13048;
wire n_13563;
wire n_17905;
wire n_7555;
wire n_19764;
wire n_12060;
wire n_18254;
wire n_10199;
wire n_8658;
wire n_11910;
wire n_15377;
wire n_15583;
wire n_13347;
wire n_8866;
wire n_8061;
wire n_16623;
wire n_17186;
wire n_13111;
wire n_15563;
wire n_10117;
wire n_12716;
wire n_16341;
wire n_16679;
wire n_13456;
wire n_10198;
wire n_7157;
wire n_13237;
wire n_15448;
wire n_7411;
wire n_19716;
wire n_16851;
wire n_7871;
wire n_12051;
wire n_6477;
wire n_15298;
wire n_11533;
wire n_8652;
wire n_7198;
wire n_9904;
wire n_17891;
wire n_19182;
wire n_6184;
wire n_10973;
wire n_11036;
wire n_17362;
wire n_10267;
wire n_10551;
wire n_18589;
wire n_17029;
wire n_17924;
wire n_18323;
wire n_13127;
wire n_18004;
wire n_11002;
wire n_19637;
wire n_14075;
wire n_9032;
wire n_6313;
wire n_18884;
wire n_16184;
wire n_7145;
wire n_12325;
wire n_9245;
wire n_9357;
wire n_19060;
wire n_15766;
wire n_18121;
wire n_16759;
wire n_14530;
wire n_17724;
wire n_19773;
wire n_7994;
wire n_14206;
wire n_17328;
wire n_7349;
wire n_9598;
wire n_14481;
wire n_17993;
wire n_15044;
wire n_12504;
wire n_12602;
wire n_12062;
wire n_15375;
wire n_16100;
wire n_12335;
wire n_12949;
wire n_13611;
wire n_15268;
wire n_10487;
wire n_10960;
wire n_6141;
wire n_18540;
wire n_20409;
wire n_10931;
wire n_19831;
wire n_11574;
wire n_15049;
wire n_15181;
wire n_8168;
wire n_7190;
wire n_14870;
wire n_12322;
wire n_14196;
wire n_10236;
wire n_11205;
wire n_11776;
wire n_20169;
wire n_11650;
wire n_19197;
wire n_12179;
wire n_14439;
wire n_20229;
wire n_9896;
wire n_11856;
wire n_14825;
wire n_20631;
wire n_11536;
wire n_14914;
wire n_10283;
wire n_19865;
wire n_6324;
wire n_13437;
wire n_15623;
wire n_16696;
wire n_20516;
wire n_18865;
wire n_8411;
wire n_16733;
wire n_18799;
wire n_13221;
wire n_11163;
wire n_13657;
wire n_14099;
wire n_15632;
wire n_16245;
wire n_11419;
wire n_12095;
wire n_9018;
wire n_13990;
wire n_16302;
wire n_13663;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_14939;
wire n_11740;
wire n_17471;
wire n_8444;
wire n_20369;
wire n_17227;
wire n_7008;
wire n_12392;
wire n_11979;
wire n_7596;
wire n_20579;
wire n_6280;
wire n_18090;
wire n_18626;
wire n_10759;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_19960;
wire n_18211;
wire n_8977;
wire n_20025;
wire n_15797;
wire n_9962;
wire n_11104;
wire n_11537;
wire n_13814;
wire n_18993;
wire n_12707;
wire n_14861;
wire n_7686;
wire n_15194;
wire n_18894;
wire n_15572;
wire n_12424;
wire n_11699;
wire n_8125;
wire n_14811;
wire n_17608;
wire n_10226;
wire n_6526;
wire n_17401;
wire n_7196;
wire n_14864;
wire n_17936;
wire n_16643;
wire n_12107;
wire n_10161;
wire n_9842;
wire n_9614;
wire n_16024;
wire n_10699;
wire n_7846;
wire n_8598;
wire n_7256;
wire n_16078;
wire n_7331;
wire n_13509;
wire n_17637;
wire n_7342;
wire n_14791;
wire n_14485;
wire n_10606;
wire n_11164;
wire n_12203;
wire n_7147;
wire n_12359;
wire n_19175;
wire n_9037;
wire n_15983;
wire n_12548;
wire n_15874;
wire n_14461;
wire n_20600;
wire n_13958;
wire n_17619;
wire n_6863;
wire n_10012;
wire n_13754;
wire n_12985;
wire n_20087;
wire n_16191;
wire n_14171;
wire n_6768;
wire n_15212;
wire n_15977;
wire n_9128;
wire n_9872;
wire n_14380;
wire n_10310;
wire n_15896;
wire n_6151;
wire n_16843;
wire n_7110;
wire n_17273;
wire n_13920;
wire n_18119;
wire n_10097;
wire n_8915;
wire n_16509;
wire n_9866;
wire n_9858;
wire n_13977;
wire n_8727;
wire n_18494;
wire n_16538;
wire n_11662;
wire n_16992;
wire n_18065;
wire n_10266;
wire n_17949;
wire n_20099;
wire n_7734;
wire n_8955;
wire n_20001;
wire n_17781;
wire n_12384;
wire n_15438;
wire n_11260;
wire n_11351;
wire n_15611;
wire n_14388;
wire n_12249;
wire n_14977;
wire n_10628;
wire n_13429;
wire n_7905;
wire n_11775;
wire n_10769;
wire n_10256;
wire n_13999;
wire n_14037;
wire n_11706;
wire n_11800;
wire n_18382;
wire n_11642;
wire n_20235;
wire n_11143;
wire n_17103;
wire n_11074;
wire n_6831;
wire n_16352;
wire n_18713;
wire n_18032;
wire n_11934;
wire n_7677;
wire n_10396;
wire n_13919;
wire n_19357;
wire n_13642;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_10693;
wire n_15872;
wire n_13240;
wire n_20336;
wire n_12578;
wire n_12194;
wire n_7519;
wire n_7400;
wire n_15649;
wire n_9724;
wire n_9281;
wire n_10101;
wire n_15863;
wire n_6581;
wire n_19690;
wire n_7013;
wire n_14150;
wire n_12125;
wire n_7290;
wire n_18830;
wire n_9687;
wire n_18052;
wire n_19108;
wire n_9426;
wire n_7889;
wire n_9102;
wire n_11526;
wire n_16115;
wire n_14128;
wire n_11851;
wire n_18983;
wire n_17323;
wire n_6965;
wire n_9144;
wire n_18191;
wire n_7461;
wire n_15133;
wire n_16885;
wire n_9521;
wire n_15288;
wire n_16900;
wire n_13040;
wire n_7278;
wire n_6509;
wire n_7454;
wire n_11253;
wire n_17102;
wire n_15527;
wire n_12861;
wire n_17443;
wire n_16146;
wire n_16654;
wire n_12918;
wire n_18332;
wire n_18145;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_16991;
wire n_18051;
wire n_19051;
wire n_13716;
wire n_7069;
wire n_7904;
wire n_11691;
wire n_14408;
wire n_9410;
wire n_12865;
wire n_10712;
wire n_7168;
wire n_17604;
wire n_18765;
wire n_7970;
wire n_7091;
wire n_10972;
wire n_6359;
wire n_20564;
wire n_10945;
wire n_8800;
wire n_10845;
wire n_8229;
wire n_18743;
wire n_14863;
wire n_6766;
wire n_7629;
wire n_9735;
wire n_18831;
wire n_20344;
wire n_20541;
wire n_14711;
wire n_9802;
wire n_14373;
wire n_8107;
wire n_11108;
wire n_12992;
wire n_11004;
wire n_6519;
wire n_15752;
wire n_11686;
wire n_6530;
wire n_10566;
wire n_17798;
wire n_19592;
wire n_16568;
wire n_17581;
wire n_18906;
wire n_12104;
wire n_17954;
wire n_6402;
wire n_12469;
wire n_19554;
wire n_15829;
wire n_19568;
wire n_7326;
wire n_17522;
wire n_7067;
wire n_14835;
wire n_15391;
wire n_16226;
wire n_14871;
wire n_8691;
wire n_14907;
wire n_6748;
wire n_11719;
wire n_19307;
wire n_16685;
wire n_19498;
wire n_16979;
wire n_18282;
wire n_15358;
wire n_14636;
wire n_8026;
wire n_7528;
wire n_9638;
wire n_16069;
wire n_20101;
wire n_8174;
wire n_13524;
wire n_11175;
wire n_10040;
wire n_8861;
wire n_8644;
wire n_12304;
wire n_15156;
wire n_13138;
wire n_7117;
wire n_18490;
wire n_6205;
wire n_20141;
wire n_7136;
wire n_6754;
wire n_12692;
wire n_7939;
wire n_13602;
wire n_17436;
wire n_16785;
wire n_9612;
wire n_10790;
wire n_14919;
wire n_16653;
wire n_9108;
wire n_6723;
wire n_16692;
wire n_7436;
wire n_6440;
wire n_14101;
wire n_9376;
wire n_8446;
wire n_17654;
wire n_20396;
wire n_12996;
wire n_15171;
wire n_19711;
wire n_13625;
wire n_12643;
wire n_6124;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_19265;
wire n_8197;
wire n_6622;
wire n_11521;
wire n_20463;
wire n_12827;
wire n_12678;
wire n_15868;
wire n_17249;
wire n_7747;
wire n_9779;
wire n_8082;
wire n_8730;
wire n_15533;
wire n_6528;
wire n_15165;
wire n_13475;
wire n_15079;
wire n_19822;
wire n_13859;
wire n_18640;
wire n_12713;
wire n_13144;
wire n_18129;
wire n_19488;
wire n_10660;
wire n_7430;
wire n_18560;
wire n_9937;
wire n_7912;
wire n_16749;
wire n_8281;
wire n_20347;
wire n_19437;
wire n_18876;
wire n_20174;
wire n_19430;
wire n_11428;
wire n_17626;
wire n_11677;
wire n_7281;
wire n_9717;
wire n_13577;
wire n_18523;
wire n_19176;
wire n_19970;
wire n_13769;
wire n_18044;
wire n_13672;
wire n_19036;
wire n_17600;
wire n_8956;
wire n_6763;
wire n_7858;
wire n_20203;
wire n_6542;
wire n_15681;
wire n_17262;
wire n_6556;
wire n_20245;
wire n_12374;
wire n_8998;
wire n_10538;
wire n_13342;
wire n_18856;
wire n_9123;
wire n_17374;
wire n_6471;
wire n_15545;
wire n_14924;
wire n_11867;
wire n_12796;
wire n_16053;
wire n_19185;
wire n_15708;
wire n_19441;
wire n_11716;
wire n_8979;
wire n_7245;
wire n_18858;
wire n_6675;
wire n_6270;
wire n_18111;
wire n_6808;
wire n_16091;
wire n_20326;
wire n_11886;
wire n_7006;
wire n_16264;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_17231;
wire n_10925;
wire n_20190;
wire n_11158;
wire n_9861;
wire n_15878;
wire n_14390;
wire n_18678;
wire n_8264;
wire n_7381;
wire n_16160;
wire n_12078;
wire n_15647;
wire n_9832;
wire n_19925;
wire n_20547;
wire n_6580;
wire n_18790;
wire n_9898;
wire n_6412;
wire n_18410;
wire n_19959;
wire n_13293;
wire n_6437;
wire n_14381;
wire n_15709;
wire n_18590;
wire n_8408;
wire n_10661;
wire n_9495;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_11771;
wire n_16870;
wire n_19082;
wire n_13833;
wire n_16518;
wire n_9867;
wire n_14441;
wire n_9688;
wire n_10967;
wire n_20620;
wire n_7870;
wire n_18377;
wire n_20208;
wire n_6117;
wire n_11828;
wire n_12326;
wire n_14264;
wire n_19317;
wire n_14115;
wire n_16635;
wire n_8963;
wire n_12309;
wire n_7399;
wire n_13953;
wire n_7482;
wire n_19830;
wire n_14847;
wire n_10312;
wire n_18308;
wire n_9223;
wire n_17465;
wire n_15930;
wire n_13226;
wire n_19416;
wire n_17943;
wire n_16433;
wire n_11244;
wire n_18577;
wire n_14432;
wire n_10209;
wire n_13253;
wire n_8183;
wire n_19936;
wire n_16098;
wire n_11245;
wire n_13354;
wire n_6085;
wire n_12422;
wire n_15616;
wire n_17614;
wire n_14422;
wire n_9694;
wire n_16636;
wire n_9948;
wire n_14630;
wire n_17048;
wire n_18966;
wire n_19390;
wire n_19729;
wire n_10887;
wire n_16876;
wire n_6554;
wire n_12146;
wire n_6560;
wire n_14055;
wire n_12136;
wire n_17046;
wire n_16138;
wire n_12399;
wire n_12342;
wire n_9744;
wire n_7414;
wire n_9548;
wire n_8973;
wire n_6448;
wire n_12378;
wire n_19155;
wire n_12533;
wire n_7431;
wire n_12178;
wire n_18871;
wire n_20192;
wire n_11346;
wire n_17210;
wire n_18206;
wire n_19851;
wire n_14810;
wire n_8249;
wire n_12257;
wire n_15770;
wire n_13394;
wire n_13391;
wire n_14680;
wire n_8234;
wire n_20442;
wire n_16835;
wire n_18438;
wire n_16863;
wire n_9280;
wire n_18285;
wire n_13263;
wire n_14877;
wire n_19815;
wire n_15203;
wire n_11491;
wire n_14048;
wire n_11772;
wire n_16063;
wire n_16237;
wire n_16112;
wire n_15891;
wire n_12769;
wire n_12641;
wire n_10765;
wire n_15263;
wire n_11792;
wire n_20076;
wire n_18776;
wire n_8558;
wire n_10489;
wire n_12421;
wire n_7274;
wire n_10159;
wire n_14351;
wire n_7466;
wire n_13310;
wire n_11568;
wire n_7429;
wire n_11766;
wire n_11038;
wire n_13798;
wire n_16894;
wire n_18890;
wire n_17294;
wire n_16932;
wire n_15842;
wire n_14822;
wire n_8813;
wire n_10356;
wire n_17461;
wire n_18216;
wire n_10173;
wire n_20010;
wire n_19162;
wire n_12311;
wire n_14374;
wire n_9448;
wire n_6555;
wire n_14815;
wire n_10739;
wire n_8470;
wire n_16480;
wire n_20062;
wire n_17657;
wire n_14831;
wire n_11170;
wire n_17683;
wire n_11758;
wire n_9396;
wire n_19486;
wire n_14450;
wire n_7061;
wire n_12480;
wire n_14192;
wire n_9053;
wire n_15504;
wire n_11893;
wire n_10573;
wire n_10850;
wire n_9185;
wire n_19697;
wire n_13376;
wire n_8092;
wire n_13864;
wire n_15279;
wire n_11456;
wire n_10546;
wire n_6574;
wire n_20270;
wire n_6571;
wire n_17484;
wire n_9151;
wire n_7824;
wire n_17202;
wire n_18080;
wire n_20444;
wire n_13236;
wire n_14299;
wire n_7094;
wire n_16320;
wire n_7036;
wire n_13777;
wire n_19359;
wire n_20467;
wire n_6260;
wire n_7413;
wire n_16803;
wire n_17229;
wire n_6286;
wire n_8267;
wire n_18929;
wire n_7175;
wire n_9978;
wire n_11914;
wire n_9670;
wire n_19964;
wire n_9334;
wire n_15131;
wire n_20064;
wire n_12531;
wire n_11302;
wire n_19931;
wire n_19006;
wire n_9413;
wire n_12727;
wire n_20043;
wire n_15509;
wire n_11707;
wire n_7697;
wire n_13835;
wire n_16260;
wire n_7547;
wire n_13815;
wire n_20515;
wire n_9557;
wire n_15957;
wire n_16319;
wire n_17259;
wire n_20355;
wire n_14039;
wire n_6348;
wire n_6744;
wire n_18578;
wire n_8582;
wire n_6293;
wire n_9762;
wire n_8957;
wire n_18646;
wire n_15793;
wire n_6558;
wire n_20323;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_18209;
wire n_9271;
wire n_17747;
wire n_13688;
wire n_11396;
wire n_15196;
wire n_16176;
wire n_20207;
wire n_9483;
wire n_19649;
wire n_19435;
wire n_19769;
wire n_14754;
wire n_19768;
wire n_15020;
wire n_6091;
wire n_14252;
wire n_15830;
wire n_12583;
wire n_7691;
wire n_6551;
wire n_8747;
wire n_9539;
wire n_9385;
wire n_13462;
wire n_9785;
wire n_8922;
wire n_9027;
wire n_12750;
wire n_6995;
wire n_19315;
wire n_9233;
wire n_20544;
wire n_16895;
wire n_10282;
wire n_17602;
wire n_15142;
wire n_10913;
wire n_18803;
wire n_18409;
wire n_17838;
wire n_15991;
wire n_13388;
wire n_13731;
wire n_10703;
wire n_9666;
wire n_14503;
wire n_12248;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_17754;
wire n_14886;
wire n_7993;
wire n_20223;
wire n_7181;
wire n_9865;
wire n_14644;
wire n_11715;
wire n_7071;
wire n_20625;
wire n_15454;
wire n_10642;
wire n_15213;
wire n_18859;
wire n_19946;
wire n_18428;
wire n_12181;
wire n_18670;
wire n_14560;
wire n_17257;
wire n_19726;
wire n_14829;
wire n_11007;
wire n_15473;
wire n_19864;
wire n_15584;
wire n_10316;
wire n_9795;
wire n_18386;
wire n_6429;
wire n_6407;
wire n_16515;
wire n_17914;
wire n_10479;
wire n_13660;
wire n_19280;
wire n_6801;
wire n_18099;
wire n_12738;
wire n_15062;
wire n_20402;
wire n_11599;
wire n_6113;
wire n_10070;
wire n_16178;
wire n_20276;
wire n_18841;
wire n_17304;
wire n_18393;
wire n_14983;
wire n_8439;
wire n_18434;
wire n_9641;
wire n_12755;
wire n_18522;
wire n_12059;
wire n_18541;
wire n_18257;
wire n_15845;
wire n_6129;
wire n_6518;
wire n_20401;
wire n_9138;
wire n_18072;
wire n_18048;
wire n_7537;
wire n_10516;
wire n_8675;
wire n_15924;
wire n_17906;
wire n_12567;
wire n_9367;
wire n_15130;
wire n_11887;
wire n_17852;
wire n_17442;
wire n_10026;
wire n_9729;
wire n_12471;
wire n_12451;
wire n_17243;
wire n_15740;
wire n_20048;
wire n_9411;
wire n_12507;
wire n_14564;
wire n_11277;
wire n_18416;
wire n_20133;
wire n_17606;
wire n_7410;
wire n_8777;
wire n_13581;
wire n_12972;
wire n_13789;
wire n_14511;
wire n_13286;
wire n_9951;
wire n_19023;
wire n_9424;
wire n_10507;
wire n_11968;
wire n_19003;
wire n_10045;
wire n_20179;
wire n_11335;
wire n_20603;
wire n_18606;
wire n_13988;
wire n_15272;
wire n_17169;
wire n_13609;
wire n_16886;
wire n_13679;
wire n_11785;
wire n_10417;
wire n_12841;
wire n_12855;
wire n_17370;
wire n_15834;
wire n_13276;
wire n_8938;
wire n_16058;
wire n_11801;
wire n_16994;
wire n_16519;
wire n_17810;
wire n_14830;
wire n_7867;
wire n_14281;
wire n_14594;
wire n_18213;
wire n_6135;
wire n_17303;
wire n_20263;
wire n_6814;
wire n_10557;
wire n_8669;
wire n_7525;
wire n_19219;
wire n_7257;
wire n_9372;
wire n_6791;
wire n_11915;
wire n_13704;
wire n_11016;
wire n_9326;
wire n_14976;
wire n_7650;
wire n_17297;
wire n_19872;
wire n_13043;
wire n_17260;
wire n_12620;
wire n_12632;
wire n_20198;
wire n_20456;
wire n_6309;
wire n_19618;
wire n_11303;
wire n_6733;
wire n_19047;
wire n_20122;
wire n_9902;
wire n_19910;
wire n_9900;
wire n_17367;
wire n_18937;
wire n_15521;
wire n_18415;
wire n_7202;
wire n_12416;
wire n_8265;
wire n_11609;
wire n_18287;
wire n_16464;
wire n_19597;
wire n_12494;
wire n_10327;
wire n_13826;
wire n_7605;
wire n_11556;
wire n_15140;
wire n_11529;
wire n_10437;
wire n_10021;
wire n_16673;
wire n_9146;
wire n_15753;
wire n_8131;
wire n_8941;
wire n_17093;
wire n_17685;
wire n_16357;
wire n_12623;
wire n_11444;
wire n_6269;
wire n_12213;
wire n_9358;
wire n_6654;
wire n_9565;
wire n_8257;
wire n_13072;
wire n_18120;
wire n_7726;
wire n_17026;
wire n_13839;
wire n_6120;
wire n_13954;
wire n_8799;
wire n_6641;
wire n_19215;
wire n_10124;
wire n_19595;
wire n_14689;
wire n_10245;
wire n_14132;
wire n_10905;
wire n_11235;
wire n_19020;
wire n_6399;
wire n_9563;
wire n_17077;
wire n_17702;
wire n_11166;
wire n_20310;
wire n_7031;
wire n_9285;
wire n_18093;
wire n_16595;
wire n_7763;
wire n_8033;
wire n_15172;
wire n_19470;
wire n_19720;
wire n_8393;
wire n_16561;
wire n_10784;
wire n_8463;
wire n_8153;
wire n_10944;
wire n_10211;
wire n_18554;
wire n_18077;
wire n_12431;
wire n_11855;
wire n_6790;
wire n_17628;
wire n_13799;
wire n_16084;
wire n_13854;
wire n_18250;
wire n_19843;
wire n_15380;
wire n_6686;
wire n_15956;
wire n_18835;
wire n_20035;
wire n_11787;
wire n_16059;
wire n_8103;
wire n_20421;
wire n_14752;
wire n_6183;
wire n_11544;
wire n_15447;
wire n_10730;
wire n_10564;
wire n_8682;
wire n_20307;
wire n_7655;
wire n_18276;
wire n_11509;
wire n_19191;
wire n_11960;
wire n_19905;
wire n_7878;
wire n_9514;
wire n_6210;
wire n_6500;
wire n_12465;
wire n_13532;
wire n_11029;
wire n_13118;
wire n_17390;
wire n_10951;
wire n_12152;
wire n_19415;
wire n_6785;
wire n_10454;
wire n_15401;
wire n_13339;
wire n_8039;
wire n_19323;
wire n_8916;
wire n_10087;
wire n_10146;
wire n_12959;
wire n_9946;
wire n_9885;
wire n_6849;
wire n_20482;
wire n_8162;
wire n_18263;
wire n_7457;
wire n_19982;
wire n_8744;
wire n_10701;
wire n_7752;
wire n_15775;
wire n_17346;
wire n_8286;
wire n_9015;
wire n_20002;
wire n_6452;
wire n_16408;
wire n_20362;
wire n_6611;
wire n_18828;
wire n_18297;
wire n_11433;
wire n_10592;
wire n_18130;
wire n_7207;
wire n_8218;
wire n_17978;
wire n_8537;
wire n_10126;
wire n_14421;
wire n_15890;
wire n_13653;
wire n_12566;
wire n_6227;
wire n_13680;
wire n_16077;
wire n_9066;
wire n_10302;
wire n_12546;
wire n_13058;
wire n_18342;
wire n_12036;
wire n_17650;
wire n_8782;
wire n_12911;
wire n_15715;
wire n_9857;
wire n_12781;
wire n_10057;
wire n_10882;
wire n_9338;
wire n_8144;
wire n_10435;
wire n_9542;
wire n_10921;
wire n_7171;
wire n_12061;
wire n_14585;
wire n_11085;
wire n_16541;
wire n_7068;
wire n_13649;
wire n_10609;
wire n_14804;
wire n_20015;
wire n_9783;
wire n_13806;
wire n_19542;
wire n_9404;
wire n_9916;
wire n_12645;
wire n_18351;
wire n_16198;
wire n_14466;
wire n_7777;
wire n_12138;
wire n_7652;
wire n_10220;
wire n_11347;
wire n_17635;
wire n_10550;
wire n_14673;
wire n_12365;
wire n_20334;
wire n_13738;
wire n_14972;
wire n_16996;
wire n_9306;
wire n_14138;
wire n_10232;
wire n_10461;
wire n_14586;
wire n_7966;
wire n_8591;
wire n_8811;
wire n_19188;
wire n_14031;
wire n_10326;
wire n_8417;
wire n_19978;
wire n_12487;
wire n_7997;
wire n_6420;
wire n_20518;
wire n_12288;
wire n_17300;
wire n_12130;
wire n_13120;
wire n_19825;
wire n_16299;
wire n_12704;
wire n_12271;
wire n_7680;
wire n_15190;
wire n_16909;
wire n_12958;
wire n_8172;
wire n_19848;
wire n_19559;
wire n_9502;
wire n_6447;
wire n_20612;
wire n_19923;
wire n_14761;
wire n_6751;
wire n_15243;
wire n_20090;
wire n_11087;
wire n_11477;
wire n_8375;
wire n_8612;
wire n_8345;
wire n_13725;
wire n_6741;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_19414;
wire n_17551;
wire n_19417;
wire n_9164;
wire n_7183;
wire n_13197;
wire n_10878;
wire n_18408;
wire n_7140;
wire n_20284;
wire n_14860;
wire n_10450;
wire n_19609;
wire n_11472;
wire n_9114;
wire n_11978;
wire n_8515;
wire n_10529;
wire n_14685;
wire n_14892;
wire n_8812;
wire n_14505;
wire n_12254;
wire n_9392;
wire n_14531;
wire n_11538;
wire n_9698;
wire n_13435;
wire n_15408;
wire n_15173;
wire n_9644;
wire n_11353;
wire n_18745;
wire n_9499;
wire n_6647;
wire n_6275;
wire n_14771;
wire n_7750;
wire n_11597;
wire n_15902;
wire n_6277;
wire n_10920;
wire n_14398;
wire n_11126;
wire n_18453;
wire n_9409;
wire n_18629;
wire n_20565;
wire n_17814;
wire n_12555;
wire n_11646;
wire n_9768;
wire n_12980;
wire n_9881;
wire n_6807;
wire n_7251;
wire n_7254;
wire n_18178;
wire n_12973;
wire n_17313;
wire n_13123;
wire n_14669;
wire n_12234;
wire n_10776;
wire n_7882;
wire n_16348;
wire n_16514;
wire n_17704;
wire n_10848;
wire n_20216;
wire n_7765;
wire n_11482;
wire n_7816;
wire n_10164;
wire n_15809;
wire n_15579;
wire n_18549;
wire n_18084;
wire n_15585;
wire n_12033;
wire n_14376;
wire n_20102;
wire n_20173;
wire n_9595;
wire n_18978;
wire n_15555;
wire n_13923;
wire n_13051;
wire n_11524;
wire n_17220;
wire n_9265;
wire n_8239;
wire n_16114;
wire n_13330;
wire n_11228;
wire n_7898;
wire n_18286;
wire n_9789;
wire n_7646;
wire n_20166;
wire n_17537;
wire n_14627;
wire n_13699;
wire n_19940;
wire n_7665;
wire n_9354;
wire n_10501;
wire n_14026;
wire n_17782;
wire n_19687;
wire n_9436;
wire n_18157;
wire n_8489;
wire n_10350;
wire n_12730;
wire n_6887;
wire n_18926;
wire n_16123;
wire n_13152;
wire n_17221;
wire n_6637;
wire n_9238;
wire n_6633;
wire n_11031;
wire n_17365;
wire n_9839;
wire n_18479;
wire n_15704;
wire n_7900;
wire n_6569;
wire n_10807;
wire n_12478;
wire n_17265;
wire n_13545;
wire n_13760;
wire n_13883;
wire n_10511;
wire n_7576;
wire n_19499;
wire n_11023;
wire n_7313;
wire n_10873;
wire n_14484;
wire n_7676;
wire n_18956;
wire n_9017;
wire n_15726;
wire n_14307;
wire n_8865;
wire n_15302;
wire n_10337;
wire n_7779;
wire n_8999;
wire n_11626;
wire n_12148;
wire n_16872;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_16312;
wire n_16204;
wire n_8820;
wire n_16793;
wire n_16443;
wire n_6090;
wire n_20071;
wire n_18456;
wire n_18281;
wire n_12132;
wire n_10593;
wire n_16801;
wire n_12182;
wire n_12043;
wire n_10636;
wire n_16478;
wire n_18489;
wire n_18723;
wire n_8992;
wire n_8880;
wire n_8690;
wire n_6234;
wire n_7818;
wire n_11721;
wire n_13573;
wire n_19019;
wire n_6608;
wire n_9109;
wire n_7896;
wire n_12482;
wire n_18839;
wire n_15208;
wire n_6860;
wire n_12137;
wire n_12306;
wire n_11328;
wire n_11200;
wire n_14442;
wire n_15210;
wire n_16536;
wire n_19917;
wire n_13418;
wire n_7996;
wire n_10533;
wire n_16681;
wire n_10176;
wire n_19707;
wire n_7517;
wire n_8080;
wire n_12345;
wire n_13551;
wire n_19135;
wire n_19178;
wire n_16060;
wire n_8772;
wire n_8786;
wire n_15597;
wire n_12694;
wire n_8083;
wire n_20060;
wire n_10155;
wire n_9805;
wire n_19799;
wire n_13593;
wire n_8157;
wire n_19660;
wire n_13902;
wire n_19792;
wire n_9110;
wire n_18358;
wire n_14468;
wire n_12550;
wire n_13861;
wire n_13350;
wire n_10051;
wire n_10414;
wire n_8344;
wire n_17597;
wire n_8120;
wire n_9075;
wire n_12961;
wire n_18882;
wire n_11496;
wire n_12225;
wire n_20118;
wire n_8621;
wire n_12884;
wire n_20350;
wire n_19171;
wire n_6246;
wire n_8868;
wire n_8134;
wire n_12207;
wire n_9975;
wire n_20595;
wire n_12011;
wire n_7252;
wire n_20031;
wire n_6843;
wire n_10626;
wire n_6901;
wire n_19014;
wire n_13273;
wire n_18855;
wire n_8101;
wire n_19751;
wire n_19954;
wire n_6489;
wire n_7402;
wire n_19552;
wire n_11273;
wire n_19089;
wire n_19993;
wire n_16954;
wire n_12472;
wire n_19526;
wire n_14035;
wire n_13218;
wire n_9081;
wire n_11762;
wire n_9236;
wire n_6844;
wire n_10156;
wire n_9607;
wire n_6779;
wire n_10774;
wire n_12332;
wire n_7216;
wire n_15990;
wire n_15364;
wire n_6543;
wire n_19585;
wire n_6178;
wire n_9621;
wire n_18075;
wire n_16117;
wire n_10398;
wire n_17947;
wire n_16459;
wire n_17987;
wire n_18165;
wire n_15661;
wire n_20185;
wire n_17932;
wire n_7706;
wire n_20304;
wire n_6458;
wire n_7642;
wire n_12506;
wire n_18356;
wire n_12718;
wire n_12638;
wire n_14116;
wire n_20391;
wire n_18710;
wire n_16453;
wire n_16645;
wire n_10470;
wire n_20156;
wire n_15034;
wire n_19808;
wire n_14240;
wire n_14504;
wire n_13449;
wire n_12747;
wire n_10625;
wire n_12561;
wire n_18420;
wire n_8388;
wire n_18469;
wire n_14730;
wire n_18732;
wire n_9589;
wire n_10445;
wire n_15110;
wire n_8988;
wire n_15025;
wire n_19329;
wire n_18161;
wire n_12900;
wire n_18761;
wire n_8569;
wire n_14598;
wire n_10679;
wire n_11323;
wire n_10799;
wire n_17228;
wire n_10585;
wire n_18519;
wire n_13696;
wire n_12948;
wire n_7931;
wire n_13322;
wire n_9092;
wire n_10034;
wire n_9451;
wire n_11148;
wire n_18729;
wire n_13934;
wire n_6899;
wire n_19880;
wire n_7373;
wire n_7895;
wire n_15331;
wire n_17109;
wire n_13254;
wire n_15191;
wire n_17617;
wire n_8951;
wire n_18783;
wire n_15676;
wire n_17044;
wire n_9011;
wire n_7613;
wire n_6101;
wire n_14440;
wire n_7556;
wire n_10528;
wire n_20168;
wire n_13875;
wire n_17319;
wire n_17774;
wire n_19255;
wire n_14076;
wire n_11220;
wire n_17709;
wire n_9012;
wire n_18150;
wire n_14638;
wire n_19803;
wire n_7238;
wire n_14936;
wire n_16469;
wire n_8047;
wire n_11596;
wire n_6273;
wire n_7572;
wire n_11955;
wire n_20535;
wire n_18818;
wire n_16156;
wire n_11654;
wire n_18361;
wire n_12982;
wire n_11619;
wire n_10649;
wire n_19638;
wire n_6311;
wire n_7590;
wire n_12275;
wire n_13742;
wire n_15177;
wire n_12376;
wire n_13114;
wire n_8583;
wire n_10447;
wire n_15063;
wire n_7176;
wire n_9353;
wire n_13054;
wire n_8948;
wire n_8295;
wire n_10522;
wire n_13793;
wire n_11782;
wire n_16532;
wire n_20590;
wire n_16618;
wire n_10278;
wire n_15384;
wire n_13882;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_15686;
wire n_9263;
wire n_11082;
wire n_15950;
wire n_19724;
wire n_6181;
wire n_7447;
wire n_17998;
wire n_19156;
wire n_18928;
wire n_12721;
wire n_18301;
wire n_16008;
wire n_11730;
wire n_6924;
wire n_9804;
wire n_9304;
wire n_8380;
wire n_12039;
wire n_10377;
wire n_9926;
wire n_15161;
wire n_10858;
wire n_16303;
wire n_9843;
wire n_16559;
wire n_13320;
wire n_6683;
wire n_10683;
wire n_9921;
wire n_19606;
wire n_6229;
wire n_13488;
wire n_15907;
wire n_7286;
wire n_13668;
wire n_13016;
wire n_6177;
wire n_16961;
wire n_14708;
wire n_17293;
wire n_12048;
wire n_10930;
wire n_17972;
wire n_8749;
wire n_18264;
wire n_12057;
wire n_6696;
wire n_17590;
wire n_9527;
wire n_16450;
wire n_19651;
wire n_18352;
wire n_14875;
wire n_15860;
wire n_15056;
wire n_19460;
wire n_17288;
wire n_16197;
wire n_14003;
wire n_9511;
wire n_6730;
wire n_17822;
wire n_13670;
wire n_11254;
wire n_15023;
wire n_11617;
wire n_18184;
wire n_18436;
wire n_6170;
wire n_9459;
wire n_14185;
wire n_6094;
wire n_9098;
wire n_14953;
wire n_15604;
wire n_16000;
wire n_12360;
wire n_9268;
wire n_17116;
wire n_20497;
wire n_15431;
wire n_8673;
wire n_18702;
wire n_19174;
wire n_10456;
wire n_13186;
wire n_18824;
wire n_15655;
wire n_11907;
wire n_10627;
wire n_10475;
wire n_20373;
wire n_15430;
wire n_20578;
wire n_8581;
wire n_15732;
wire n_12457;
wire n_16070;
wire n_16045;
wire n_17772;
wire n_14170;
wire n_13496;
wire n_8058;
wire n_9308;
wire n_11838;
wire n_10508;
wire n_18008;
wire n_10811;
wire n_18696;
wire n_8333;
wire n_17152;
wire n_7619;
wire n_6985;
wire n_18551;
wire n_7170;
wire n_13853;
wire n_8823;
wire n_11457;
wire n_12751;
wire n_15284;
wire n_20374;
wire n_17901;
wire n_15443;
wire n_18228;
wire n_17833;
wire n_18471;
wire n_16852;
wire n_18817;
wire n_6916;
wire n_15524;
wire n_10725;
wire n_7845;
wire n_12688;
wire n_18354;
wire n_8290;
wire n_7536;
wire n_18152;
wire n_6230;
wire n_16108;
wire n_11107;
wire n_12757;
wire n_14379;
wire n_8840;
wire n_16284;
wire n_16001;
wire n_18873;
wire n_13189;
wire n_18915;
wire n_19492;
wire n_12328;
wire n_9083;
wire n_17271;
wire n_6483;
wire n_10994;
wire n_14004;
wire n_17023;
wire n_16221;
wire n_8036;
wire n_11485;
wire n_7300;
wire n_6975;
wire n_14666;
wire n_13605;
wire n_17387;
wire n_11048;
wire n_14237;
wire n_6729;
wire n_11240;
wire n_13841;
wire n_11634;
wire n_12580;
wire n_10013;
wire n_17166;
wire n_20608;
wire n_16119;
wire n_6076;
wire n_8933;
wire n_19344;
wire n_15876;
wire n_18819;
wire n_15231;
wire n_11287;
wire n_9774;
wire n_6390;
wire n_19846;
wire n_13409;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_9720;
wire n_15727;
wire n_10169;
wire n_12690;
wire n_7563;
wire n_12475;
wire n_11765;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_19510;
wire n_14414;
wire n_15565;
wire n_17823;
wire n_9149;
wire n_7035;
wire n_6193;
wire n_16858;
wire n_16980;
wire n_9345;
wire n_11550;
wire n_17315;
wire n_7527;
wire n_13061;
wire n_9682;
wire n_17719;
wire n_6582;
wire n_18432;
wire n_12545;
wire n_20390;
wire n_18320;
wire n_18078;
wire n_9924;
wire n_14744;
wire n_15091;
wire n_17527;
wire n_12753;
wire n_7090;
wire n_9254;
wire n_11641;
wire n_7415;
wire n_11211;
wire n_13691;
wire n_13375;
wire n_6745;
wire n_6972;
wire n_18526;
wire n_16913;
wire n_16663;
wire n_11857;
wire n_6240;
wire n_13482;
wire n_18069;
wire n_15778;
wire n_7121;
wire n_9469;
wire n_15869;
wire n_15598;
wire n_15988;
wire n_16593;
wire n_6515;
wire n_16604;
wire n_13873;
wire n_15805;
wire n_17836;
wire n_18769;
wire n_11201;
wire n_10531;
wire n_14964;
wire n_8918;
wire n_12878;
wire n_19273;
wire n_8932;
wire n_17756;
wire n_16603;
wire n_9249;
wire n_8180;
wire n_20624;
wire n_20191;
wire n_15580;
wire n_9444;
wire n_10772;
wire n_7114;
wire n_15984;
wire n_6770;
wire n_20237;
wire n_20124;
wire n_17730;
wire n_15151;
wire n_16626;
wire n_8943;
wire n_14767;
wire n_18463;
wire n_20343;
wire n_14773;
wire n_10127;
wire n_13654;
wire n_11814;
wire n_12255;
wire n_9723;
wire n_19446;
wire n_19669;
wire n_19834;
wire n_19577;
wire n_7199;
wire n_10039;
wire n_10854;
wire n_11358;
wire n_13366;
wire n_7940;
wire n_16467;
wire n_6782;
wire n_18746;
wire n_17669;
wire n_6503;
wire n_19423;
wire n_12017;
wire n_17357;
wire n_15381;
wire n_18477;
wire n_11958;
wire n_6621;
wire n_15624;
wire n_16103;
wire n_19041;
wire n_16460;
wire n_8271;
wire n_20303;
wire n_12728;
wire n_16651;
wire n_6783;
wire n_19963;
wire n_12259;
wire n_8699;
wire n_16305;
wire n_19409;
wire n_19932;
wire n_15861;
wire n_8225;
wire n_9536;
wire n_14250;
wire n_16818;
wire n_16573;
wire n_18671;
wire n_16562;
wire n_6296;
wire n_7708;
wire n_11671;
wire n_10328;
wire n_6497;
wire n_15705;
wire n_16816;
wire n_7333;
wire n_15376;
wire n_8546;
wire n_10963;
wire n_16358;
wire n_18035;
wire n_7371;
wire n_17547;
wire n_8152;
wire n_15050;
wire n_10826;
wire n_7463;
wire n_8525;
wire n_17767;
wire n_18680;
wire n_12160;
wire n_9620;
wire n_17145;
wire n_11119;
wire n_7954;
wire n_7951;
wire n_8096;
wire n_13901;
wire n_7231;
wire n_15252;
wire n_18043;
wire n_20465;
wire n_16238;
wire n_14050;
wire n_15763;
wire n_17983;
wire n_15317;
wire n_7772;
wire n_14197;
wire n_18159;
wire n_19364;
wire n_8996;
wire n_12070;
wire n_9714;
wire n_14898;
wire n_15672;
wire n_20532;
wire n_20623;
wire n_15920;
wire n_11928;
wire n_14395;
wire n_13528;
wire n_8292;
wire n_8601;
wire n_9377;
wire n_11932;
wire n_6970;
wire n_19328;
wire n_13027;
wire n_20342;
wire n_12607;
wire n_7272;
wire n_15782;
wire n_19553;
wire n_12075;
wire n_13489;
wire n_18887;
wire n_19693;
wire n_19797;
wire n_13877;
wire n_6209;
wire n_11922;
wire n_14020;
wire n_12358;
wire n_7408;
wire n_10488;
wire n_8969;
wire n_14187;
wire n_11577;
wire n_17840;
wire n_16914;
wire n_18513;
wire n_19165;
wire n_17907;
wire n_11475;
wire n_9048;
wire n_10274;
wire n_6694;
wire n_15318;
wire n_9168;
wire n_14220;
wire n_13837;
wire n_20640;
wire n_18570;
wire n_15559;
wire n_16871;
wire n_14221;
wire n_13964;
wire n_10832;
wire n_18829;
wire n_6856;
wire n_6466;
wire n_16039;
wire n_7864;
wire n_18295;
wire n_6727;
wire n_14360;
wire n_10584;
wire n_13601;
wire n_17457;
wire n_17115;
wire n_19281;
wire n_18155;
wire n_6820;
wire n_17083;
wire n_19007;
wire n_13392;
wire n_17563;
wire n_9169;
wire n_10229;
wire n_7512;
wire n_19008;
wire n_18401;
wire n_6469;
wire n_6700;
wire n_20494;
wire n_6223;
wire n_11398;
wire n_8798;
wire n_9600;
wire n_8085;
wire n_11274;
wire n_8123;
wire n_17997;
wire n_12512;
wire n_9927;
wire n_16973;
wire n_15657;
wire n_17571;
wire n_7127;
wire n_15513;
wire n_8666;
wire n_12284;
wire n_18322;
wire n_7801;
wire n_9155;
wire n_10416;
wire n_15837;
wire n_14370;
wire n_7959;
wire n_13430;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_10583;
wire n_10806;
wire n_7546;
wire n_6272;
wire n_14274;
wire n_6588;
wire n_18125;
wire n_15403;
wire n_13081;
wire n_15602;
wire n_12252;
wire n_16743;
wire n_10439;
wire n_12627;
wire n_19378;
wire n_16730;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_20012;
wire n_18868;
wire n_6222;
wire n_15012;
wire n_20451;
wire n_14551;
wire n_15720;
wire n_11181;
wire n_13651;
wire n_7521;
wire n_12968;
wire n_10663;
wire n_15517;
wire n_13974;
wire n_12277;
wire n_14917;
wire n_16075;
wire n_6625;
wire n_15680;
wire n_17441;
wire n_14855;
wire n_16757;
wire n_8487;
wire n_18601;
wire n_8141;
wire n_14058;
wire n_11020;
wire n_13141;
wire n_16461;
wire n_14065;
wire n_11920;
wire n_19756;
wire n_17299;
wire n_14366;
wire n_10481;
wire n_19250;
wire n_6876;
wire n_16022;
wire n_19001;
wire n_19627;
wire n_9573;
wire n_7636;
wire n_9799;
wire n_17235;
wire n_6954;
wire n_6938;
wire n_15143;
wire n_11198;
wire n_18932;
wire n_18346;
wire n_18238;
wire n_19794;
wire n_11840;
wire n_13157;
wire n_10261;
wire n_14084;
wire n_9827;
wire n_13334;
wire n_10907;
wire n_14002;
wire n_19842;
wire n_19892;
wire n_7214;
wire n_16205;
wire n_13399;
wire n_19984;
wire n_7075;
wire n_19503;
wire n_14697;
wire n_7124;
wire n_13967;
wire n_20506;
wire n_7799;
wire n_11092;
wire n_14310;
wire n_15792;
wire n_15281;
wire n_15675;
wire n_8917;
wire n_9647;
wire n_15515;
wire n_15106;
wire n_12067;
wire n_9214;
wire n_17030;
wire n_19537;
wire n_7776;
wire n_19621;
wire n_14309;
wire n_9864;
wire n_16256;
wire n_17416;
wire n_16741;
wire n_11770;
wire n_19201;
wire n_13996;
wire n_19904;
wire n_19853;
wire n_17944;
wire n_17679;
wire n_9000;
wire n_18442;
wire n_18505;
wire n_10864;
wire n_18412;
wire n_14704;
wire n_8307;
wire n_9383;
wire n_17692;
wire n_15258;
wire n_12174;
wire n_16322;
wire n_15220;
wire n_6400;
wire n_19611;
wire n_16304;
wire n_18417;
wire n_7543;
wire n_13504;
wire n_16787;
wire n_13169;
wire n_7877;
wire n_9672;
wire n_15291;
wire n_8855;
wire n_18375;
wire n_8885;
wire n_15345;
wire n_14721;
wire n_13265;
wire n_12153;
wire n_7284;
wire n_7264;
wire n_13666;
wire n_19192;
wire n_6537;
wire n_20408;
wire n_10702;
wire n_20613;
wire n_13730;
wire n_12405;
wire n_10319;
wire n_9654;
wire n_8802;
wire n_9859;
wire n_6092;
wire n_6241;
wire n_8667;
wire n_18996;
wire n_8121;
wire n_9645;
wire n_7754;
wire n_15549;
wire n_18777;
wire n_12792;
wire n_19661;
wire n_9796;
wire n_8320;
wire n_18219;
wire n_18231;
wire n_15889;
wire n_11830;
wire n_12438;
wire n_8766;
wire n_16173;
wire n_16665;
wire n_9165;
wire n_19555;
wire n_12539;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_18461;
wire n_14369;
wire n_7240;
wire n_15354;
wire n_10476;
wire n_9966;
wire n_16794;
wire n_11486;
wire n_15999;
wire n_15280;
wire n_12677;
wire n_7237;
wire n_17867;
wire n_16456;
wire n_6877;
wire n_12873;
wire n_16364;
wire n_6949;
wire n_20531;
wire n_19356;
wire n_17036;
wire n_19698;
wire n_13401;
wire n_12276;
wire n_9893;
wire n_14122;
wire n_17565;
wire n_8126;
wire n_15819;
wire n_10362;
wire n_9239;
wire n_15603;
wire n_12352;
wire n_17267;
wire n_18528;
wire n_10099;
wire n_9961;
wire n_16833;
wire n_14895;
wire n_7163;
wire n_16582;
wire n_18028;
wire n_15270;
wire n_17964;
wire n_10181;
wire n_15670;
wire n_19974;
wire n_7201;
wire n_16825;
wire n_20274;
wire n_10949;
wire n_18197;
wire n_13969;
wire n_16548;
wire n_12693;
wire n_6792;
wire n_20594;
wire n_9316;
wire n_13259;
wire n_19164;
wire n_14954;
wire n_12648;
wire n_9914;
wire n_8132;
wire n_19541;
wire n_20433;
wire n_10917;
wire n_16050;
wire n_18006;
wire n_7821;
wire n_12407;
wire n_11284;
wire n_20100;
wire n_14668;
wire n_14776;
wire n_10458;
wire n_11656;
wire n_13134;
wire n_10271;
wire n_15415;
wire n_20315;
wire n_16808;
wire n_18902;
wire n_6673;
wire n_20026;
wire n_18207;
wire n_11909;
wire n_12637;
wire n_7887;
wire n_15414;
wire n_15783;
wire n_12009;
wire n_13612;
wire n_19388;
wire n_10648;
wire n_7550;
wire n_17498;
wire n_15077;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_15733;
wire n_15864;
wire n_14207;
wire n_19080;
wire n_19736;
wire n_13863;
wire n_14305;
wire n_9863;
wire n_15330;
wire n_10500;
wire n_15261;
wire n_11929;
wire n_11075;
wire n_7851;
wire n_16605;
wire n_20372;
wire n_9791;
wire n_19228;
wire n_11177;
wire n_19761;
wire n_13667;
wire n_18056;
wire n_13126;
wire n_7798;
wire n_10857;
wire n_18491;
wire n_11310;
wire n_13275;
wire n_11165;
wire n_14411;
wire n_20503;
wire n_12823;
wire n_15412;
wire n_20331;
wire n_12193;
wire n_6088;
wire n_15257;
wire n_19701;
wire n_8528;
wire n_8204;
wire n_11733;
wire n_15646;
wire n_18214;
wire n_7100;
wire n_18347;
wire n_14738;
wire n_12242;
wire n_20108;
wire n_13796;
wire n_10502;
wire n_15522;
wire n_17577;
wire n_17874;
wire n_6722;
wire n_17892;
wire n_7622;
wire n_11123;
wire n_8512;
wire n_14464;
wire n_8635;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_15535;
wire n_16633;
wire n_7831;
wire n_10227;
wire n_10574;
wire n_19271;
wire n_16323;
wire n_18624;
wire n_6201;
wire n_12218;
wire n_12343;
wire n_8919;
wire n_17014;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_11478;
wire n_16067;
wire n_15650;
wire n_12236;
wire n_12902;
wire n_16230;
wire n_7784;
wire n_9272;
wire n_13038;
wire n_12892;
wire n_17768;
wire n_11294;
wire n_15667;
wire n_19861;
wire n_10289;
wire n_6565;
wire n_6942;
wire n_11819;
wire n_19389;
wire n_13420;
wire n_6862;
wire n_17200;
wire n_15053;
wire n_13005;
wire n_14805;
wire n_20575;
wire n_11844;
wire n_15390;
wire n_6635;
wire n_13184;
wire n_13535;
wire n_14982;
wire n_12247;
wire n_14770;
wire n_11100;
wire n_19350;
wire n_7167;
wire n_6480;
wire n_15105;
wire n_18927;
wire n_18383;
wire n_12765;
wire n_7865;
wire n_15690;
wire n_9289;
wire n_11315;
wire n_6561;
wire n_12706;
wire n_19949;
wire n_11153;
wire n_17128;
wire n_6875;
wire n_10934;
wire n_10197;
wire n_18999;
wire n_19584;
wire n_11949;
wire n_8402;
wire n_9690;
wire n_11746;
wire n_9371;
wire n_19689;
wire n_19990;
wire n_16837;
wire n_20095;
wire n_7267;
wire n_12315;
wire n_18668;
wire n_7850;
wire n_14100;
wire n_12998;
wire n_7812;
wire n_13143;
wire n_9080;
wire n_14549;
wire n_8133;
wire n_6176;
wire n_14717;
wire n_16426;
wire n_14459;
wire n_11530;
wire n_13411;
wire n_7056;
wire n_8193;
wire n_12445;
wire n_12856;
wire n_19520;
wire n_7813;
wire n_7514;
wire n_7649;
wire n_18734;
wire n_12525;
wire n_16116;
wire n_6078;
wire n_15823;
wire n_13758;
wire n_7688;
wire n_16820;
wire n_8707;
wire n_12357;
wire n_9208;
wire n_11791;
wire n_19525;
wire n_7611;
wire n_19778;
wire n_17218;
wire n_15216;
wire n_11848;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_12180;
wire n_15608;
wire n_10935;
wire n_20044;
wire n_7723;
wire n_11621;
wire n_19448;
wire n_16171;
wire n_7450;
wire n_11667;
wire n_17311;
wire n_7362;
wire n_17455;
wire n_12208;
wire n_14565;
wire n_17248;
wire n_11298;
wire n_15796;
wire n_8993;
wire n_6204;
wire n_13314;
wire n_11741;
wire n_15537;
wire n_12773;
wire n_9044;
wire n_12381;
wire n_19885;
wire n_19302;
wire n_18174;
wire n_14883;
wire n_17024;
wire n_6451;
wire n_9813;
wire n_18482;
wire n_20217;
wire n_17322;
wire n_9244;
wire n_15304;
wire n_7049;
wire n_15271;
wire n_14865;
wire n_8278;
wire n_11644;
wire n_6345;
wire n_15893;
wire n_9094;
wire n_15432;
wire n_13108;
wire n_13170;
wire n_14471;
wire n_11357;
wire n_19387;
wire n_9985;
wire n_12089;
wire n_20104;
wire n_7057;
wire n_17888;
wire n_11959;
wire n_19586;
wire n_12987;
wire n_8529;
wire n_10254;
wire n_18625;
wire n_14715;
wire n_15970;
wire n_11208;
wire n_15978;
wire n_12452;
wire n_20495;
wire n_15961;
wire n_8574;
wire n_12292;
wire n_12818;
wire n_11420;
wire n_12500;
wire n_8044;
wire n_16330;
wire n_9439;
wire n_15239;
wire n_11630;
wire n_19759;
wire n_15444;
wire n_15289;
wire n_13172;
wire n_16234;
wire n_9120;
wire n_17335;
wire n_17610;
wire n_19522;
wire n_12168;
wire n_16496;
wire n_8903;
wire n_16057;
wire n_16401;
wire n_15781;
wire n_14448;
wire n_11017;
wire n_7247;
wire n_14622;
wire n_7893;
wire n_6213;
wire n_19924;
wire n_14739;
wire n_16649;
wire n_12613;
wire n_14365;
wire n_9325;
wire n_16448;
wire n_17173;
wire n_9384;
wire n_6216;
wire n_7340;
wire n_12695;
wire n_15467;
wire n_14219;
wire n_11576;
wire n_12006;
wire n_10128;
wire n_18319;
wire n_12246;
wire n_18220;
wire n_9955;
wire n_19477;
wire n_9007;
wire n_10143;
wire n_18715;
wire n_17884;
wire n_13085;
wire n_19260;
wire n_7780;
wire n_20413;
wire n_8452;
wire n_11518;
wire n_8557;
wire n_10303;
wire n_16189;
wire n_15097;
wire n_18892;
wire n_11252;
wire n_8012;
wire n_17055;
wire n_6472;
wire n_18067;
wire n_8114;
wire n_16227;
wire n_14563;
wire n_16329;
wire n_11256;
wire n_6166;
wire n_12370;
wire n_9136;
wire n_12860;
wire n_16278;
wire n_17404;
wire n_19635;
wire n_7063;
wire n_14768;
wire n_13885;
wire n_20364;
wire n_13631;
wire n_18103;
wire n_6081;
wire n_16746;
wire n_15929;
wire n_6724;
wire n_11336;
wire n_12758;
wire n_17410;
wire n_19248;
wire n_11849;
wire n_9204;
wire n_9476;
wire n_12142;
wire n_9689;
wire n_16711;
wire n_10659;
wire n_7585;
wire n_6946;
wire n_12983;
wire n_6424;
wire n_11210;
wire n_7599;
wire n_16271;
wire n_15541;
wire n_13980;
wire n_16366;
wire n_11191;
wire n_10547;
wire n_6778;
wire n_17359;
wire n_13205;
wire n_20629;
wire n_15283;
wire n_12396;
wire n_15407;
wire n_7614;
wire n_19381;
wire n_7839;
wire n_9837;
wire n_10896;
wire n_17761;
wire n_10562;
wire n_16042;
wire n_14417;
wire n_6340;
wire n_10054;
wire n_10355;
wire n_16893;
wire n_6706;
wire n_13034;
wire n_16828;
wire n_10007;
wire n_11751;
wire n_17550;
wire n_17185;
wire n_20286;
wire n_20597;
wire n_14637;
wire n_11495;
wire n_17015;
wire n_7372;
wire n_19617;
wire n_17980;
wire n_17535;
wire n_16822;
wire n_10704;
wire n_11520;
wire n_19614;
wire n_12169;
wire n_16788;
wire n_15088;
wire n_17976;
wire n_16383;
wire n_17538;
wire n_11012;
wire n_6111;
wire n_11502;
wire n_15348;
wire n_11631;
wire n_13588;
wire n_13570;
wire n_20176;
wire n_20038;
wire n_11842;
wire n_14710;
wire n_13737;
wire n_16590;
wire n_18188;
wire n_16640;
wire n_11389;
wire n_7226;
wire n_9013;
wire n_18373;
wire n_9634;
wire n_17846;
wire n_10916;
wire n_8584;
wire n_11557;
wire n_17113;
wire n_16748;
wire n_15363;
wire n_7810;
wire n_14955;
wire n_9364;
wire n_8228;
wire n_16015;
wire n_15642;
wire n_10929;
wire n_18854;
wire n_19372;
wire n_13862;
wire n_8100;
wire n_13446;
wire n_13086;
wire n_8091;
wire n_17155;
wire n_20236;
wire n_14965;
wire n_13887;
wire n_12787;
wire n_12799;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_15205;
wire n_8158;
wire n_8469;
wire n_18718;
wire n_18481;
wire n_10102;
wire n_11825;
wire n_14354;
wire n_7684;
wire n_15532;
wire n_16083;
wire n_10589;
wire n_11611;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_18221;
wire n_12408;
wire n_16287;
wire n_16169;
wire n_19314;
wire n_17556;
wire n_10110;
wire n_11230;
wire n_11688;
wire n_12715;
wire n_12434;
wire n_11709;
wire n_14328;
wire n_6095;
wire n_17049;
wire n_18938;
wire n_16540;
wire n_14429;
wire n_12979;
wire n_16901;
wire n_6559;
wire n_15799;
wire n_19733;
wire n_17195;
wire n_19050;
wire n_14270;
wire n_15238;
wire n_10190;
wire n_19656;
wire n_6287;
wire n_13614;
wire n_8347;
wire n_17703;
wire n_19440;
wire n_14208;
wire n_9330;
wire n_20399;
wire n_15693;
wire n_12029;
wire n_9523;
wire n_14584;
wire n_19636;
wire n_10060;
wire n_18192;
wire n_9686;
wire n_20434;
wire n_17130;
wire n_19375;
wire n_10162;
wire n_15002;
wire n_9964;
wire n_17515;
wire n_13842;
wire n_7510;
wire n_6662;
wire n_11291;
wire n_9154;
wire n_13107;
wire n_14501;
wire n_7109;
wire n_8822;
wire n_14790;
wire n_17204;
wire n_12187;
wire n_19662;
wire n_20121;
wire n_18772;
wire n_7253;
wire n_17201;
wire n_8476;
wire n_17745;
wire n_11927;
wire n_16674;
wire n_16326;
wire n_16571;
wire n_8359;
wire n_15808;
wire n_16497;
wire n_16752;
wire n_14574;
wire n_14451;
wire n_9455;
wire n_8708;
wire n_14092;
wire n_14509;
wire n_11882;
wire n_17649;
wire n_11647;
wire n_15027;
wire n_15404;
wire n_10706;
wire n_19129;
wire n_8872;
wire n_20120;
wire n_19746;
wire n_8238;
wire n_20626;
wire n_15465;
wire n_20318;
wire n_11222;
wire n_9200;
wire n_16279;
wire n_15858;
wire n_18946;
wire n_14765;
wire n_7704;
wire n_18893;
wire n_16170;
wire n_14995;
wire n_6302;
wire n_17479;
wire n_7203;
wire n_11259;
wire n_7670;
wire n_18258;
wire n_16010;
wire n_9673;
wire n_14434;
wire n_20252;
wire n_8642;
wire n_11875;
wire n_18567;
wire n_12111;
wire n_8912;
wire n_19067;
wire n_14275;
wire n_19309;
wire n_12903;
wire n_6343;
wire n_12593;
wire n_20051;
wire n_17849;
wire n_20588;
wire n_11602;
wire n_15689;
wire n_19850;
wire n_12413;
wire n_17474;
wire n_13813;
wire n_16190;
wire n_8111;
wire n_18315;
wire n_10432;
wire n_19227;
wire n_16888;
wire n_8056;
wire n_18376;
wire n_9674;
wire n_6433;
wire n_18253;
wire n_15469;
wire n_17140;
wire n_18407;
wire n_18816;
wire n_13636;
wire n_19332;
wire n_19456;
wire n_18920;
wire n_11341;
wire n_10787;
wire n_13256;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_16308;
wire n_6279;
wire n_13905;
wire n_12290;
wire n_20558;
wire n_7881;
wire n_9369;
wire n_18896;
wire n_16986;
wire n_17872;
wire n_9583;
wire n_19422;
wire n_19858;
wire n_15119;
wire n_19117;
wire n_12150;
wire n_15256;
wire n_18366;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_15982;
wire n_19643;
wire n_18647;
wire n_15452;
wire n_13615;
wire n_15625;
wire n_12633;
wire n_14779;
wire n_15114;
wire n_10277;
wire n_17934;
wire n_8163;
wire n_16632;
wire n_16028;
wire n_19862;
wire n_10948;
wire n_10525;
wire n_14287;
wire n_9507;
wire n_11528;
wire n_15296;
wire n_15828;
wire n_18107;
wire n_19211;
wire n_16126;
wire n_18102;
wire n_19699;
wire n_18545;
wire n_16168;
wire n_15915;
wire n_10049;
wire n_15551;
wire n_9457;
wire n_16738;
wire n_6084;
wire n_11039;
wire n_14342;
wire n_13693;
wire n_18992;
wire n_12606;
wire n_10900;
wire n_14107;
wire n_14781;
wire n_13333;
wire n_13229;
wire n_17336;
wire n_11380;
wire n_15737;
wire n_19567;
wire n_10792;
wire n_15573;
wire n_13296;
wire n_20617;
wire n_14611;
wire n_17863;
wire n_20165;
wire n_20196;
wire n_17088;
wire n_19100;
wire n_15051;
wire n_6548;
wire n_20383;
wire n_6993;
wire n_15916;
wire n_16468;
wire n_10241;
wire n_19598;
wire n_15639;
wire n_8702;
wire n_17158;
wire n_8116;
wire n_7946;
wire n_8195;
wire n_14069;
wire n_18452;
wire n_19786;
wire n_9991;
wire n_11366;
wire n_11872;
wire n_19901;
wire n_10823;
wire n_19685;
wire n_14766;
wire n_11106;
wire n_14592;
wire n_15109;
wire n_11132;
wire n_17625;
wire n_18546;
wire n_18034;
wire n_18181;
wire n_17126;
wire n_10824;
wire n_19566;
wire n_16216;
wire n_19398;
wire n_14277;
wire n_19565;
wire n_13493;
wire n_16389;
wire n_9047;
wire n_12842;
wire n_18569;
wire n_12481;
wire n_18168;
wire n_11316;
wire n_9599;
wire n_11559;
wire n_9072;
wire n_19811;
wire n_9428;
wire n_10340;
wire n_17463;
wire n_15817;
wire n_15344;
wire n_13669;
wire n_17245;
wire n_17179;
wire n_11109;
wire n_13840;
wire n_16601;
wire n_20199;
wire n_11591;
wire n_19710;
wire n_14251;
wire n_11225;
wire n_6765;
wire n_8883;
wire n_10634;
wire n_11058;
wire n_15888;
wire n_7336;
wire n_11471;
wire n_7446;
wire n_14679;
wire n_10961;
wire n_7357;
wire n_20301;
wire n_17064;
wire n_8737;
wire n_13925;
wire n_18334;
wire n_10379;
wire n_16704;
wire n_18223;
wire n_13368;
wire n_14507;
wire n_9484;
wire n_10989;
wire n_17725;
wire n_10939;
wire n_19557;
wire n_11144;
wire n_14857;
wire n_6406;
wire n_14034;
wire n_10962;
wire n_11128;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_11025;
wire n_12007;
wire n_15901;
wire n_13481;
wire n_12018;
wire n_18040;
wire n_17393;
wire n_14457;
wire n_16931;
wire n_12872;
wire n_18189;
wire n_6492;
wire n_14517;
wire n_11460;
wire n_13713;
wire n_12372;
wire n_13608;
wire n_7046;
wire n_19059;
wire n_10956;
wire n_7468;
wire n_18785;
wire n_14934;
wire n_19663;
wire n_18844;
wire n_12572;
wire n_12453;
wire n_19968;
wire n_19752;
wire n_17870;
wire n_15652;
wire n_19466;
wire n_16713;
wire n_14578;
wire n_15653;
wire n_12955;
wire n_9321;
wire n_16856;
wire n_18555;
wire n_15016;
wire n_18493;
wire n_9161;
wire n_7836;
wire n_10737;
wire n_17910;
wire n_17750;
wire n_15865;
wire n_13448;
wire n_16928;
wire n_13767;
wire n_11055;
wire n_16616;
wire n_14832;
wire n_10982;
wire n_17599;
wire n_14571;
wire n_6631;
wire n_12369;
wire n_7577;
wire n_7308;
wire n_8927;
wire n_17985;
wire n_16396;
wire n_17531;
wire n_15155;
wire n_12686;
wire n_6228;
wire n_19336;
wire n_14881;
wire n_18588;
wire n_14527;
wire n_12822;
wire n_13307;
wire n_7279;
wire n_17460;
wire n_13312;
wire n_11761;
wire n_8474;
wire n_9984;
wire n_10600;
wire n_6102;
wire n_10833;
wire n_18329;
wire n_18649;
wire n_13023;
wire n_20382;
wire n_19343;
wire n_15315;
wire n_19210;
wire n_11185;
wire n_13440;
wire n_13436;
wire n_19615;
wire n_19133;
wire n_16982;
wire n_11081;
wire n_16687;
wire n_14858;
wire n_8787;
wire n_13911;
wire n_17544;
wire n_20241;
wire n_10941;
wire n_14617;
wire n_9816;
wire n_17132;
wire n_14263;
wire n_8605;
wire n_10358;
wire n_17593;
wire n_9944;
wire n_6998;
wire n_16158;
wire n_20105;
wire n_12338;
wire n_7615;
wire n_9605;
wire n_7591;
wire n_11404;
wire n_16488;
wire n_20584;
wire n_15994;
wire n_15685;
wire n_9788;
wire n_16273;
wire n_10785;
wire n_18262;
wire n_13872;
wire n_17646;
wire n_12341;
wire n_18389;
wire n_14475;
wire n_10815;
wire n_8784;
wire n_7382;
wire n_13955;
wire n_17708;
wire n_14400;
wire n_16904;
wire n_16725;
wire n_16432;
wire n_12085;
wire n_18190;
wire n_13554;
wire n_18421;
wire n_6780;
wire n_11582;
wire n_20083;
wire n_11705;
wire n_7673;
wire n_6830;
wire n_17391;
wire n_19782;
wire n_17682;
wire n_7282;
wire n_9968;
wire n_11474;
wire n_10657;
wire n_13595;
wire n_10687;
wire n_13283;
wire n_19543;
wire n_15615;
wire n_12110;
wire n_8363;
wire n_19445;
wire n_17802;
wire n_9669;
wire n_17775;
wire n_8282;
wire n_6510;
wire n_15972;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_17446;
wire n_18573;
wire n_14975;
wire n_7581;
wire n_6360;
wire n_17960;
wire n_15217;
wire n_13308;
wire n_19049;
wire n_9952;
wire n_15323;
wire n_12183;
wire n_19857;
wire n_9256;
wire n_10668;
wire n_14007;
wire n_7346;
wire n_13373;
wire n_7428;
wire n_12221;
wire n_9195;
wire n_16236;
wire n_17787;
wire n_7283;
wire n_6314;
wire n_10632;
wire n_18861;
wire n_9623;
wire n_6964;
wire n_19027;
wire n_19561;
wire n_18912;
wire n_19322;
wire n_16702;
wire n_11329;
wire n_6495;
wire n_17280;
wire n_9516;
wire n_13241;
wire n_16027;
wire n_8976;
wire n_17844;
wire n_18136;
wire n_10130;
wire n_11661;
wire n_9222;
wire n_8435;
wire n_8882;
wire n_16391;
wire n_15949;
wire n_10622;
wire n_19840;
wire n_6797;
wire n_15673;
wire n_14012;
wire n_8759;
wire n_16941;
wire n_7177;
wire n_13066;
wire n_13665;
wire n_12993;
wire n_19604;
wire n_11314;
wire n_17784;
wire n_15678;
wire n_8235;
wire n_13083;
wire n_19093;
wire n_16164;
wire n_6152;
wire n_16444;
wire n_9820;
wire n_14071;
wire n_12749;
wire n_8448;
wire n_12066;
wire n_6513;
wire n_15908;
wire n_11184;
wire n_11945;
wire n_11368;
wire n_6330;
wire n_17842;
wire n_19628;
wire n_8457;
wire n_19200;
wire n_18605;
wire n_18837;
wire n_9339;
wire n_14312;
wire n_9601;
wire n_15045;
wire n_11409;
wire n_18995;
wire n_20393;
wire n_18737;
wire n_12437;
wire n_10840;
wire n_6263;
wire n_10515;
wire n_15501;
wire n_6490;
wire n_15751;
wire n_11605;
wire n_10242;
wire n_10144;
wire n_9684;
wire n_15741;
wire n_16195;
wire n_14793;
wire n_18754;
wire n_13472;
wire n_15596;
wire n_18316;
wire n_15379;
wire n_16272;
wire n_14884;
wire n_8964;
wire n_16629;
wire n_9814;
wire n_14423;
wire n_16280;
wire n_16414;
wire n_13443;
wire n_14626;
wire n_20058;
wire n_8960;
wire n_19899;
wire n_15402;
wire n_20563;
wire n_18026;
wire n_8443;
wire n_7715;
wire n_8683;
wire n_18558;
wire n_6349;
wire n_10510;
wire n_15306;
wire n_15981;
wire n_19994;
wire n_16367;

CKINVDCx20_ASAP7_75t_R g6076 ( 
.A(n_3396),
.Y(n_6076)
);

INVx1_ASAP7_75t_SL g6077 ( 
.A(n_385),
.Y(n_6077)
);

CKINVDCx5p33_ASAP7_75t_R g6078 ( 
.A(n_4452),
.Y(n_6078)
);

CKINVDCx5p33_ASAP7_75t_R g6079 ( 
.A(n_3187),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_1373),
.Y(n_6080)
);

CKINVDCx5p33_ASAP7_75t_R g6081 ( 
.A(n_178),
.Y(n_6081)
);

CKINVDCx5p33_ASAP7_75t_R g6082 ( 
.A(n_5327),
.Y(n_6082)
);

CKINVDCx5p33_ASAP7_75t_R g6083 ( 
.A(n_1832),
.Y(n_6083)
);

CKINVDCx5p33_ASAP7_75t_R g6084 ( 
.A(n_615),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_4926),
.Y(n_6085)
);

CKINVDCx5p33_ASAP7_75t_R g6086 ( 
.A(n_5238),
.Y(n_6086)
);

BUFx6f_ASAP7_75t_L g6087 ( 
.A(n_2968),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_3627),
.Y(n_6088)
);

CKINVDCx20_ASAP7_75t_R g6089 ( 
.A(n_832),
.Y(n_6089)
);

BUFx6f_ASAP7_75t_L g6090 ( 
.A(n_1134),
.Y(n_6090)
);

CKINVDCx20_ASAP7_75t_R g6091 ( 
.A(n_2502),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_3675),
.Y(n_6092)
);

BUFx2_ASAP7_75t_L g6093 ( 
.A(n_4395),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_1627),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5277),
.Y(n_6095)
);

CKINVDCx5p33_ASAP7_75t_R g6096 ( 
.A(n_3348),
.Y(n_6096)
);

CKINVDCx5p33_ASAP7_75t_R g6097 ( 
.A(n_1304),
.Y(n_6097)
);

CKINVDCx5p33_ASAP7_75t_R g6098 ( 
.A(n_3414),
.Y(n_6098)
);

CKINVDCx5p33_ASAP7_75t_R g6099 ( 
.A(n_3802),
.Y(n_6099)
);

CKINVDCx20_ASAP7_75t_R g6100 ( 
.A(n_4429),
.Y(n_6100)
);

CKINVDCx5p33_ASAP7_75t_R g6101 ( 
.A(n_2918),
.Y(n_6101)
);

CKINVDCx5p33_ASAP7_75t_R g6102 ( 
.A(n_4929),
.Y(n_6102)
);

BUFx10_ASAP7_75t_L g6103 ( 
.A(n_1913),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_4434),
.Y(n_6104)
);

CKINVDCx5p33_ASAP7_75t_R g6105 ( 
.A(n_5335),
.Y(n_6105)
);

CKINVDCx5p33_ASAP7_75t_R g6106 ( 
.A(n_2726),
.Y(n_6106)
);

INVx1_ASAP7_75t_SL g6107 ( 
.A(n_3010),
.Y(n_6107)
);

BUFx6f_ASAP7_75t_L g6108 ( 
.A(n_675),
.Y(n_6108)
);

CKINVDCx5p33_ASAP7_75t_R g6109 ( 
.A(n_4247),
.Y(n_6109)
);

INVx2_ASAP7_75t_L g6110 ( 
.A(n_26),
.Y(n_6110)
);

CKINVDCx5p33_ASAP7_75t_R g6111 ( 
.A(n_924),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_992),
.Y(n_6112)
);

BUFx6f_ASAP7_75t_L g6113 ( 
.A(n_3874),
.Y(n_6113)
);

CKINVDCx5p33_ASAP7_75t_R g6114 ( 
.A(n_1131),
.Y(n_6114)
);

CKINVDCx5p33_ASAP7_75t_R g6115 ( 
.A(n_6055),
.Y(n_6115)
);

CKINVDCx20_ASAP7_75t_R g6116 ( 
.A(n_4570),
.Y(n_6116)
);

BUFx3_ASAP7_75t_L g6117 ( 
.A(n_5907),
.Y(n_6117)
);

CKINVDCx5p33_ASAP7_75t_R g6118 ( 
.A(n_3421),
.Y(n_6118)
);

CKINVDCx5p33_ASAP7_75t_R g6119 ( 
.A(n_5734),
.Y(n_6119)
);

CKINVDCx5p33_ASAP7_75t_R g6120 ( 
.A(n_6070),
.Y(n_6120)
);

BUFx2_ASAP7_75t_L g6121 ( 
.A(n_951),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5954),
.Y(n_6122)
);

CKINVDCx5p33_ASAP7_75t_R g6123 ( 
.A(n_4717),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_4365),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_2704),
.Y(n_6125)
);

CKINVDCx16_ASAP7_75t_R g6126 ( 
.A(n_1184),
.Y(n_6126)
);

INVx1_ASAP7_75t_SL g6127 ( 
.A(n_4472),
.Y(n_6127)
);

CKINVDCx5p33_ASAP7_75t_R g6128 ( 
.A(n_4579),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_4351),
.Y(n_6129)
);

BUFx5_ASAP7_75t_L g6130 ( 
.A(n_1610),
.Y(n_6130)
);

CKINVDCx5p33_ASAP7_75t_R g6131 ( 
.A(n_5704),
.Y(n_6131)
);

CKINVDCx5p33_ASAP7_75t_R g6132 ( 
.A(n_5442),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_1343),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_804),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_4186),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_4799),
.Y(n_6136)
);

CKINVDCx20_ASAP7_75t_R g6137 ( 
.A(n_253),
.Y(n_6137)
);

CKINVDCx5p33_ASAP7_75t_R g6138 ( 
.A(n_4612),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_859),
.Y(n_6139)
);

CKINVDCx5p33_ASAP7_75t_R g6140 ( 
.A(n_1507),
.Y(n_6140)
);

CKINVDCx5p33_ASAP7_75t_R g6141 ( 
.A(n_2795),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_1893),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_4500),
.Y(n_6143)
);

CKINVDCx5p33_ASAP7_75t_R g6144 ( 
.A(n_4451),
.Y(n_6144)
);

CKINVDCx5p33_ASAP7_75t_R g6145 ( 
.A(n_4143),
.Y(n_6145)
);

INVx1_ASAP7_75t_SL g6146 ( 
.A(n_3138),
.Y(n_6146)
);

CKINVDCx5p33_ASAP7_75t_R g6147 ( 
.A(n_1242),
.Y(n_6147)
);

CKINVDCx5p33_ASAP7_75t_R g6148 ( 
.A(n_4405),
.Y(n_6148)
);

CKINVDCx5p33_ASAP7_75t_R g6149 ( 
.A(n_4620),
.Y(n_6149)
);

CKINVDCx5p33_ASAP7_75t_R g6150 ( 
.A(n_1581),
.Y(n_6150)
);

BUFx6f_ASAP7_75t_L g6151 ( 
.A(n_1042),
.Y(n_6151)
);

CKINVDCx5p33_ASAP7_75t_R g6152 ( 
.A(n_4366),
.Y(n_6152)
);

CKINVDCx5p33_ASAP7_75t_R g6153 ( 
.A(n_5473),
.Y(n_6153)
);

CKINVDCx5p33_ASAP7_75t_R g6154 ( 
.A(n_4742),
.Y(n_6154)
);

CKINVDCx5p33_ASAP7_75t_R g6155 ( 
.A(n_5710),
.Y(n_6155)
);

CKINVDCx5p33_ASAP7_75t_R g6156 ( 
.A(n_2739),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5984),
.Y(n_6157)
);

CKINVDCx5p33_ASAP7_75t_R g6158 ( 
.A(n_2113),
.Y(n_6158)
);

CKINVDCx5p33_ASAP7_75t_R g6159 ( 
.A(n_4353),
.Y(n_6159)
);

INVx1_ASAP7_75t_SL g6160 ( 
.A(n_924),
.Y(n_6160)
);

CKINVDCx5p33_ASAP7_75t_R g6161 ( 
.A(n_232),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_4418),
.Y(n_6162)
);

CKINVDCx5p33_ASAP7_75t_R g6163 ( 
.A(n_5986),
.Y(n_6163)
);

CKINVDCx5p33_ASAP7_75t_R g6164 ( 
.A(n_1951),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_5831),
.Y(n_6165)
);

INVx1_ASAP7_75t_SL g6166 ( 
.A(n_2154),
.Y(n_6166)
);

BUFx6f_ASAP7_75t_L g6167 ( 
.A(n_4317),
.Y(n_6167)
);

CKINVDCx5p33_ASAP7_75t_R g6168 ( 
.A(n_1284),
.Y(n_6168)
);

CKINVDCx5p33_ASAP7_75t_R g6169 ( 
.A(n_4215),
.Y(n_6169)
);

CKINVDCx5p33_ASAP7_75t_R g6170 ( 
.A(n_4479),
.Y(n_6170)
);

CKINVDCx5p33_ASAP7_75t_R g6171 ( 
.A(n_2170),
.Y(n_6171)
);

INVx2_ASAP7_75t_SL g6172 ( 
.A(n_4490),
.Y(n_6172)
);

INVx2_ASAP7_75t_L g6173 ( 
.A(n_1485),
.Y(n_6173)
);

CKINVDCx5p33_ASAP7_75t_R g6174 ( 
.A(n_5086),
.Y(n_6174)
);

CKINVDCx5p33_ASAP7_75t_R g6175 ( 
.A(n_4381),
.Y(n_6175)
);

INVx1_ASAP7_75t_SL g6176 ( 
.A(n_5839),
.Y(n_6176)
);

BUFx5_ASAP7_75t_L g6177 ( 
.A(n_4357),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_6038),
.Y(n_6178)
);

CKINVDCx5p33_ASAP7_75t_R g6179 ( 
.A(n_2784),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_3895),
.Y(n_6180)
);

CKINVDCx5p33_ASAP7_75t_R g6181 ( 
.A(n_804),
.Y(n_6181)
);

CKINVDCx5p33_ASAP7_75t_R g6182 ( 
.A(n_4993),
.Y(n_6182)
);

CKINVDCx5p33_ASAP7_75t_R g6183 ( 
.A(n_195),
.Y(n_6183)
);

CKINVDCx5p33_ASAP7_75t_R g6184 ( 
.A(n_6059),
.Y(n_6184)
);

BUFx5_ASAP7_75t_L g6185 ( 
.A(n_6042),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_1494),
.Y(n_6186)
);

CKINVDCx5p33_ASAP7_75t_R g6187 ( 
.A(n_3413),
.Y(n_6187)
);

CKINVDCx5p33_ASAP7_75t_R g6188 ( 
.A(n_5209),
.Y(n_6188)
);

CKINVDCx20_ASAP7_75t_R g6189 ( 
.A(n_2410),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_1046),
.Y(n_6190)
);

CKINVDCx5p33_ASAP7_75t_R g6191 ( 
.A(n_560),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_3705),
.Y(n_6192)
);

BUFx6f_ASAP7_75t_L g6193 ( 
.A(n_5256),
.Y(n_6193)
);

CKINVDCx5p33_ASAP7_75t_R g6194 ( 
.A(n_244),
.Y(n_6194)
);

INVx2_ASAP7_75t_L g6195 ( 
.A(n_4841),
.Y(n_6195)
);

INVxp67_ASAP7_75t_SL g6196 ( 
.A(n_2782),
.Y(n_6196)
);

CKINVDCx5p33_ASAP7_75t_R g6197 ( 
.A(n_3865),
.Y(n_6197)
);

CKINVDCx5p33_ASAP7_75t_R g6198 ( 
.A(n_2221),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_1221),
.Y(n_6199)
);

CKINVDCx5p33_ASAP7_75t_R g6200 ( 
.A(n_4535),
.Y(n_6200)
);

INVx2_ASAP7_75t_SL g6201 ( 
.A(n_5700),
.Y(n_6201)
);

CKINVDCx5p33_ASAP7_75t_R g6202 ( 
.A(n_2850),
.Y(n_6202)
);

CKINVDCx20_ASAP7_75t_R g6203 ( 
.A(n_4852),
.Y(n_6203)
);

CKINVDCx20_ASAP7_75t_R g6204 ( 
.A(n_611),
.Y(n_6204)
);

CKINVDCx20_ASAP7_75t_R g6205 ( 
.A(n_4623),
.Y(n_6205)
);

CKINVDCx5p33_ASAP7_75t_R g6206 ( 
.A(n_4400),
.Y(n_6206)
);

CKINVDCx5p33_ASAP7_75t_R g6207 ( 
.A(n_4751),
.Y(n_6207)
);

CKINVDCx5p33_ASAP7_75t_R g6208 ( 
.A(n_2613),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_5705),
.Y(n_6209)
);

CKINVDCx5p33_ASAP7_75t_R g6210 ( 
.A(n_903),
.Y(n_6210)
);

BUFx10_ASAP7_75t_L g6211 ( 
.A(n_1422),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_886),
.Y(n_6212)
);

CKINVDCx5p33_ASAP7_75t_R g6213 ( 
.A(n_4475),
.Y(n_6213)
);

CKINVDCx5p33_ASAP7_75t_R g6214 ( 
.A(n_5241),
.Y(n_6214)
);

CKINVDCx5p33_ASAP7_75t_R g6215 ( 
.A(n_4462),
.Y(n_6215)
);

CKINVDCx5p33_ASAP7_75t_R g6216 ( 
.A(n_4878),
.Y(n_6216)
);

CKINVDCx5p33_ASAP7_75t_R g6217 ( 
.A(n_4402),
.Y(n_6217)
);

CKINVDCx5p33_ASAP7_75t_R g6218 ( 
.A(n_6037),
.Y(n_6218)
);

CKINVDCx5p33_ASAP7_75t_R g6219 ( 
.A(n_1023),
.Y(n_6219)
);

CKINVDCx5p33_ASAP7_75t_R g6220 ( 
.A(n_5272),
.Y(n_6220)
);

INVx1_ASAP7_75t_L g6221 ( 
.A(n_5680),
.Y(n_6221)
);

CKINVDCx5p33_ASAP7_75t_R g6222 ( 
.A(n_4475),
.Y(n_6222)
);

CKINVDCx5p33_ASAP7_75t_R g6223 ( 
.A(n_4705),
.Y(n_6223)
);

CKINVDCx5p33_ASAP7_75t_R g6224 ( 
.A(n_2909),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_3694),
.Y(n_6225)
);

CKINVDCx5p33_ASAP7_75t_R g6226 ( 
.A(n_4187),
.Y(n_6226)
);

INVxp67_ASAP7_75t_L g6227 ( 
.A(n_4539),
.Y(n_6227)
);

CKINVDCx20_ASAP7_75t_R g6228 ( 
.A(n_769),
.Y(n_6228)
);

CKINVDCx5p33_ASAP7_75t_R g6229 ( 
.A(n_2162),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5249),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5167),
.Y(n_6231)
);

CKINVDCx5p33_ASAP7_75t_R g6232 ( 
.A(n_4521),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_4700),
.Y(n_6233)
);

CKINVDCx20_ASAP7_75t_R g6234 ( 
.A(n_4566),
.Y(n_6234)
);

CKINVDCx5p33_ASAP7_75t_R g6235 ( 
.A(n_4670),
.Y(n_6235)
);

CKINVDCx5p33_ASAP7_75t_R g6236 ( 
.A(n_5542),
.Y(n_6236)
);

INVx1_ASAP7_75t_SL g6237 ( 
.A(n_1037),
.Y(n_6237)
);

CKINVDCx5p33_ASAP7_75t_R g6238 ( 
.A(n_43),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_3601),
.Y(n_6239)
);

CKINVDCx5p33_ASAP7_75t_R g6240 ( 
.A(n_2515),
.Y(n_6240)
);

BUFx5_ASAP7_75t_L g6241 ( 
.A(n_2939),
.Y(n_6241)
);

INVx1_ASAP7_75t_L g6242 ( 
.A(n_964),
.Y(n_6242)
);

CKINVDCx5p33_ASAP7_75t_R g6243 ( 
.A(n_1454),
.Y(n_6243)
);

CKINVDCx5p33_ASAP7_75t_R g6244 ( 
.A(n_4414),
.Y(n_6244)
);

INVx2_ASAP7_75t_L g6245 ( 
.A(n_3503),
.Y(n_6245)
);

BUFx3_ASAP7_75t_L g6246 ( 
.A(n_1418),
.Y(n_6246)
);

INVx2_ASAP7_75t_L g6247 ( 
.A(n_1050),
.Y(n_6247)
);

CKINVDCx5p33_ASAP7_75t_R g6248 ( 
.A(n_19),
.Y(n_6248)
);

CKINVDCx5p33_ASAP7_75t_R g6249 ( 
.A(n_5259),
.Y(n_6249)
);

CKINVDCx20_ASAP7_75t_R g6250 ( 
.A(n_2903),
.Y(n_6250)
);

CKINVDCx11_ASAP7_75t_R g6251 ( 
.A(n_4503),
.Y(n_6251)
);

CKINVDCx5p33_ASAP7_75t_R g6252 ( 
.A(n_2079),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_36),
.Y(n_6253)
);

INVx1_ASAP7_75t_SL g6254 ( 
.A(n_593),
.Y(n_6254)
);

CKINVDCx5p33_ASAP7_75t_R g6255 ( 
.A(n_4849),
.Y(n_6255)
);

CKINVDCx5p33_ASAP7_75t_R g6256 ( 
.A(n_2809),
.Y(n_6256)
);

INVx1_ASAP7_75t_SL g6257 ( 
.A(n_5647),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_2953),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_3507),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_468),
.Y(n_6260)
);

INVx1_ASAP7_75t_L g6261 ( 
.A(n_4403),
.Y(n_6261)
);

CKINVDCx5p33_ASAP7_75t_R g6262 ( 
.A(n_3982),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_4706),
.Y(n_6263)
);

CKINVDCx16_ASAP7_75t_R g6264 ( 
.A(n_4983),
.Y(n_6264)
);

CKINVDCx5p33_ASAP7_75t_R g6265 ( 
.A(n_5388),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_4455),
.Y(n_6266)
);

BUFx6f_ASAP7_75t_L g6267 ( 
.A(n_1212),
.Y(n_6267)
);

CKINVDCx5p33_ASAP7_75t_R g6268 ( 
.A(n_4444),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_6054),
.Y(n_6269)
);

BUFx5_ASAP7_75t_L g6270 ( 
.A(n_2682),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_1802),
.Y(n_6271)
);

CKINVDCx5p33_ASAP7_75t_R g6272 ( 
.A(n_2474),
.Y(n_6272)
);

CKINVDCx5p33_ASAP7_75t_R g6273 ( 
.A(n_3765),
.Y(n_6273)
);

CKINVDCx5p33_ASAP7_75t_R g6274 ( 
.A(n_3253),
.Y(n_6274)
);

CKINVDCx5p33_ASAP7_75t_R g6275 ( 
.A(n_1823),
.Y(n_6275)
);

INVx1_ASAP7_75t_L g6276 ( 
.A(n_1381),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_4147),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_1971),
.Y(n_6278)
);

CKINVDCx20_ASAP7_75t_R g6279 ( 
.A(n_4359),
.Y(n_6279)
);

CKINVDCx5p33_ASAP7_75t_R g6280 ( 
.A(n_3800),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_2774),
.Y(n_6281)
);

CKINVDCx5p33_ASAP7_75t_R g6282 ( 
.A(n_954),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_5834),
.Y(n_6283)
);

CKINVDCx5p33_ASAP7_75t_R g6284 ( 
.A(n_970),
.Y(n_6284)
);

BUFx10_ASAP7_75t_L g6285 ( 
.A(n_88),
.Y(n_6285)
);

CKINVDCx5p33_ASAP7_75t_R g6286 ( 
.A(n_4663),
.Y(n_6286)
);

CKINVDCx20_ASAP7_75t_R g6287 ( 
.A(n_4545),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_4148),
.Y(n_6288)
);

INVx2_ASAP7_75t_L g6289 ( 
.A(n_42),
.Y(n_6289)
);

CKINVDCx5p33_ASAP7_75t_R g6290 ( 
.A(n_2572),
.Y(n_6290)
);

CKINVDCx5p33_ASAP7_75t_R g6291 ( 
.A(n_815),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_498),
.Y(n_6292)
);

CKINVDCx5p33_ASAP7_75t_R g6293 ( 
.A(n_2804),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_72),
.Y(n_6294)
);

CKINVDCx5p33_ASAP7_75t_R g6295 ( 
.A(n_198),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_3595),
.Y(n_6296)
);

CKINVDCx5p33_ASAP7_75t_R g6297 ( 
.A(n_3561),
.Y(n_6297)
);

CKINVDCx5p33_ASAP7_75t_R g6298 ( 
.A(n_5780),
.Y(n_6298)
);

CKINVDCx20_ASAP7_75t_R g6299 ( 
.A(n_2748),
.Y(n_6299)
);

CKINVDCx5p33_ASAP7_75t_R g6300 ( 
.A(n_2903),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5151),
.Y(n_6301)
);

CKINVDCx5p33_ASAP7_75t_R g6302 ( 
.A(n_382),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_6057),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_3815),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_894),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_1641),
.Y(n_6306)
);

CKINVDCx5p33_ASAP7_75t_R g6307 ( 
.A(n_4014),
.Y(n_6307)
);

CKINVDCx5p33_ASAP7_75t_R g6308 ( 
.A(n_941),
.Y(n_6308)
);

BUFx5_ASAP7_75t_L g6309 ( 
.A(n_3202),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_869),
.Y(n_6310)
);

CKINVDCx5p33_ASAP7_75t_R g6311 ( 
.A(n_4909),
.Y(n_6311)
);

BUFx10_ASAP7_75t_L g6312 ( 
.A(n_5678),
.Y(n_6312)
);

BUFx3_ASAP7_75t_L g6313 ( 
.A(n_5281),
.Y(n_6313)
);

INVx2_ASAP7_75t_L g6314 ( 
.A(n_342),
.Y(n_6314)
);

CKINVDCx5p33_ASAP7_75t_R g6315 ( 
.A(n_5610),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_771),
.Y(n_6316)
);

CKINVDCx5p33_ASAP7_75t_R g6317 ( 
.A(n_4648),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_10),
.Y(n_6318)
);

CKINVDCx20_ASAP7_75t_R g6319 ( 
.A(n_5382),
.Y(n_6319)
);

CKINVDCx5p33_ASAP7_75t_R g6320 ( 
.A(n_3581),
.Y(n_6320)
);

CKINVDCx5p33_ASAP7_75t_R g6321 ( 
.A(n_5471),
.Y(n_6321)
);

HB1xp67_ASAP7_75t_L g6322 ( 
.A(n_1725),
.Y(n_6322)
);

CKINVDCx5p33_ASAP7_75t_R g6323 ( 
.A(n_2734),
.Y(n_6323)
);

BUFx2_ASAP7_75t_L g6324 ( 
.A(n_1916),
.Y(n_6324)
);

CKINVDCx5p33_ASAP7_75t_R g6325 ( 
.A(n_3894),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_730),
.Y(n_6326)
);

CKINVDCx5p33_ASAP7_75t_R g6327 ( 
.A(n_6073),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_2149),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_4085),
.Y(n_6329)
);

BUFx6f_ASAP7_75t_L g6330 ( 
.A(n_317),
.Y(n_6330)
);

CKINVDCx20_ASAP7_75t_R g6331 ( 
.A(n_2367),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_4457),
.Y(n_6332)
);

BUFx8_ASAP7_75t_SL g6333 ( 
.A(n_5144),
.Y(n_6333)
);

BUFx6f_ASAP7_75t_L g6334 ( 
.A(n_6040),
.Y(n_6334)
);

CKINVDCx5p33_ASAP7_75t_R g6335 ( 
.A(n_1742),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_5075),
.Y(n_6336)
);

CKINVDCx5p33_ASAP7_75t_R g6337 ( 
.A(n_769),
.Y(n_6337)
);

CKINVDCx5p33_ASAP7_75t_R g6338 ( 
.A(n_4392),
.Y(n_6338)
);

CKINVDCx5p33_ASAP7_75t_R g6339 ( 
.A(n_2246),
.Y(n_6339)
);

CKINVDCx5p33_ASAP7_75t_R g6340 ( 
.A(n_4059),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_1584),
.Y(n_6341)
);

CKINVDCx5p33_ASAP7_75t_R g6342 ( 
.A(n_3730),
.Y(n_6342)
);

CKINVDCx20_ASAP7_75t_R g6343 ( 
.A(n_4497),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_2864),
.Y(n_6344)
);

CKINVDCx5p33_ASAP7_75t_R g6345 ( 
.A(n_3520),
.Y(n_6345)
);

INVx1_ASAP7_75t_L g6346 ( 
.A(n_997),
.Y(n_6346)
);

BUFx3_ASAP7_75t_L g6347 ( 
.A(n_2306),
.Y(n_6347)
);

CKINVDCx5p33_ASAP7_75t_R g6348 ( 
.A(n_665),
.Y(n_6348)
);

INVx1_ASAP7_75t_L g6349 ( 
.A(n_2858),
.Y(n_6349)
);

CKINVDCx5p33_ASAP7_75t_R g6350 ( 
.A(n_5672),
.Y(n_6350)
);

CKINVDCx5p33_ASAP7_75t_R g6351 ( 
.A(n_4374),
.Y(n_6351)
);

CKINVDCx5p33_ASAP7_75t_R g6352 ( 
.A(n_2853),
.Y(n_6352)
);

CKINVDCx5p33_ASAP7_75t_R g6353 ( 
.A(n_5854),
.Y(n_6353)
);

INVx1_ASAP7_75t_L g6354 ( 
.A(n_5440),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_1503),
.Y(n_6355)
);

CKINVDCx5p33_ASAP7_75t_R g6356 ( 
.A(n_4563),
.Y(n_6356)
);

BUFx6f_ASAP7_75t_L g6357 ( 
.A(n_3909),
.Y(n_6357)
);

CKINVDCx5p33_ASAP7_75t_R g6358 ( 
.A(n_3290),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_1322),
.Y(n_6359)
);

CKINVDCx20_ASAP7_75t_R g6360 ( 
.A(n_2339),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_491),
.Y(n_6361)
);

CKINVDCx5p33_ASAP7_75t_R g6362 ( 
.A(n_5460),
.Y(n_6362)
);

INVx2_ASAP7_75t_L g6363 ( 
.A(n_4529),
.Y(n_6363)
);

CKINVDCx5p33_ASAP7_75t_R g6364 ( 
.A(n_3786),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_431),
.Y(n_6365)
);

CKINVDCx5p33_ASAP7_75t_R g6366 ( 
.A(n_4581),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_1433),
.Y(n_6367)
);

CKINVDCx5p33_ASAP7_75t_R g6368 ( 
.A(n_5882),
.Y(n_6368)
);

CKINVDCx5p33_ASAP7_75t_R g6369 ( 
.A(n_229),
.Y(n_6369)
);

CKINVDCx5p33_ASAP7_75t_R g6370 ( 
.A(n_830),
.Y(n_6370)
);

CKINVDCx5p33_ASAP7_75t_R g6371 ( 
.A(n_3580),
.Y(n_6371)
);

CKINVDCx5p33_ASAP7_75t_R g6372 ( 
.A(n_3608),
.Y(n_6372)
);

BUFx6f_ASAP7_75t_L g6373 ( 
.A(n_4658),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_658),
.Y(n_6374)
);

CKINVDCx5p33_ASAP7_75t_R g6375 ( 
.A(n_1056),
.Y(n_6375)
);

CKINVDCx5p33_ASAP7_75t_R g6376 ( 
.A(n_749),
.Y(n_6376)
);

CKINVDCx5p33_ASAP7_75t_R g6377 ( 
.A(n_1053),
.Y(n_6377)
);

CKINVDCx5p33_ASAP7_75t_R g6378 ( 
.A(n_2628),
.Y(n_6378)
);

CKINVDCx5p33_ASAP7_75t_R g6379 ( 
.A(n_779),
.Y(n_6379)
);

CKINVDCx5p33_ASAP7_75t_R g6380 ( 
.A(n_68),
.Y(n_6380)
);

BUFx5_ASAP7_75t_L g6381 ( 
.A(n_4454),
.Y(n_6381)
);

BUFx3_ASAP7_75t_L g6382 ( 
.A(n_4177),
.Y(n_6382)
);

BUFx3_ASAP7_75t_L g6383 ( 
.A(n_1653),
.Y(n_6383)
);

INVx1_ASAP7_75t_L g6384 ( 
.A(n_3453),
.Y(n_6384)
);

CKINVDCx5p33_ASAP7_75t_R g6385 ( 
.A(n_5684),
.Y(n_6385)
);

CKINVDCx5p33_ASAP7_75t_R g6386 ( 
.A(n_1448),
.Y(n_6386)
);

CKINVDCx5p33_ASAP7_75t_R g6387 ( 
.A(n_3893),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5221),
.Y(n_6388)
);

CKINVDCx5p33_ASAP7_75t_R g6389 ( 
.A(n_2935),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_124),
.Y(n_6390)
);

CKINVDCx5p33_ASAP7_75t_R g6391 ( 
.A(n_4765),
.Y(n_6391)
);

CKINVDCx5p33_ASAP7_75t_R g6392 ( 
.A(n_1060),
.Y(n_6392)
);

CKINVDCx5p33_ASAP7_75t_R g6393 ( 
.A(n_3161),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_4419),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_1257),
.Y(n_6395)
);

CKINVDCx5p33_ASAP7_75t_R g6396 ( 
.A(n_971),
.Y(n_6396)
);

INVx1_ASAP7_75t_SL g6397 ( 
.A(n_881),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_4438),
.Y(n_6398)
);

INVx2_ASAP7_75t_L g6399 ( 
.A(n_131),
.Y(n_6399)
);

HB1xp67_ASAP7_75t_L g6400 ( 
.A(n_4522),
.Y(n_6400)
);

CKINVDCx5p33_ASAP7_75t_R g6401 ( 
.A(n_1464),
.Y(n_6401)
);

CKINVDCx14_ASAP7_75t_R g6402 ( 
.A(n_264),
.Y(n_6402)
);

CKINVDCx5p33_ASAP7_75t_R g6403 ( 
.A(n_3646),
.Y(n_6403)
);

CKINVDCx5p33_ASAP7_75t_R g6404 ( 
.A(n_3003),
.Y(n_6404)
);

CKINVDCx5p33_ASAP7_75t_R g6405 ( 
.A(n_4523),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_3596),
.Y(n_6406)
);

CKINVDCx5p33_ASAP7_75t_R g6407 ( 
.A(n_6067),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_1509),
.Y(n_6408)
);

CKINVDCx5p33_ASAP7_75t_R g6409 ( 
.A(n_3170),
.Y(n_6409)
);

CKINVDCx5p33_ASAP7_75t_R g6410 ( 
.A(n_1777),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_5694),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_1780),
.Y(n_6412)
);

BUFx10_ASAP7_75t_L g6413 ( 
.A(n_3835),
.Y(n_6413)
);

INVx1_ASAP7_75t_SL g6414 ( 
.A(n_2507),
.Y(n_6414)
);

CKINVDCx16_ASAP7_75t_R g6415 ( 
.A(n_3875),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_3287),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_1114),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_694),
.Y(n_6418)
);

CKINVDCx5p33_ASAP7_75t_R g6419 ( 
.A(n_1170),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_2041),
.Y(n_6420)
);

CKINVDCx5p33_ASAP7_75t_R g6421 ( 
.A(n_3259),
.Y(n_6421)
);

CKINVDCx5p33_ASAP7_75t_R g6422 ( 
.A(n_4443),
.Y(n_6422)
);

INVxp67_ASAP7_75t_L g6423 ( 
.A(n_2227),
.Y(n_6423)
);

HB1xp67_ASAP7_75t_L g6424 ( 
.A(n_2108),
.Y(n_6424)
);

CKINVDCx5p33_ASAP7_75t_R g6425 ( 
.A(n_4358),
.Y(n_6425)
);

CKINVDCx5p33_ASAP7_75t_R g6426 ( 
.A(n_4439),
.Y(n_6426)
);

CKINVDCx5p33_ASAP7_75t_R g6427 ( 
.A(n_1178),
.Y(n_6427)
);

CKINVDCx20_ASAP7_75t_R g6428 ( 
.A(n_4279),
.Y(n_6428)
);

CKINVDCx5p33_ASAP7_75t_R g6429 ( 
.A(n_1853),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_5632),
.Y(n_6430)
);

INVx1_ASAP7_75t_SL g6431 ( 
.A(n_4546),
.Y(n_6431)
);

INVx2_ASAP7_75t_L g6432 ( 
.A(n_3298),
.Y(n_6432)
);

CKINVDCx5p33_ASAP7_75t_R g6433 ( 
.A(n_1993),
.Y(n_6433)
);

CKINVDCx5p33_ASAP7_75t_R g6434 ( 
.A(n_6075),
.Y(n_6434)
);

CKINVDCx5p33_ASAP7_75t_R g6435 ( 
.A(n_485),
.Y(n_6435)
);

CKINVDCx5p33_ASAP7_75t_R g6436 ( 
.A(n_5416),
.Y(n_6436)
);

INVxp33_ASAP7_75t_R g6437 ( 
.A(n_1364),
.Y(n_6437)
);

CKINVDCx16_ASAP7_75t_R g6438 ( 
.A(n_2626),
.Y(n_6438)
);

INVx1_ASAP7_75t_SL g6439 ( 
.A(n_3071),
.Y(n_6439)
);

CKINVDCx5p33_ASAP7_75t_R g6440 ( 
.A(n_4369),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_4300),
.Y(n_6441)
);

CKINVDCx5p33_ASAP7_75t_R g6442 ( 
.A(n_5682),
.Y(n_6442)
);

CKINVDCx5p33_ASAP7_75t_R g6443 ( 
.A(n_3109),
.Y(n_6443)
);

CKINVDCx20_ASAP7_75t_R g6444 ( 
.A(n_1176),
.Y(n_6444)
);

INVxp67_ASAP7_75t_L g6445 ( 
.A(n_112),
.Y(n_6445)
);

CKINVDCx5p33_ASAP7_75t_R g6446 ( 
.A(n_4506),
.Y(n_6446)
);

INVx2_ASAP7_75t_L g6447 ( 
.A(n_4542),
.Y(n_6447)
);

CKINVDCx5p33_ASAP7_75t_R g6448 ( 
.A(n_5519),
.Y(n_6448)
);

BUFx8_ASAP7_75t_SL g6449 ( 
.A(n_942),
.Y(n_6449)
);

CKINVDCx5p33_ASAP7_75t_R g6450 ( 
.A(n_4404),
.Y(n_6450)
);

INVx2_ASAP7_75t_L g6451 ( 
.A(n_105),
.Y(n_6451)
);

INVx2_ASAP7_75t_SL g6452 ( 
.A(n_990),
.Y(n_6452)
);

CKINVDCx5p33_ASAP7_75t_R g6453 ( 
.A(n_5692),
.Y(n_6453)
);

BUFx3_ASAP7_75t_L g6454 ( 
.A(n_5091),
.Y(n_6454)
);

CKINVDCx5p33_ASAP7_75t_R g6455 ( 
.A(n_2534),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_2633),
.Y(n_6456)
);

CKINVDCx20_ASAP7_75t_R g6457 ( 
.A(n_2266),
.Y(n_6457)
);

CKINVDCx5p33_ASAP7_75t_R g6458 ( 
.A(n_2328),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_4382),
.Y(n_6459)
);

CKINVDCx5p33_ASAP7_75t_R g6460 ( 
.A(n_6058),
.Y(n_6460)
);

CKINVDCx5p33_ASAP7_75t_R g6461 ( 
.A(n_1801),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_4478),
.Y(n_6462)
);

CKINVDCx5p33_ASAP7_75t_R g6463 ( 
.A(n_4423),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_5182),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_3673),
.Y(n_6465)
);

CKINVDCx20_ASAP7_75t_R g6466 ( 
.A(n_4674),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_1216),
.Y(n_6467)
);

CKINVDCx5p33_ASAP7_75t_R g6468 ( 
.A(n_5072),
.Y(n_6468)
);

INVx2_ASAP7_75t_SL g6469 ( 
.A(n_3640),
.Y(n_6469)
);

BUFx3_ASAP7_75t_L g6470 ( 
.A(n_1564),
.Y(n_6470)
);

INVx1_ASAP7_75t_SL g6471 ( 
.A(n_5747),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_846),
.Y(n_6472)
);

CKINVDCx16_ASAP7_75t_R g6473 ( 
.A(n_2299),
.Y(n_6473)
);

INVx2_ASAP7_75t_L g6474 ( 
.A(n_4449),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_2727),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_3537),
.Y(n_6476)
);

CKINVDCx14_ASAP7_75t_R g6477 ( 
.A(n_5673),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_342),
.Y(n_6478)
);

CKINVDCx20_ASAP7_75t_R g6479 ( 
.A(n_4534),
.Y(n_6479)
);

CKINVDCx5p33_ASAP7_75t_R g6480 ( 
.A(n_4299),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_3768),
.Y(n_6481)
);

CKINVDCx5p33_ASAP7_75t_R g6482 ( 
.A(n_3109),
.Y(n_6482)
);

CKINVDCx5p33_ASAP7_75t_R g6483 ( 
.A(n_5466),
.Y(n_6483)
);

BUFx8_ASAP7_75t_SL g6484 ( 
.A(n_289),
.Y(n_6484)
);

CKINVDCx5p33_ASAP7_75t_R g6485 ( 
.A(n_1584),
.Y(n_6485)
);

CKINVDCx5p33_ASAP7_75t_R g6486 ( 
.A(n_850),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_1722),
.Y(n_6487)
);

CKINVDCx5p33_ASAP7_75t_R g6488 ( 
.A(n_1694),
.Y(n_6488)
);

CKINVDCx5p33_ASAP7_75t_R g6489 ( 
.A(n_5280),
.Y(n_6489)
);

CKINVDCx14_ASAP7_75t_R g6490 ( 
.A(n_4205),
.Y(n_6490)
);

CKINVDCx5p33_ASAP7_75t_R g6491 ( 
.A(n_351),
.Y(n_6491)
);

CKINVDCx5p33_ASAP7_75t_R g6492 ( 
.A(n_2655),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_3941),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_4853),
.Y(n_6494)
);

HB1xp67_ASAP7_75t_L g6495 ( 
.A(n_1221),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_5828),
.Y(n_6496)
);

CKINVDCx5p33_ASAP7_75t_R g6497 ( 
.A(n_1268),
.Y(n_6497)
);

CKINVDCx14_ASAP7_75t_R g6498 ( 
.A(n_6072),
.Y(n_6498)
);

CKINVDCx5p33_ASAP7_75t_R g6499 ( 
.A(n_4262),
.Y(n_6499)
);

INVx2_ASAP7_75t_SL g6500 ( 
.A(n_5732),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_175),
.Y(n_6501)
);

CKINVDCx20_ASAP7_75t_R g6502 ( 
.A(n_4639),
.Y(n_6502)
);

CKINVDCx5p33_ASAP7_75t_R g6503 ( 
.A(n_1369),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_2024),
.Y(n_6504)
);

CKINVDCx5p33_ASAP7_75t_R g6505 ( 
.A(n_681),
.Y(n_6505)
);

CKINVDCx5p33_ASAP7_75t_R g6506 ( 
.A(n_3322),
.Y(n_6506)
);

INVx1_ASAP7_75t_SL g6507 ( 
.A(n_13),
.Y(n_6507)
);

CKINVDCx5p33_ASAP7_75t_R g6508 ( 
.A(n_2642),
.Y(n_6508)
);

INVx1_ASAP7_75t_L g6509 ( 
.A(n_4768),
.Y(n_6509)
);

CKINVDCx5p33_ASAP7_75t_R g6510 ( 
.A(n_1948),
.Y(n_6510)
);

INVxp67_ASAP7_75t_L g6511 ( 
.A(n_9),
.Y(n_6511)
);

CKINVDCx5p33_ASAP7_75t_R g6512 ( 
.A(n_569),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_5608),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_5926),
.Y(n_6514)
);

CKINVDCx5p33_ASAP7_75t_R g6515 ( 
.A(n_591),
.Y(n_6515)
);

CKINVDCx5p33_ASAP7_75t_R g6516 ( 
.A(n_4131),
.Y(n_6516)
);

BUFx10_ASAP7_75t_L g6517 ( 
.A(n_5573),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_4477),
.Y(n_6518)
);

INVx1_ASAP7_75t_L g6519 ( 
.A(n_4433),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_2583),
.Y(n_6520)
);

CKINVDCx20_ASAP7_75t_R g6521 ( 
.A(n_4501),
.Y(n_6521)
);

CKINVDCx5p33_ASAP7_75t_R g6522 ( 
.A(n_5087),
.Y(n_6522)
);

CKINVDCx5p33_ASAP7_75t_R g6523 ( 
.A(n_4446),
.Y(n_6523)
);

CKINVDCx5p33_ASAP7_75t_R g6524 ( 
.A(n_2210),
.Y(n_6524)
);

CKINVDCx5p33_ASAP7_75t_R g6525 ( 
.A(n_1028),
.Y(n_6525)
);

CKINVDCx5p33_ASAP7_75t_R g6526 ( 
.A(n_1025),
.Y(n_6526)
);

CKINVDCx5p33_ASAP7_75t_R g6527 ( 
.A(n_2359),
.Y(n_6527)
);

CKINVDCx5p33_ASAP7_75t_R g6528 ( 
.A(n_2144),
.Y(n_6528)
);

CKINVDCx5p33_ASAP7_75t_R g6529 ( 
.A(n_4394),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_1980),
.Y(n_6530)
);

CKINVDCx5p33_ASAP7_75t_R g6531 ( 
.A(n_4375),
.Y(n_6531)
);

CKINVDCx5p33_ASAP7_75t_R g6532 ( 
.A(n_4476),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_4510),
.Y(n_6533)
);

CKINVDCx5p33_ASAP7_75t_R g6534 ( 
.A(n_4736),
.Y(n_6534)
);

BUFx6f_ASAP7_75t_L g6535 ( 
.A(n_4413),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_699),
.Y(n_6536)
);

INVx4_ASAP7_75t_R g6537 ( 
.A(n_4601),
.Y(n_6537)
);

INVx1_ASAP7_75t_SL g6538 ( 
.A(n_5216),
.Y(n_6538)
);

CKINVDCx5p33_ASAP7_75t_R g6539 ( 
.A(n_1575),
.Y(n_6539)
);

CKINVDCx5p33_ASAP7_75t_R g6540 ( 
.A(n_3626),
.Y(n_6540)
);

INVxp67_ASAP7_75t_L g6541 ( 
.A(n_1905),
.Y(n_6541)
);

CKINVDCx5p33_ASAP7_75t_R g6542 ( 
.A(n_5570),
.Y(n_6542)
);

CKINVDCx5p33_ASAP7_75t_R g6543 ( 
.A(n_854),
.Y(n_6543)
);

CKINVDCx5p33_ASAP7_75t_R g6544 ( 
.A(n_4517),
.Y(n_6544)
);

CKINVDCx20_ASAP7_75t_R g6545 ( 
.A(n_2949),
.Y(n_6545)
);

INVx2_ASAP7_75t_SL g6546 ( 
.A(n_1690),
.Y(n_6546)
);

CKINVDCx5p33_ASAP7_75t_R g6547 ( 
.A(n_2250),
.Y(n_6547)
);

CKINVDCx5p33_ASAP7_75t_R g6548 ( 
.A(n_4370),
.Y(n_6548)
);

CKINVDCx16_ASAP7_75t_R g6549 ( 
.A(n_2310),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_6056),
.Y(n_6550)
);

CKINVDCx20_ASAP7_75t_R g6551 ( 
.A(n_876),
.Y(n_6551)
);

CKINVDCx16_ASAP7_75t_R g6552 ( 
.A(n_3106),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_5399),
.Y(n_6553)
);

CKINVDCx5p33_ASAP7_75t_R g6554 ( 
.A(n_2507),
.Y(n_6554)
);

INVx1_ASAP7_75t_L g6555 ( 
.A(n_2823),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_3076),
.Y(n_6556)
);

CKINVDCx5p33_ASAP7_75t_R g6557 ( 
.A(n_4485),
.Y(n_6557)
);

BUFx10_ASAP7_75t_L g6558 ( 
.A(n_2847),
.Y(n_6558)
);

INVx1_ASAP7_75t_L g6559 ( 
.A(n_4149),
.Y(n_6559)
);

CKINVDCx5p33_ASAP7_75t_R g6560 ( 
.A(n_4908),
.Y(n_6560)
);

INVx1_ASAP7_75t_L g6561 ( 
.A(n_5605),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_706),
.Y(n_6562)
);

CKINVDCx5p33_ASAP7_75t_R g6563 ( 
.A(n_4122),
.Y(n_6563)
);

CKINVDCx5p33_ASAP7_75t_R g6564 ( 
.A(n_4928),
.Y(n_6564)
);

INVx1_ASAP7_75t_L g6565 ( 
.A(n_2328),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_352),
.Y(n_6566)
);

INVx2_ASAP7_75t_L g6567 ( 
.A(n_4778),
.Y(n_6567)
);

BUFx3_ASAP7_75t_L g6568 ( 
.A(n_1844),
.Y(n_6568)
);

CKINVDCx5p33_ASAP7_75t_R g6569 ( 
.A(n_4482),
.Y(n_6569)
);

CKINVDCx5p33_ASAP7_75t_R g6570 ( 
.A(n_5522),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_3539),
.Y(n_6571)
);

CKINVDCx5p33_ASAP7_75t_R g6572 ( 
.A(n_6043),
.Y(n_6572)
);

BUFx3_ASAP7_75t_L g6573 ( 
.A(n_161),
.Y(n_6573)
);

CKINVDCx5p33_ASAP7_75t_R g6574 ( 
.A(n_2421),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_314),
.Y(n_6575)
);

CKINVDCx5p33_ASAP7_75t_R g6576 ( 
.A(n_1708),
.Y(n_6576)
);

CKINVDCx5p33_ASAP7_75t_R g6577 ( 
.A(n_3619),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_3697),
.Y(n_6578)
);

CKINVDCx5p33_ASAP7_75t_R g6579 ( 
.A(n_860),
.Y(n_6579)
);

CKINVDCx20_ASAP7_75t_R g6580 ( 
.A(n_1262),
.Y(n_6580)
);

CKINVDCx5p33_ASAP7_75t_R g6581 ( 
.A(n_3988),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_3398),
.Y(n_6582)
);

CKINVDCx20_ASAP7_75t_R g6583 ( 
.A(n_5127),
.Y(n_6583)
);

CKINVDCx20_ASAP7_75t_R g6584 ( 
.A(n_3324),
.Y(n_6584)
);

INVx1_ASAP7_75t_L g6585 ( 
.A(n_4364),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_281),
.Y(n_6586)
);

INVx2_ASAP7_75t_SL g6587 ( 
.A(n_4806),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_2143),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_1327),
.Y(n_6589)
);

CKINVDCx5p33_ASAP7_75t_R g6590 ( 
.A(n_702),
.Y(n_6590)
);

CKINVDCx5p33_ASAP7_75t_R g6591 ( 
.A(n_4445),
.Y(n_6591)
);

CKINVDCx5p33_ASAP7_75t_R g6592 ( 
.A(n_1189),
.Y(n_6592)
);

CKINVDCx5p33_ASAP7_75t_R g6593 ( 
.A(n_4673),
.Y(n_6593)
);

BUFx6f_ASAP7_75t_L g6594 ( 
.A(n_1590),
.Y(n_6594)
);

BUFx10_ASAP7_75t_L g6595 ( 
.A(n_4493),
.Y(n_6595)
);

BUFx3_ASAP7_75t_L g6596 ( 
.A(n_206),
.Y(n_6596)
);

CKINVDCx5p33_ASAP7_75t_R g6597 ( 
.A(n_5310),
.Y(n_6597)
);

INVx1_ASAP7_75t_SL g6598 ( 
.A(n_1109),
.Y(n_6598)
);

CKINVDCx20_ASAP7_75t_R g6599 ( 
.A(n_4531),
.Y(n_6599)
);

CKINVDCx5p33_ASAP7_75t_R g6600 ( 
.A(n_787),
.Y(n_6600)
);

CKINVDCx5p33_ASAP7_75t_R g6601 ( 
.A(n_236),
.Y(n_6601)
);

CKINVDCx5p33_ASAP7_75t_R g6602 ( 
.A(n_225),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_847),
.Y(n_6603)
);

INVx2_ASAP7_75t_L g6604 ( 
.A(n_4488),
.Y(n_6604)
);

CKINVDCx5p33_ASAP7_75t_R g6605 ( 
.A(n_5575),
.Y(n_6605)
);

CKINVDCx5p33_ASAP7_75t_R g6606 ( 
.A(n_3641),
.Y(n_6606)
);

CKINVDCx5p33_ASAP7_75t_R g6607 ( 
.A(n_1455),
.Y(n_6607)
);

INVx2_ASAP7_75t_L g6608 ( 
.A(n_3522),
.Y(n_6608)
);

CKINVDCx5p33_ASAP7_75t_R g6609 ( 
.A(n_5365),
.Y(n_6609)
);

CKINVDCx5p33_ASAP7_75t_R g6610 ( 
.A(n_1188),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_4380),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_870),
.Y(n_6612)
);

CKINVDCx5p33_ASAP7_75t_R g6613 ( 
.A(n_4626),
.Y(n_6613)
);

CKINVDCx5p33_ASAP7_75t_R g6614 ( 
.A(n_5215),
.Y(n_6614)
);

INVx2_ASAP7_75t_L g6615 ( 
.A(n_5514),
.Y(n_6615)
);

CKINVDCx5p33_ASAP7_75t_R g6616 ( 
.A(n_3431),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_474),
.Y(n_6617)
);

CKINVDCx5p33_ASAP7_75t_R g6618 ( 
.A(n_2296),
.Y(n_6618)
);

CKINVDCx5p33_ASAP7_75t_R g6619 ( 
.A(n_2752),
.Y(n_6619)
);

BUFx10_ASAP7_75t_L g6620 ( 
.A(n_3597),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_2957),
.Y(n_6621)
);

CKINVDCx5p33_ASAP7_75t_R g6622 ( 
.A(n_5043),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_4414),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_4460),
.Y(n_6624)
);

CKINVDCx5p33_ASAP7_75t_R g6625 ( 
.A(n_1707),
.Y(n_6625)
);

CKINVDCx5p33_ASAP7_75t_R g6626 ( 
.A(n_1353),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6064),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_2160),
.Y(n_6628)
);

BUFx10_ASAP7_75t_L g6629 ( 
.A(n_2108),
.Y(n_6629)
);

CKINVDCx5p33_ASAP7_75t_R g6630 ( 
.A(n_2252),
.Y(n_6630)
);

CKINVDCx5p33_ASAP7_75t_R g6631 ( 
.A(n_4680),
.Y(n_6631)
);

CKINVDCx20_ASAP7_75t_R g6632 ( 
.A(n_6009),
.Y(n_6632)
);

CKINVDCx5p33_ASAP7_75t_R g6633 ( 
.A(n_4879),
.Y(n_6633)
);

CKINVDCx16_ASAP7_75t_R g6634 ( 
.A(n_4540),
.Y(n_6634)
);

CKINVDCx5p33_ASAP7_75t_R g6635 ( 
.A(n_4471),
.Y(n_6635)
);

CKINVDCx5p33_ASAP7_75t_R g6636 ( 
.A(n_991),
.Y(n_6636)
);

CKINVDCx5p33_ASAP7_75t_R g6637 ( 
.A(n_6050),
.Y(n_6637)
);

BUFx6f_ASAP7_75t_L g6638 ( 
.A(n_2183),
.Y(n_6638)
);

INVx2_ASAP7_75t_SL g6639 ( 
.A(n_1203),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_922),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_4672),
.Y(n_6641)
);

INVx2_ASAP7_75t_SL g6642 ( 
.A(n_4533),
.Y(n_6642)
);

CKINVDCx5p33_ASAP7_75t_R g6643 ( 
.A(n_5324),
.Y(n_6643)
);

CKINVDCx5p33_ASAP7_75t_R g6644 ( 
.A(n_3083),
.Y(n_6644)
);

INVx1_ASAP7_75t_SL g6645 ( 
.A(n_5034),
.Y(n_6645)
);

CKINVDCx5p33_ASAP7_75t_R g6646 ( 
.A(n_31),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_595),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_5624),
.Y(n_6648)
);

CKINVDCx11_ASAP7_75t_R g6649 ( 
.A(n_5531),
.Y(n_6649)
);

CKINVDCx5p33_ASAP7_75t_R g6650 ( 
.A(n_1727),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_2887),
.Y(n_6651)
);

CKINVDCx5p33_ASAP7_75t_R g6652 ( 
.A(n_6065),
.Y(n_6652)
);

CKINVDCx20_ASAP7_75t_R g6653 ( 
.A(n_2486),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_3771),
.Y(n_6654)
);

BUFx6f_ASAP7_75t_L g6655 ( 
.A(n_4547),
.Y(n_6655)
);

CKINVDCx20_ASAP7_75t_R g6656 ( 
.A(n_3418),
.Y(n_6656)
);

INVx1_ASAP7_75t_L g6657 ( 
.A(n_2840),
.Y(n_6657)
);

CKINVDCx5p33_ASAP7_75t_R g6658 ( 
.A(n_4398),
.Y(n_6658)
);

CKINVDCx20_ASAP7_75t_R g6659 ( 
.A(n_4284),
.Y(n_6659)
);

CKINVDCx5p33_ASAP7_75t_R g6660 ( 
.A(n_2508),
.Y(n_6660)
);

CKINVDCx5p33_ASAP7_75t_R g6661 ( 
.A(n_4939),
.Y(n_6661)
);

CKINVDCx5p33_ASAP7_75t_R g6662 ( 
.A(n_5746),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_916),
.Y(n_6663)
);

CKINVDCx5p33_ASAP7_75t_R g6664 ( 
.A(n_4373),
.Y(n_6664)
);

INVx1_ASAP7_75t_SL g6665 ( 
.A(n_1260),
.Y(n_6665)
);

INVxp67_ASAP7_75t_L g6666 ( 
.A(n_2450),
.Y(n_6666)
);

BUFx2_ASAP7_75t_L g6667 ( 
.A(n_1285),
.Y(n_6667)
);

CKINVDCx5p33_ASAP7_75t_R g6668 ( 
.A(n_2287),
.Y(n_6668)
);

CKINVDCx5p33_ASAP7_75t_R g6669 ( 
.A(n_2062),
.Y(n_6669)
);

CKINVDCx5p33_ASAP7_75t_R g6670 ( 
.A(n_5779),
.Y(n_6670)
);

CKINVDCx5p33_ASAP7_75t_R g6671 ( 
.A(n_658),
.Y(n_6671)
);

CKINVDCx5p33_ASAP7_75t_R g6672 ( 
.A(n_1136),
.Y(n_6672)
);

CKINVDCx5p33_ASAP7_75t_R g6673 ( 
.A(n_3612),
.Y(n_6673)
);

CKINVDCx5p33_ASAP7_75t_R g6674 ( 
.A(n_2235),
.Y(n_6674)
);

INVx2_ASAP7_75t_L g6675 ( 
.A(n_3925),
.Y(n_6675)
);

HB1xp67_ASAP7_75t_L g6676 ( 
.A(n_5441),
.Y(n_6676)
);

CKINVDCx5p33_ASAP7_75t_R g6677 ( 
.A(n_5364),
.Y(n_6677)
);

INVx2_ASAP7_75t_L g6678 ( 
.A(n_1979),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_1095),
.Y(n_6679)
);

INVx2_ASAP7_75t_L g6680 ( 
.A(n_2724),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_1178),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_1370),
.Y(n_6682)
);

CKINVDCx5p33_ASAP7_75t_R g6683 ( 
.A(n_5121),
.Y(n_6683)
);

CKINVDCx5p33_ASAP7_75t_R g6684 ( 
.A(n_632),
.Y(n_6684)
);

CKINVDCx5p33_ASAP7_75t_R g6685 ( 
.A(n_3731),
.Y(n_6685)
);

CKINVDCx5p33_ASAP7_75t_R g6686 ( 
.A(n_4208),
.Y(n_6686)
);

CKINVDCx5p33_ASAP7_75t_R g6687 ( 
.A(n_3746),
.Y(n_6687)
);

BUFx6f_ASAP7_75t_L g6688 ( 
.A(n_4598),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_1422),
.Y(n_6689)
);

CKINVDCx5p33_ASAP7_75t_R g6690 ( 
.A(n_4286),
.Y(n_6690)
);

CKINVDCx5p33_ASAP7_75t_R g6691 ( 
.A(n_3984),
.Y(n_6691)
);

BUFx6f_ASAP7_75t_L g6692 ( 
.A(n_641),
.Y(n_6692)
);

CKINVDCx5p33_ASAP7_75t_R g6693 ( 
.A(n_5495),
.Y(n_6693)
);

CKINVDCx20_ASAP7_75t_R g6694 ( 
.A(n_6046),
.Y(n_6694)
);

CKINVDCx5p33_ASAP7_75t_R g6695 ( 
.A(n_4489),
.Y(n_6695)
);

BUFx10_ASAP7_75t_L g6696 ( 
.A(n_4518),
.Y(n_6696)
);

INVx1_ASAP7_75t_L g6697 ( 
.A(n_5613),
.Y(n_6697)
);

CKINVDCx5p33_ASAP7_75t_R g6698 ( 
.A(n_5904),
.Y(n_6698)
);

BUFx5_ASAP7_75t_L g6699 ( 
.A(n_1613),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_4499),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_4473),
.Y(n_6701)
);

CKINVDCx20_ASAP7_75t_R g6702 ( 
.A(n_3530),
.Y(n_6702)
);

CKINVDCx5p33_ASAP7_75t_R g6703 ( 
.A(n_4470),
.Y(n_6703)
);

CKINVDCx5p33_ASAP7_75t_R g6704 ( 
.A(n_265),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_2376),
.Y(n_6705)
);

CKINVDCx5p33_ASAP7_75t_R g6706 ( 
.A(n_3508),
.Y(n_6706)
);

HB1xp67_ASAP7_75t_L g6707 ( 
.A(n_2977),
.Y(n_6707)
);

CKINVDCx5p33_ASAP7_75t_R g6708 ( 
.A(n_3275),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_695),
.Y(n_6709)
);

CKINVDCx5p33_ASAP7_75t_R g6710 ( 
.A(n_734),
.Y(n_6710)
);

CKINVDCx5p33_ASAP7_75t_R g6711 ( 
.A(n_4031),
.Y(n_6711)
);

CKINVDCx5p33_ASAP7_75t_R g6712 ( 
.A(n_6029),
.Y(n_6712)
);

CKINVDCx5p33_ASAP7_75t_R g6713 ( 
.A(n_3724),
.Y(n_6713)
);

CKINVDCx5p33_ASAP7_75t_R g6714 ( 
.A(n_3766),
.Y(n_6714)
);

CKINVDCx5p33_ASAP7_75t_R g6715 ( 
.A(n_2697),
.Y(n_6715)
);

INVx2_ASAP7_75t_L g6716 ( 
.A(n_4463),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_3475),
.Y(n_6717)
);

CKINVDCx5p33_ASAP7_75t_R g6718 ( 
.A(n_5670),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_4424),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_2931),
.Y(n_6720)
);

CKINVDCx5p33_ASAP7_75t_R g6721 ( 
.A(n_3565),
.Y(n_6721)
);

CKINVDCx5p33_ASAP7_75t_R g6722 ( 
.A(n_667),
.Y(n_6722)
);

CKINVDCx5p33_ASAP7_75t_R g6723 ( 
.A(n_393),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_3794),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_4422),
.Y(n_6725)
);

CKINVDCx5p33_ASAP7_75t_R g6726 ( 
.A(n_3855),
.Y(n_6726)
);

CKINVDCx5p33_ASAP7_75t_R g6727 ( 
.A(n_2854),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_3045),
.Y(n_6728)
);

CKINVDCx5p33_ASAP7_75t_R g6729 ( 
.A(n_1106),
.Y(n_6729)
);

CKINVDCx5p33_ASAP7_75t_R g6730 ( 
.A(n_4391),
.Y(n_6730)
);

BUFx2_ASAP7_75t_L g6731 ( 
.A(n_2590),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_777),
.Y(n_6732)
);

CKINVDCx5p33_ASAP7_75t_R g6733 ( 
.A(n_2654),
.Y(n_6733)
);

CKINVDCx20_ASAP7_75t_R g6734 ( 
.A(n_2557),
.Y(n_6734)
);

INVxp67_ASAP7_75t_L g6735 ( 
.A(n_2952),
.Y(n_6735)
);

INVx1_ASAP7_75t_L g6736 ( 
.A(n_2844),
.Y(n_6736)
);

BUFx10_ASAP7_75t_L g6737 ( 
.A(n_877),
.Y(n_6737)
);

CKINVDCx5p33_ASAP7_75t_R g6738 ( 
.A(n_3723),
.Y(n_6738)
);

CKINVDCx5p33_ASAP7_75t_R g6739 ( 
.A(n_3869),
.Y(n_6739)
);

CKINVDCx5p33_ASAP7_75t_R g6740 ( 
.A(n_2848),
.Y(n_6740)
);

CKINVDCx5p33_ASAP7_75t_R g6741 ( 
.A(n_3070),
.Y(n_6741)
);

CKINVDCx5p33_ASAP7_75t_R g6742 ( 
.A(n_3086),
.Y(n_6742)
);

CKINVDCx5p33_ASAP7_75t_R g6743 ( 
.A(n_5630),
.Y(n_6743)
);

INVx1_ASAP7_75t_L g6744 ( 
.A(n_4182),
.Y(n_6744)
);

CKINVDCx5p33_ASAP7_75t_R g6745 ( 
.A(n_6049),
.Y(n_6745)
);

CKINVDCx14_ASAP7_75t_R g6746 ( 
.A(n_5289),
.Y(n_6746)
);

CKINVDCx5p33_ASAP7_75t_R g6747 ( 
.A(n_3984),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_3113),
.Y(n_6748)
);

INVx2_ASAP7_75t_L g6749 ( 
.A(n_1052),
.Y(n_6749)
);

CKINVDCx20_ASAP7_75t_R g6750 ( 
.A(n_288),
.Y(n_6750)
);

CKINVDCx5p33_ASAP7_75t_R g6751 ( 
.A(n_1404),
.Y(n_6751)
);

CKINVDCx5p33_ASAP7_75t_R g6752 ( 
.A(n_5679),
.Y(n_6752)
);

CKINVDCx5p33_ASAP7_75t_R g6753 ( 
.A(n_345),
.Y(n_6753)
);

CKINVDCx5p33_ASAP7_75t_R g6754 ( 
.A(n_5775),
.Y(n_6754)
);

INVx1_ASAP7_75t_L g6755 ( 
.A(n_914),
.Y(n_6755)
);

CKINVDCx5p33_ASAP7_75t_R g6756 ( 
.A(n_3339),
.Y(n_6756)
);

CKINVDCx5p33_ASAP7_75t_R g6757 ( 
.A(n_5484),
.Y(n_6757)
);

CKINVDCx16_ASAP7_75t_R g6758 ( 
.A(n_1811),
.Y(n_6758)
);

INVx2_ASAP7_75t_L g6759 ( 
.A(n_901),
.Y(n_6759)
);

CKINVDCx5p33_ASAP7_75t_R g6760 ( 
.A(n_3163),
.Y(n_6760)
);

CKINVDCx5p33_ASAP7_75t_R g6761 ( 
.A(n_4416),
.Y(n_6761)
);

CKINVDCx5p33_ASAP7_75t_R g6762 ( 
.A(n_3061),
.Y(n_6762)
);

CKINVDCx5p33_ASAP7_75t_R g6763 ( 
.A(n_3040),
.Y(n_6763)
);

CKINVDCx5p33_ASAP7_75t_R g6764 ( 
.A(n_5848),
.Y(n_6764)
);

INVx1_ASAP7_75t_SL g6765 ( 
.A(n_6025),
.Y(n_6765)
);

CKINVDCx5p33_ASAP7_75t_R g6766 ( 
.A(n_3675),
.Y(n_6766)
);

CKINVDCx5p33_ASAP7_75t_R g6767 ( 
.A(n_2590),
.Y(n_6767)
);

CKINVDCx5p33_ASAP7_75t_R g6768 ( 
.A(n_4496),
.Y(n_6768)
);

CKINVDCx20_ASAP7_75t_R g6769 ( 
.A(n_3018),
.Y(n_6769)
);

CKINVDCx5p33_ASAP7_75t_R g6770 ( 
.A(n_5293),
.Y(n_6770)
);

BUFx10_ASAP7_75t_L g6771 ( 
.A(n_4530),
.Y(n_6771)
);

CKINVDCx5p33_ASAP7_75t_R g6772 ( 
.A(n_4492),
.Y(n_6772)
);

CKINVDCx5p33_ASAP7_75t_R g6773 ( 
.A(n_2217),
.Y(n_6773)
);

CKINVDCx5p33_ASAP7_75t_R g6774 ( 
.A(n_3602),
.Y(n_6774)
);

CKINVDCx5p33_ASAP7_75t_R g6775 ( 
.A(n_2066),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_4456),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_4307),
.Y(n_6777)
);

CKINVDCx20_ASAP7_75t_R g6778 ( 
.A(n_3911),
.Y(n_6778)
);

CKINVDCx5p33_ASAP7_75t_R g6779 ( 
.A(n_4426),
.Y(n_6779)
);

CKINVDCx5p33_ASAP7_75t_R g6780 ( 
.A(n_5017),
.Y(n_6780)
);

INVxp67_ASAP7_75t_L g6781 ( 
.A(n_2319),
.Y(n_6781)
);

CKINVDCx5p33_ASAP7_75t_R g6782 ( 
.A(n_4440),
.Y(n_6782)
);

CKINVDCx5p33_ASAP7_75t_R g6783 ( 
.A(n_482),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_3226),
.Y(n_6784)
);

CKINVDCx5p33_ASAP7_75t_R g6785 ( 
.A(n_437),
.Y(n_6785)
);

INVx1_ASAP7_75t_SL g6786 ( 
.A(n_5486),
.Y(n_6786)
);

CKINVDCx20_ASAP7_75t_R g6787 ( 
.A(n_4057),
.Y(n_6787)
);

CKINVDCx16_ASAP7_75t_R g6788 ( 
.A(n_4481),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_4468),
.Y(n_6789)
);

CKINVDCx5p33_ASAP7_75t_R g6790 ( 
.A(n_3637),
.Y(n_6790)
);

BUFx3_ASAP7_75t_L g6791 ( 
.A(n_2067),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_4518),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_3585),
.Y(n_6793)
);

INVx1_ASAP7_75t_SL g6794 ( 
.A(n_4149),
.Y(n_6794)
);

CKINVDCx16_ASAP7_75t_R g6795 ( 
.A(n_4223),
.Y(n_6795)
);

CKINVDCx5p33_ASAP7_75t_R g6796 ( 
.A(n_5468),
.Y(n_6796)
);

INVx1_ASAP7_75t_L g6797 ( 
.A(n_2029),
.Y(n_6797)
);

CKINVDCx5p33_ASAP7_75t_R g6798 ( 
.A(n_529),
.Y(n_6798)
);

CKINVDCx5p33_ASAP7_75t_R g6799 ( 
.A(n_1595),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_5717),
.Y(n_6800)
);

CKINVDCx20_ASAP7_75t_R g6801 ( 
.A(n_307),
.Y(n_6801)
);

CKINVDCx5p33_ASAP7_75t_R g6802 ( 
.A(n_4720),
.Y(n_6802)
);

INVx2_ASAP7_75t_SL g6803 ( 
.A(n_6074),
.Y(n_6803)
);

CKINVDCx5p33_ASAP7_75t_R g6804 ( 
.A(n_1236),
.Y(n_6804)
);

CKINVDCx5p33_ASAP7_75t_R g6805 ( 
.A(n_5998),
.Y(n_6805)
);

CKINVDCx5p33_ASAP7_75t_R g6806 ( 
.A(n_3661),
.Y(n_6806)
);

BUFx6f_ASAP7_75t_L g6807 ( 
.A(n_3662),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_5933),
.Y(n_6808)
);

CKINVDCx16_ASAP7_75t_R g6809 ( 
.A(n_3734),
.Y(n_6809)
);

CKINVDCx5p33_ASAP7_75t_R g6810 ( 
.A(n_1277),
.Y(n_6810)
);

CKINVDCx5p33_ASAP7_75t_R g6811 ( 
.A(n_1865),
.Y(n_6811)
);

CKINVDCx5p33_ASAP7_75t_R g6812 ( 
.A(n_6068),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_4270),
.Y(n_6813)
);

CKINVDCx5p33_ASAP7_75t_R g6814 ( 
.A(n_1467),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_3942),
.Y(n_6815)
);

CKINVDCx5p33_ASAP7_75t_R g6816 ( 
.A(n_4525),
.Y(n_6816)
);

CKINVDCx20_ASAP7_75t_R g6817 ( 
.A(n_1314),
.Y(n_6817)
);

CKINVDCx20_ASAP7_75t_R g6818 ( 
.A(n_3904),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_2230),
.Y(n_6819)
);

CKINVDCx5p33_ASAP7_75t_R g6820 ( 
.A(n_1391),
.Y(n_6820)
);

CKINVDCx16_ASAP7_75t_R g6821 ( 
.A(n_534),
.Y(n_6821)
);

CKINVDCx5p33_ASAP7_75t_R g6822 ( 
.A(n_4450),
.Y(n_6822)
);

CKINVDCx5p33_ASAP7_75t_R g6823 ( 
.A(n_3519),
.Y(n_6823)
);

INVxp67_ASAP7_75t_L g6824 ( 
.A(n_5611),
.Y(n_6824)
);

INVx1_ASAP7_75t_L g6825 ( 
.A(n_5246),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_3050),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_919),
.Y(n_6827)
);

CKINVDCx5p33_ASAP7_75t_R g6828 ( 
.A(n_4320),
.Y(n_6828)
);

CKINVDCx5p33_ASAP7_75t_R g6829 ( 
.A(n_3427),
.Y(n_6829)
);

INVx1_ASAP7_75t_L g6830 ( 
.A(n_1442),
.Y(n_6830)
);

CKINVDCx5p33_ASAP7_75t_R g6831 ( 
.A(n_1731),
.Y(n_6831)
);

CKINVDCx5p33_ASAP7_75t_R g6832 ( 
.A(n_4437),
.Y(n_6832)
);

CKINVDCx5p33_ASAP7_75t_R g6833 ( 
.A(n_5499),
.Y(n_6833)
);

INVx1_ASAP7_75t_L g6834 ( 
.A(n_307),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_4461),
.Y(n_6835)
);

CKINVDCx5p33_ASAP7_75t_R g6836 ( 
.A(n_4956),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_368),
.Y(n_6837)
);

BUFx3_ASAP7_75t_L g6838 ( 
.A(n_102),
.Y(n_6838)
);

BUFx10_ASAP7_75t_L g6839 ( 
.A(n_1767),
.Y(n_6839)
);

CKINVDCx5p33_ASAP7_75t_R g6840 ( 
.A(n_2062),
.Y(n_6840)
);

CKINVDCx5p33_ASAP7_75t_R g6841 ( 
.A(n_711),
.Y(n_6841)
);

INVx2_ASAP7_75t_L g6842 ( 
.A(n_3114),
.Y(n_6842)
);

CKINVDCx5p33_ASAP7_75t_R g6843 ( 
.A(n_3983),
.Y(n_6843)
);

CKINVDCx5p33_ASAP7_75t_R g6844 ( 
.A(n_3007),
.Y(n_6844)
);

CKINVDCx5p33_ASAP7_75t_R g6845 ( 
.A(n_3778),
.Y(n_6845)
);

CKINVDCx5p33_ASAP7_75t_R g6846 ( 
.A(n_1884),
.Y(n_6846)
);

INVx2_ASAP7_75t_L g6847 ( 
.A(n_5571),
.Y(n_6847)
);

CKINVDCx5p33_ASAP7_75t_R g6848 ( 
.A(n_2381),
.Y(n_6848)
);

CKINVDCx5p33_ASAP7_75t_R g6849 ( 
.A(n_3581),
.Y(n_6849)
);

INVx1_ASAP7_75t_L g6850 ( 
.A(n_3),
.Y(n_6850)
);

CKINVDCx5p33_ASAP7_75t_R g6851 ( 
.A(n_319),
.Y(n_6851)
);

CKINVDCx5p33_ASAP7_75t_R g6852 ( 
.A(n_5232),
.Y(n_6852)
);

CKINVDCx16_ASAP7_75t_R g6853 ( 
.A(n_2554),
.Y(n_6853)
);

CKINVDCx5p33_ASAP7_75t_R g6854 ( 
.A(n_1417),
.Y(n_6854)
);

CKINVDCx5p33_ASAP7_75t_R g6855 ( 
.A(n_4410),
.Y(n_6855)
);

INVx1_ASAP7_75t_SL g6856 ( 
.A(n_1596),
.Y(n_6856)
);

INVx2_ASAP7_75t_L g6857 ( 
.A(n_5593),
.Y(n_6857)
);

CKINVDCx5p33_ASAP7_75t_R g6858 ( 
.A(n_5133),
.Y(n_6858)
);

INVx1_ASAP7_75t_SL g6859 ( 
.A(n_5868),
.Y(n_6859)
);

CKINVDCx5p33_ASAP7_75t_R g6860 ( 
.A(n_5965),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_4967),
.Y(n_6861)
);

CKINVDCx20_ASAP7_75t_R g6862 ( 
.A(n_4876),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_1343),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6048),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_4360),
.Y(n_6865)
);

CKINVDCx5p33_ASAP7_75t_R g6866 ( 
.A(n_341),
.Y(n_6866)
);

CKINVDCx5p33_ASAP7_75t_R g6867 ( 
.A(n_4415),
.Y(n_6867)
);

INVx2_ASAP7_75t_L g6868 ( 
.A(n_4594),
.Y(n_6868)
);

CKINVDCx5p33_ASAP7_75t_R g6869 ( 
.A(n_2708),
.Y(n_6869)
);

BUFx6f_ASAP7_75t_L g6870 ( 
.A(n_5124),
.Y(n_6870)
);

BUFx2_ASAP7_75t_SL g6871 ( 
.A(n_3236),
.Y(n_6871)
);

CKINVDCx5p33_ASAP7_75t_R g6872 ( 
.A(n_1926),
.Y(n_6872)
);

CKINVDCx5p33_ASAP7_75t_R g6873 ( 
.A(n_749),
.Y(n_6873)
);

BUFx3_ASAP7_75t_L g6874 ( 
.A(n_1395),
.Y(n_6874)
);

CKINVDCx5p33_ASAP7_75t_R g6875 ( 
.A(n_1492),
.Y(n_6875)
);

CKINVDCx5p33_ASAP7_75t_R g6876 ( 
.A(n_596),
.Y(n_6876)
);

CKINVDCx5p33_ASAP7_75t_R g6877 ( 
.A(n_4702),
.Y(n_6877)
);

CKINVDCx5p33_ASAP7_75t_R g6878 ( 
.A(n_2515),
.Y(n_6878)
);

INVx2_ASAP7_75t_L g6879 ( 
.A(n_586),
.Y(n_6879)
);

CKINVDCx5p33_ASAP7_75t_R g6880 ( 
.A(n_5905),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_3672),
.Y(n_6881)
);

CKINVDCx5p33_ASAP7_75t_R g6882 ( 
.A(n_850),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_3934),
.Y(n_6883)
);

CKINVDCx5p33_ASAP7_75t_R g6884 ( 
.A(n_3113),
.Y(n_6884)
);

CKINVDCx5p33_ASAP7_75t_R g6885 ( 
.A(n_998),
.Y(n_6885)
);

CKINVDCx5p33_ASAP7_75t_R g6886 ( 
.A(n_1445),
.Y(n_6886)
);

CKINVDCx20_ASAP7_75t_R g6887 ( 
.A(n_1913),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_593),
.Y(n_6888)
);

INVx1_ASAP7_75t_L g6889 ( 
.A(n_909),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_529),
.Y(n_6890)
);

INVxp67_ASAP7_75t_SL g6891 ( 
.A(n_1346),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_2939),
.Y(n_6892)
);

CKINVDCx5p33_ASAP7_75t_R g6893 ( 
.A(n_5218),
.Y(n_6893)
);

CKINVDCx5p33_ASAP7_75t_R g6894 ( 
.A(n_1638),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_3611),
.Y(n_6895)
);

CKINVDCx5p33_ASAP7_75t_R g6896 ( 
.A(n_3409),
.Y(n_6896)
);

CKINVDCx5p33_ASAP7_75t_R g6897 ( 
.A(n_5572),
.Y(n_6897)
);

CKINVDCx5p33_ASAP7_75t_R g6898 ( 
.A(n_2107),
.Y(n_6898)
);

INVx1_ASAP7_75t_SL g6899 ( 
.A(n_4138),
.Y(n_6899)
);

CKINVDCx5p33_ASAP7_75t_R g6900 ( 
.A(n_5564),
.Y(n_6900)
);

INVx1_ASAP7_75t_L g6901 ( 
.A(n_4385),
.Y(n_6901)
);

INVx2_ASAP7_75t_SL g6902 ( 
.A(n_5949),
.Y(n_6902)
);

CKINVDCx5p33_ASAP7_75t_R g6903 ( 
.A(n_2906),
.Y(n_6903)
);

CKINVDCx5p33_ASAP7_75t_R g6904 ( 
.A(n_2900),
.Y(n_6904)
);

CKINVDCx5p33_ASAP7_75t_R g6905 ( 
.A(n_1303),
.Y(n_6905)
);

CKINVDCx5p33_ASAP7_75t_R g6906 ( 
.A(n_4142),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_2772),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_3487),
.Y(n_6908)
);

CKINVDCx5p33_ASAP7_75t_R g6909 ( 
.A(n_3324),
.Y(n_6909)
);

CKINVDCx5p33_ASAP7_75t_R g6910 ( 
.A(n_158),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_1490),
.Y(n_6911)
);

BUFx6f_ASAP7_75t_L g6912 ( 
.A(n_1190),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_644),
.Y(n_6913)
);

CKINVDCx5p33_ASAP7_75t_R g6914 ( 
.A(n_3553),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_4985),
.Y(n_6915)
);

CKINVDCx5p33_ASAP7_75t_R g6916 ( 
.A(n_2408),
.Y(n_6916)
);

CKINVDCx5p33_ASAP7_75t_R g6917 ( 
.A(n_4014),
.Y(n_6917)
);

CKINVDCx5p33_ASAP7_75t_R g6918 ( 
.A(n_2435),
.Y(n_6918)
);

CKINVDCx5p33_ASAP7_75t_R g6919 ( 
.A(n_3030),
.Y(n_6919)
);

CKINVDCx5p33_ASAP7_75t_R g6920 ( 
.A(n_6071),
.Y(n_6920)
);

CKINVDCx5p33_ASAP7_75t_R g6921 ( 
.A(n_4715),
.Y(n_6921)
);

CKINVDCx5p33_ASAP7_75t_R g6922 ( 
.A(n_2404),
.Y(n_6922)
);

CKINVDCx5p33_ASAP7_75t_R g6923 ( 
.A(n_5357),
.Y(n_6923)
);

CKINVDCx20_ASAP7_75t_R g6924 ( 
.A(n_1881),
.Y(n_6924)
);

CKINVDCx5p33_ASAP7_75t_R g6925 ( 
.A(n_5929),
.Y(n_6925)
);

CKINVDCx20_ASAP7_75t_R g6926 ( 
.A(n_2365),
.Y(n_6926)
);

CKINVDCx5p33_ASAP7_75t_R g6927 ( 
.A(n_3785),
.Y(n_6927)
);

INVx2_ASAP7_75t_SL g6928 ( 
.A(n_1386),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_3465),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_1835),
.Y(n_6930)
);

CKINVDCx5p33_ASAP7_75t_R g6931 ( 
.A(n_5307),
.Y(n_6931)
);

CKINVDCx5p33_ASAP7_75t_R g6932 ( 
.A(n_2006),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_3202),
.Y(n_6933)
);

CKINVDCx5p33_ASAP7_75t_R g6934 ( 
.A(n_3234),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_4511),
.Y(n_6935)
);

CKINVDCx20_ASAP7_75t_R g6936 ( 
.A(n_2276),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_4883),
.Y(n_6937)
);

CKINVDCx5p33_ASAP7_75t_R g6938 ( 
.A(n_501),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_11),
.Y(n_6939)
);

CKINVDCx20_ASAP7_75t_R g6940 ( 
.A(n_3052),
.Y(n_6940)
);

CKINVDCx5p33_ASAP7_75t_R g6941 ( 
.A(n_4685),
.Y(n_6941)
);

CKINVDCx5p33_ASAP7_75t_R g6942 ( 
.A(n_2725),
.Y(n_6942)
);

CKINVDCx5p33_ASAP7_75t_R g6943 ( 
.A(n_6066),
.Y(n_6943)
);

CKINVDCx5p33_ASAP7_75t_R g6944 ( 
.A(n_1353),
.Y(n_6944)
);

BUFx2_ASAP7_75t_L g6945 ( 
.A(n_1053),
.Y(n_6945)
);

CKINVDCx20_ASAP7_75t_R g6946 ( 
.A(n_1812),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_4509),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_2247),
.Y(n_6948)
);

BUFx3_ASAP7_75t_L g6949 ( 
.A(n_2319),
.Y(n_6949)
);

CKINVDCx5p33_ASAP7_75t_R g6950 ( 
.A(n_5968),
.Y(n_6950)
);

CKINVDCx5p33_ASAP7_75t_R g6951 ( 
.A(n_1084),
.Y(n_6951)
);

INVx1_ASAP7_75t_SL g6952 ( 
.A(n_5972),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_5266),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_243),
.Y(n_6954)
);

CKINVDCx5p33_ASAP7_75t_R g6955 ( 
.A(n_2578),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_4671),
.Y(n_6956)
);

CKINVDCx16_ASAP7_75t_R g6957 ( 
.A(n_4538),
.Y(n_6957)
);

CKINVDCx5p33_ASAP7_75t_R g6958 ( 
.A(n_3730),
.Y(n_6958)
);

BUFx3_ASAP7_75t_L g6959 ( 
.A(n_793),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_3919),
.Y(n_6960)
);

CKINVDCx5p33_ASAP7_75t_R g6961 ( 
.A(n_3432),
.Y(n_6961)
);

CKINVDCx5p33_ASAP7_75t_R g6962 ( 
.A(n_4527),
.Y(n_6962)
);

BUFx10_ASAP7_75t_L g6963 ( 
.A(n_4851),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_1364),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_5749),
.Y(n_6965)
);

CKINVDCx5p33_ASAP7_75t_R g6966 ( 
.A(n_5917),
.Y(n_6966)
);

CKINVDCx5p33_ASAP7_75t_R g6967 ( 
.A(n_947),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_1446),
.Y(n_6968)
);

CKINVDCx5p33_ASAP7_75t_R g6969 ( 
.A(n_4369),
.Y(n_6969)
);

CKINVDCx5p33_ASAP7_75t_R g6970 ( 
.A(n_3491),
.Y(n_6970)
);

CKINVDCx20_ASAP7_75t_R g6971 ( 
.A(n_1185),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_4420),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_4480),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_2540),
.Y(n_6974)
);

BUFx3_ASAP7_75t_L g6975 ( 
.A(n_4399),
.Y(n_6975)
);

INVx1_ASAP7_75t_L g6976 ( 
.A(n_93),
.Y(n_6976)
);

BUFx3_ASAP7_75t_L g6977 ( 
.A(n_5511),
.Y(n_6977)
);

CKINVDCx5p33_ASAP7_75t_R g6978 ( 
.A(n_1114),
.Y(n_6978)
);

CKINVDCx5p33_ASAP7_75t_R g6979 ( 
.A(n_4794),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_2342),
.Y(n_6980)
);

CKINVDCx5p33_ASAP7_75t_R g6981 ( 
.A(n_107),
.Y(n_6981)
);

CKINVDCx5p33_ASAP7_75t_R g6982 ( 
.A(n_271),
.Y(n_6982)
);

CKINVDCx5p33_ASAP7_75t_R g6983 ( 
.A(n_4095),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_4017),
.Y(n_6984)
);

CKINVDCx20_ASAP7_75t_R g6985 ( 
.A(n_4431),
.Y(n_6985)
);

CKINVDCx5p33_ASAP7_75t_R g6986 ( 
.A(n_4428),
.Y(n_6986)
);

CKINVDCx5p33_ASAP7_75t_R g6987 ( 
.A(n_156),
.Y(n_6987)
);

CKINVDCx5p33_ASAP7_75t_R g6988 ( 
.A(n_3863),
.Y(n_6988)
);

CKINVDCx5p33_ASAP7_75t_R g6989 ( 
.A(n_4508),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_5057),
.Y(n_6990)
);

CKINVDCx5p33_ASAP7_75t_R g6991 ( 
.A(n_2798),
.Y(n_6991)
);

CKINVDCx5p33_ASAP7_75t_R g6992 ( 
.A(n_896),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_4378),
.Y(n_6993)
);

CKINVDCx5p33_ASAP7_75t_R g6994 ( 
.A(n_516),
.Y(n_6994)
);

CKINVDCx5p33_ASAP7_75t_R g6995 ( 
.A(n_5543),
.Y(n_6995)
);

CKINVDCx5p33_ASAP7_75t_R g6996 ( 
.A(n_3365),
.Y(n_6996)
);

CKINVDCx5p33_ASAP7_75t_R g6997 ( 
.A(n_2096),
.Y(n_6997)
);

CKINVDCx5p33_ASAP7_75t_R g6998 ( 
.A(n_5383),
.Y(n_6998)
);

CKINVDCx20_ASAP7_75t_R g6999 ( 
.A(n_5751),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_1194),
.Y(n_7000)
);

BUFx3_ASAP7_75t_L g7001 ( 
.A(n_5222),
.Y(n_7001)
);

CKINVDCx5p33_ASAP7_75t_R g7002 ( 
.A(n_2215),
.Y(n_7002)
);

CKINVDCx5p33_ASAP7_75t_R g7003 ( 
.A(n_4411),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6062),
.Y(n_7004)
);

CKINVDCx5p33_ASAP7_75t_R g7005 ( 
.A(n_627),
.Y(n_7005)
);

CKINVDCx5p33_ASAP7_75t_R g7006 ( 
.A(n_4361),
.Y(n_7006)
);

INVx1_ASAP7_75t_L g7007 ( 
.A(n_4172),
.Y(n_7007)
);

INVx1_ASAP7_75t_SL g7008 ( 
.A(n_9),
.Y(n_7008)
);

CKINVDCx5p33_ASAP7_75t_R g7009 ( 
.A(n_4426),
.Y(n_7009)
);

CKINVDCx5p33_ASAP7_75t_R g7010 ( 
.A(n_3159),
.Y(n_7010)
);

CKINVDCx5p33_ASAP7_75t_R g7011 ( 
.A(n_5827),
.Y(n_7011)
);

INVx1_ASAP7_75t_SL g7012 ( 
.A(n_4512),
.Y(n_7012)
);

CKINVDCx20_ASAP7_75t_R g7013 ( 
.A(n_1128),
.Y(n_7013)
);

CKINVDCx5p33_ASAP7_75t_R g7014 ( 
.A(n_4429),
.Y(n_7014)
);

INVx2_ASAP7_75t_SL g7015 ( 
.A(n_3271),
.Y(n_7015)
);

CKINVDCx5p33_ASAP7_75t_R g7016 ( 
.A(n_5019),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_3812),
.Y(n_7017)
);

INVxp67_ASAP7_75t_L g7018 ( 
.A(n_4453),
.Y(n_7018)
);

INVxp67_ASAP7_75t_L g7019 ( 
.A(n_1436),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_2894),
.Y(n_7020)
);

BUFx3_ASAP7_75t_L g7021 ( 
.A(n_3922),
.Y(n_7021)
);

BUFx5_ASAP7_75t_L g7022 ( 
.A(n_5261),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_1296),
.Y(n_7023)
);

CKINVDCx5p33_ASAP7_75t_R g7024 ( 
.A(n_460),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_5538),
.Y(n_7025)
);

CKINVDCx5p33_ASAP7_75t_R g7026 ( 
.A(n_2292),
.Y(n_7026)
);

INVx1_ASAP7_75t_SL g7027 ( 
.A(n_4406),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_5617),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_5620),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_4502),
.Y(n_7030)
);

CKINVDCx5p33_ASAP7_75t_R g7031 ( 
.A(n_3438),
.Y(n_7031)
);

CKINVDCx5p33_ASAP7_75t_R g7032 ( 
.A(n_6045),
.Y(n_7032)
);

CKINVDCx5p33_ASAP7_75t_R g7033 ( 
.A(n_4524),
.Y(n_7033)
);

INVx2_ASAP7_75t_L g7034 ( 
.A(n_5411),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_4390),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_997),
.Y(n_7036)
);

CKINVDCx5p33_ASAP7_75t_R g7037 ( 
.A(n_1556),
.Y(n_7037)
);

CKINVDCx5p33_ASAP7_75t_R g7038 ( 
.A(n_4938),
.Y(n_7038)
);

CKINVDCx5p33_ASAP7_75t_R g7039 ( 
.A(n_4409),
.Y(n_7039)
);

CKINVDCx5p33_ASAP7_75t_R g7040 ( 
.A(n_2971),
.Y(n_7040)
);

CKINVDCx5p33_ASAP7_75t_R g7041 ( 
.A(n_4895),
.Y(n_7041)
);

CKINVDCx5p33_ASAP7_75t_R g7042 ( 
.A(n_4935),
.Y(n_7042)
);

INVx1_ASAP7_75t_SL g7043 ( 
.A(n_1572),
.Y(n_7043)
);

CKINVDCx14_ASAP7_75t_R g7044 ( 
.A(n_6039),
.Y(n_7044)
);

INVx1_ASAP7_75t_SL g7045 ( 
.A(n_4363),
.Y(n_7045)
);

CKINVDCx16_ASAP7_75t_R g7046 ( 
.A(n_5740),
.Y(n_7046)
);

CKINVDCx5p33_ASAP7_75t_R g7047 ( 
.A(n_419),
.Y(n_7047)
);

HB1xp67_ASAP7_75t_L g7048 ( 
.A(n_5236),
.Y(n_7048)
);

CKINVDCx20_ASAP7_75t_R g7049 ( 
.A(n_4653),
.Y(n_7049)
);

CKINVDCx5p33_ASAP7_75t_R g7050 ( 
.A(n_3373),
.Y(n_7050)
);

CKINVDCx20_ASAP7_75t_R g7051 ( 
.A(n_3629),
.Y(n_7051)
);

CKINVDCx5p33_ASAP7_75t_R g7052 ( 
.A(n_3834),
.Y(n_7052)
);

CKINVDCx5p33_ASAP7_75t_R g7053 ( 
.A(n_5859),
.Y(n_7053)
);

CKINVDCx5p33_ASAP7_75t_R g7054 ( 
.A(n_4978),
.Y(n_7054)
);

CKINVDCx5p33_ASAP7_75t_R g7055 ( 
.A(n_251),
.Y(n_7055)
);

INVx1_ASAP7_75t_L g7056 ( 
.A(n_3604),
.Y(n_7056)
);

CKINVDCx5p33_ASAP7_75t_R g7057 ( 
.A(n_3678),
.Y(n_7057)
);

CKINVDCx5p33_ASAP7_75t_R g7058 ( 
.A(n_1284),
.Y(n_7058)
);

CKINVDCx5p33_ASAP7_75t_R g7059 ( 
.A(n_4544),
.Y(n_7059)
);

CKINVDCx5p33_ASAP7_75t_R g7060 ( 
.A(n_4364),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_3672),
.Y(n_7061)
);

BUFx6f_ASAP7_75t_L g7062 ( 
.A(n_4015),
.Y(n_7062)
);

INVx1_ASAP7_75t_SL g7063 ( 
.A(n_3002),
.Y(n_7063)
);

CKINVDCx16_ASAP7_75t_R g7064 ( 
.A(n_2037),
.Y(n_7064)
);

CKINVDCx5p33_ASAP7_75t_R g7065 ( 
.A(n_359),
.Y(n_7065)
);

CKINVDCx5p33_ASAP7_75t_R g7066 ( 
.A(n_4464),
.Y(n_7066)
);

CKINVDCx5p33_ASAP7_75t_R g7067 ( 
.A(n_3787),
.Y(n_7067)
);

CKINVDCx20_ASAP7_75t_R g7068 ( 
.A(n_2978),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_1877),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_1886),
.Y(n_7070)
);

CKINVDCx5p33_ASAP7_75t_R g7071 ( 
.A(n_4254),
.Y(n_7071)
);

INVx1_ASAP7_75t_L g7072 ( 
.A(n_150),
.Y(n_7072)
);

CKINVDCx5p33_ASAP7_75t_R g7073 ( 
.A(n_5788),
.Y(n_7073)
);

CKINVDCx5p33_ASAP7_75t_R g7074 ( 
.A(n_3575),
.Y(n_7074)
);

CKINVDCx20_ASAP7_75t_R g7075 ( 
.A(n_4459),
.Y(n_7075)
);

CKINVDCx16_ASAP7_75t_R g7076 ( 
.A(n_3224),
.Y(n_7076)
);

CKINVDCx5p33_ASAP7_75t_R g7077 ( 
.A(n_4197),
.Y(n_7077)
);

CKINVDCx5p33_ASAP7_75t_R g7078 ( 
.A(n_1647),
.Y(n_7078)
);

BUFx2_ASAP7_75t_L g7079 ( 
.A(n_3971),
.Y(n_7079)
);

HB1xp67_ASAP7_75t_L g7080 ( 
.A(n_5892),
.Y(n_7080)
);

INVx1_ASAP7_75t_L g7081 ( 
.A(n_1000),
.Y(n_7081)
);

INVx1_ASAP7_75t_L g7082 ( 
.A(n_608),
.Y(n_7082)
);

BUFx10_ASAP7_75t_L g7083 ( 
.A(n_4479),
.Y(n_7083)
);

CKINVDCx5p33_ASAP7_75t_R g7084 ( 
.A(n_2610),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_509),
.Y(n_7085)
);

BUFx6f_ASAP7_75t_L g7086 ( 
.A(n_4595),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_3215),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_1988),
.Y(n_7088)
);

BUFx2_ASAP7_75t_L g7089 ( 
.A(n_4497),
.Y(n_7089)
);

CKINVDCx5p33_ASAP7_75t_R g7090 ( 
.A(n_2756),
.Y(n_7090)
);

CKINVDCx5p33_ASAP7_75t_R g7091 ( 
.A(n_3137),
.Y(n_7091)
);

CKINVDCx5p33_ASAP7_75t_R g7092 ( 
.A(n_2729),
.Y(n_7092)
);

INVx1_ASAP7_75t_SL g7093 ( 
.A(n_4318),
.Y(n_7093)
);

CKINVDCx5p33_ASAP7_75t_R g7094 ( 
.A(n_3396),
.Y(n_7094)
);

INVx1_ASAP7_75t_L g7095 ( 
.A(n_3132),
.Y(n_7095)
);

CKINVDCx5p33_ASAP7_75t_R g7096 ( 
.A(n_1052),
.Y(n_7096)
);

CKINVDCx20_ASAP7_75t_R g7097 ( 
.A(n_2944),
.Y(n_7097)
);

HB1xp67_ASAP7_75t_L g7098 ( 
.A(n_5439),
.Y(n_7098)
);

CKINVDCx5p33_ASAP7_75t_R g7099 ( 
.A(n_3435),
.Y(n_7099)
);

CKINVDCx16_ASAP7_75t_R g7100 ( 
.A(n_4436),
.Y(n_7100)
);

INVx1_ASAP7_75t_L g7101 ( 
.A(n_4379),
.Y(n_7101)
);

CKINVDCx5p33_ASAP7_75t_R g7102 ( 
.A(n_243),
.Y(n_7102)
);

CKINVDCx5p33_ASAP7_75t_R g7103 ( 
.A(n_4407),
.Y(n_7103)
);

CKINVDCx14_ASAP7_75t_R g7104 ( 
.A(n_4487),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_4393),
.Y(n_7105)
);

CKINVDCx5p33_ASAP7_75t_R g7106 ( 
.A(n_5648),
.Y(n_7106)
);

CKINVDCx5p33_ASAP7_75t_R g7107 ( 
.A(n_1528),
.Y(n_7107)
);

INVx1_ASAP7_75t_SL g7108 ( 
.A(n_6069),
.Y(n_7108)
);

CKINVDCx5p33_ASAP7_75t_R g7109 ( 
.A(n_6051),
.Y(n_7109)
);

INVx2_ASAP7_75t_L g7110 ( 
.A(n_5351),
.Y(n_7110)
);

CKINVDCx20_ASAP7_75t_R g7111 ( 
.A(n_4474),
.Y(n_7111)
);

CKINVDCx5p33_ASAP7_75t_R g7112 ( 
.A(n_4714),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_426),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_3005),
.Y(n_7114)
);

INVx2_ASAP7_75t_L g7115 ( 
.A(n_3938),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_4430),
.Y(n_7116)
);

CKINVDCx5p33_ASAP7_75t_R g7117 ( 
.A(n_5790),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_4507),
.Y(n_7118)
);

CKINVDCx5p33_ASAP7_75t_R g7119 ( 
.A(n_28),
.Y(n_7119)
);

CKINVDCx5p33_ASAP7_75t_R g7120 ( 
.A(n_5379),
.Y(n_7120)
);

CKINVDCx5p33_ASAP7_75t_R g7121 ( 
.A(n_903),
.Y(n_7121)
);

BUFx6f_ASAP7_75t_L g7122 ( 
.A(n_4845),
.Y(n_7122)
);

CKINVDCx5p33_ASAP7_75t_R g7123 ( 
.A(n_4057),
.Y(n_7123)
);

CKINVDCx5p33_ASAP7_75t_R g7124 ( 
.A(n_1215),
.Y(n_7124)
);

BUFx10_ASAP7_75t_L g7125 ( 
.A(n_3180),
.Y(n_7125)
);

CKINVDCx20_ASAP7_75t_R g7126 ( 
.A(n_3429),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_661),
.Y(n_7127)
);

CKINVDCx5p33_ASAP7_75t_R g7128 ( 
.A(n_4469),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_4260),
.Y(n_7129)
);

CKINVDCx5p33_ASAP7_75t_R g7130 ( 
.A(n_4661),
.Y(n_7130)
);

CKINVDCx5p33_ASAP7_75t_R g7131 ( 
.A(n_1892),
.Y(n_7131)
);

CKINVDCx5p33_ASAP7_75t_R g7132 ( 
.A(n_3366),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_4486),
.Y(n_7133)
);

CKINVDCx5p33_ASAP7_75t_R g7134 ( 
.A(n_4458),
.Y(n_7134)
);

INVx1_ASAP7_75t_SL g7135 ( 
.A(n_4146),
.Y(n_7135)
);

INVx2_ASAP7_75t_SL g7136 ( 
.A(n_5596),
.Y(n_7136)
);

CKINVDCx5p33_ASAP7_75t_R g7137 ( 
.A(n_1583),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_1611),
.Y(n_7138)
);

CKINVDCx5p33_ASAP7_75t_R g7139 ( 
.A(n_4465),
.Y(n_7139)
);

INVx1_ASAP7_75t_L g7140 ( 
.A(n_1848),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_4494),
.Y(n_7141)
);

CKINVDCx5p33_ASAP7_75t_R g7142 ( 
.A(n_4448),
.Y(n_7142)
);

CKINVDCx20_ASAP7_75t_R g7143 ( 
.A(n_5812),
.Y(n_7143)
);

INVx2_ASAP7_75t_L g7144 ( 
.A(n_4811),
.Y(n_7144)
);

INVx1_ASAP7_75t_L g7145 ( 
.A(n_1947),
.Y(n_7145)
);

INVx2_ASAP7_75t_L g7146 ( 
.A(n_4530),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_1032),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_2849),
.Y(n_7148)
);

CKINVDCx16_ASAP7_75t_R g7149 ( 
.A(n_2437),
.Y(n_7149)
);

CKINVDCx5p33_ASAP7_75t_R g7150 ( 
.A(n_5363),
.Y(n_7150)
);

CKINVDCx16_ASAP7_75t_R g7151 ( 
.A(n_2257),
.Y(n_7151)
);

CKINVDCx5p33_ASAP7_75t_R g7152 ( 
.A(n_463),
.Y(n_7152)
);

CKINVDCx5p33_ASAP7_75t_R g7153 ( 
.A(n_4904),
.Y(n_7153)
);

INVx2_ASAP7_75t_L g7154 ( 
.A(n_398),
.Y(n_7154)
);

CKINVDCx5p33_ASAP7_75t_R g7155 ( 
.A(n_2110),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_2369),
.Y(n_7156)
);

CKINVDCx5p33_ASAP7_75t_R g7157 ( 
.A(n_2431),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_5425),
.Y(n_7158)
);

INVx1_ASAP7_75t_L g7159 ( 
.A(n_1012),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_5445),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_5404),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6044),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_4435),
.Y(n_7163)
);

CKINVDCx16_ASAP7_75t_R g7164 ( 
.A(n_4371),
.Y(n_7164)
);

CKINVDCx5p33_ASAP7_75t_R g7165 ( 
.A(n_4077),
.Y(n_7165)
);

CKINVDCx5p33_ASAP7_75t_R g7166 ( 
.A(n_383),
.Y(n_7166)
);

BUFx2_ASAP7_75t_SL g7167 ( 
.A(n_589),
.Y(n_7167)
);

CKINVDCx5p33_ASAP7_75t_R g7168 ( 
.A(n_1192),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_698),
.Y(n_7169)
);

INVx1_ASAP7_75t_L g7170 ( 
.A(n_2633),
.Y(n_7170)
);

CKINVDCx20_ASAP7_75t_R g7171 ( 
.A(n_1300),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_2244),
.Y(n_7172)
);

CKINVDCx5p33_ASAP7_75t_R g7173 ( 
.A(n_4536),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_4436),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_2158),
.Y(n_7175)
);

CKINVDCx5p33_ASAP7_75t_R g7176 ( 
.A(n_2352),
.Y(n_7176)
);

CKINVDCx5p33_ASAP7_75t_R g7177 ( 
.A(n_636),
.Y(n_7177)
);

CKINVDCx5p33_ASAP7_75t_R g7178 ( 
.A(n_120),
.Y(n_7178)
);

CKINVDCx5p33_ASAP7_75t_R g7179 ( 
.A(n_4513),
.Y(n_7179)
);

CKINVDCx5p33_ASAP7_75t_R g7180 ( 
.A(n_4446),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_1008),
.Y(n_7181)
);

CKINVDCx5p33_ASAP7_75t_R g7182 ( 
.A(n_1764),
.Y(n_7182)
);

BUFx3_ASAP7_75t_L g7183 ( 
.A(n_6060),
.Y(n_7183)
);

CKINVDCx5p33_ASAP7_75t_R g7184 ( 
.A(n_3406),
.Y(n_7184)
);

CKINVDCx5p33_ASAP7_75t_R g7185 ( 
.A(n_3811),
.Y(n_7185)
);

CKINVDCx5p33_ASAP7_75t_R g7186 ( 
.A(n_1657),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_3937),
.Y(n_7187)
);

CKINVDCx5p33_ASAP7_75t_R g7188 ( 
.A(n_4466),
.Y(n_7188)
);

CKINVDCx20_ASAP7_75t_R g7189 ( 
.A(n_380),
.Y(n_7189)
);

CKINVDCx5p33_ASAP7_75t_R g7190 ( 
.A(n_4537),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_5427),
.Y(n_7191)
);

CKINVDCx5p33_ASAP7_75t_R g7192 ( 
.A(n_6047),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_1021),
.Y(n_7193)
);

CKINVDCx20_ASAP7_75t_R g7194 ( 
.A(n_4417),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_3514),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_1491),
.Y(n_7196)
);

INVx1_ASAP7_75t_SL g7197 ( 
.A(n_3826),
.Y(n_7197)
);

BUFx10_ASAP7_75t_L g7198 ( 
.A(n_5361),
.Y(n_7198)
);

CKINVDCx5p33_ASAP7_75t_R g7199 ( 
.A(n_4652),
.Y(n_7199)
);

CKINVDCx5p33_ASAP7_75t_R g7200 ( 
.A(n_2079),
.Y(n_7200)
);

CKINVDCx5p33_ASAP7_75t_R g7201 ( 
.A(n_4307),
.Y(n_7201)
);

CKINVDCx5p33_ASAP7_75t_R g7202 ( 
.A(n_1457),
.Y(n_7202)
);

CKINVDCx20_ASAP7_75t_R g7203 ( 
.A(n_201),
.Y(n_7203)
);

CKINVDCx5p33_ASAP7_75t_R g7204 ( 
.A(n_2752),
.Y(n_7204)
);

CKINVDCx20_ASAP7_75t_R g7205 ( 
.A(n_5977),
.Y(n_7205)
);

CKINVDCx5p33_ASAP7_75t_R g7206 ( 
.A(n_1718),
.Y(n_7206)
);

CKINVDCx5p33_ASAP7_75t_R g7207 ( 
.A(n_5210),
.Y(n_7207)
);

HB1xp67_ASAP7_75t_L g7208 ( 
.A(n_5964),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_517),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_2684),
.Y(n_7210)
);

INVx1_ASAP7_75t_L g7211 ( 
.A(n_4350),
.Y(n_7211)
);

CKINVDCx5p33_ASAP7_75t_R g7212 ( 
.A(n_2173),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_685),
.Y(n_7213)
);

CKINVDCx5p33_ASAP7_75t_R g7214 ( 
.A(n_4483),
.Y(n_7214)
);

BUFx6f_ASAP7_75t_L g7215 ( 
.A(n_2387),
.Y(n_7215)
);

CKINVDCx5p33_ASAP7_75t_R g7216 ( 
.A(n_4355),
.Y(n_7216)
);

CKINVDCx5p33_ASAP7_75t_R g7217 ( 
.A(n_98),
.Y(n_7217)
);

CKINVDCx5p33_ASAP7_75t_R g7218 ( 
.A(n_5444),
.Y(n_7218)
);

CKINVDCx5p33_ASAP7_75t_R g7219 ( 
.A(n_2846),
.Y(n_7219)
);

CKINVDCx5p33_ASAP7_75t_R g7220 ( 
.A(n_4367),
.Y(n_7220)
);

CKINVDCx5p33_ASAP7_75t_R g7221 ( 
.A(n_5789),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_4088),
.Y(n_7222)
);

CKINVDCx5p33_ASAP7_75t_R g7223 ( 
.A(n_4484),
.Y(n_7223)
);

CKINVDCx20_ASAP7_75t_R g7224 ( 
.A(n_548),
.Y(n_7224)
);

CKINVDCx5p33_ASAP7_75t_R g7225 ( 
.A(n_1251),
.Y(n_7225)
);

CKINVDCx5p33_ASAP7_75t_R g7226 ( 
.A(n_3794),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_3044),
.Y(n_7227)
);

CKINVDCx5p33_ASAP7_75t_R g7228 ( 
.A(n_1249),
.Y(n_7228)
);

CKINVDCx5p33_ASAP7_75t_R g7229 ( 
.A(n_4516),
.Y(n_7229)
);

CKINVDCx5p33_ASAP7_75t_R g7230 ( 
.A(n_4293),
.Y(n_7230)
);

CKINVDCx5p33_ASAP7_75t_R g7231 ( 
.A(n_5555),
.Y(n_7231)
);

CKINVDCx5p33_ASAP7_75t_R g7232 ( 
.A(n_3554),
.Y(n_7232)
);

HB1xp67_ASAP7_75t_L g7233 ( 
.A(n_1849),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_4677),
.Y(n_7234)
);

CKINVDCx16_ASAP7_75t_R g7235 ( 
.A(n_5106),
.Y(n_7235)
);

CKINVDCx20_ASAP7_75t_R g7236 ( 
.A(n_4389),
.Y(n_7236)
);

CKINVDCx5p33_ASAP7_75t_R g7237 ( 
.A(n_1787),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_3849),
.Y(n_7238)
);

CKINVDCx20_ASAP7_75t_R g7239 ( 
.A(n_180),
.Y(n_7239)
);

CKINVDCx5p33_ASAP7_75t_R g7240 ( 
.A(n_4115),
.Y(n_7240)
);

CKINVDCx5p33_ASAP7_75t_R g7241 ( 
.A(n_3896),
.Y(n_7241)
);

INVx2_ASAP7_75t_L g7242 ( 
.A(n_4467),
.Y(n_7242)
);

CKINVDCx5p33_ASAP7_75t_R g7243 ( 
.A(n_4495),
.Y(n_7243)
);

INVx2_ASAP7_75t_SL g7244 ( 
.A(n_887),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_5540),
.Y(n_7245)
);

CKINVDCx5p33_ASAP7_75t_R g7246 ( 
.A(n_2988),
.Y(n_7246)
);

CKINVDCx5p33_ASAP7_75t_R g7247 ( 
.A(n_2625),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_4396),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_4442),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_2217),
.Y(n_7250)
);

BUFx10_ASAP7_75t_L g7251 ( 
.A(n_3517),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_4362),
.Y(n_7252)
);

BUFx6f_ASAP7_75t_L g7253 ( 
.A(n_4498),
.Y(n_7253)
);

BUFx2_ASAP7_75t_L g7254 ( 
.A(n_1577),
.Y(n_7254)
);

CKINVDCx5p33_ASAP7_75t_R g7255 ( 
.A(n_3139),
.Y(n_7255)
);

BUFx6f_ASAP7_75t_L g7256 ( 
.A(n_3940),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_13),
.Y(n_7257)
);

CKINVDCx5p33_ASAP7_75t_R g7258 ( 
.A(n_2607),
.Y(n_7258)
);

CKINVDCx5p33_ASAP7_75t_R g7259 ( 
.A(n_3617),
.Y(n_7259)
);

CKINVDCx5p33_ASAP7_75t_R g7260 ( 
.A(n_879),
.Y(n_7260)
);

CKINVDCx5p33_ASAP7_75t_R g7261 ( 
.A(n_3355),
.Y(n_7261)
);

CKINVDCx5p33_ASAP7_75t_R g7262 ( 
.A(n_1362),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_780),
.Y(n_7263)
);

CKINVDCx5p33_ASAP7_75t_R g7264 ( 
.A(n_4372),
.Y(n_7264)
);

BUFx3_ASAP7_75t_L g7265 ( 
.A(n_5194),
.Y(n_7265)
);

BUFx2_ASAP7_75t_L g7266 ( 
.A(n_1710),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_6063),
.Y(n_7267)
);

CKINVDCx5p33_ASAP7_75t_R g7268 ( 
.A(n_4094),
.Y(n_7268)
);

CKINVDCx5p33_ASAP7_75t_R g7269 ( 
.A(n_2723),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_4624),
.Y(n_7270)
);

CKINVDCx5p33_ASAP7_75t_R g7271 ( 
.A(n_490),
.Y(n_7271)
);

CKINVDCx5p33_ASAP7_75t_R g7272 ( 
.A(n_4356),
.Y(n_7272)
);

INVx1_ASAP7_75t_SL g7273 ( 
.A(n_253),
.Y(n_7273)
);

CKINVDCx5p33_ASAP7_75t_R g7274 ( 
.A(n_3924),
.Y(n_7274)
);

CKINVDCx5p33_ASAP7_75t_R g7275 ( 
.A(n_2154),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_401),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_3834),
.Y(n_7277)
);

CKINVDCx5p33_ASAP7_75t_R g7278 ( 
.A(n_3252),
.Y(n_7278)
);

CKINVDCx5p33_ASAP7_75t_R g7279 ( 
.A(n_2628),
.Y(n_7279)
);

BUFx2_ASAP7_75t_L g7280 ( 
.A(n_4771),
.Y(n_7280)
);

CKINVDCx5p33_ASAP7_75t_R g7281 ( 
.A(n_388),
.Y(n_7281)
);

CKINVDCx5p33_ASAP7_75t_R g7282 ( 
.A(n_4140),
.Y(n_7282)
);

CKINVDCx5p33_ASAP7_75t_R g7283 ( 
.A(n_4387),
.Y(n_7283)
);

CKINVDCx20_ASAP7_75t_R g7284 ( 
.A(n_4543),
.Y(n_7284)
);

CKINVDCx5p33_ASAP7_75t_R g7285 ( 
.A(n_3689),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_2324),
.Y(n_7286)
);

HB1xp67_ASAP7_75t_L g7287 ( 
.A(n_4278),
.Y(n_7287)
);

BUFx2_ASAP7_75t_L g7288 ( 
.A(n_4504),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_3773),
.Y(n_7289)
);

CKINVDCx5p33_ASAP7_75t_R g7290 ( 
.A(n_5192),
.Y(n_7290)
);

CKINVDCx5p33_ASAP7_75t_R g7291 ( 
.A(n_2546),
.Y(n_7291)
);

CKINVDCx5p33_ASAP7_75t_R g7292 ( 
.A(n_4548),
.Y(n_7292)
);

CKINVDCx5p33_ASAP7_75t_R g7293 ( 
.A(n_3228),
.Y(n_7293)
);

CKINVDCx5p33_ASAP7_75t_R g7294 ( 
.A(n_4613),
.Y(n_7294)
);

CKINVDCx20_ASAP7_75t_R g7295 ( 
.A(n_4520),
.Y(n_7295)
);

CKINVDCx5p33_ASAP7_75t_R g7296 ( 
.A(n_2128),
.Y(n_7296)
);

CKINVDCx5p33_ASAP7_75t_R g7297 ( 
.A(n_3772),
.Y(n_7297)
);

CKINVDCx20_ASAP7_75t_R g7298 ( 
.A(n_931),
.Y(n_7298)
);

CKINVDCx5p33_ASAP7_75t_R g7299 ( 
.A(n_1010),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_1613),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_224),
.Y(n_7301)
);

INVx2_ASAP7_75t_L g7302 ( 
.A(n_1600),
.Y(n_7302)
);

CKINVDCx5p33_ASAP7_75t_R g7303 ( 
.A(n_1943),
.Y(n_7303)
);

CKINVDCx5p33_ASAP7_75t_R g7304 ( 
.A(n_4512),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_3774),
.Y(n_7305)
);

CKINVDCx5p33_ASAP7_75t_R g7306 ( 
.A(n_1619),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_4141),
.Y(n_7307)
);

CKINVDCx5p33_ASAP7_75t_R g7308 ( 
.A(n_4380),
.Y(n_7308)
);

INVx2_ASAP7_75t_L g7309 ( 
.A(n_5141),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_1756),
.Y(n_7310)
);

INVx1_ASAP7_75t_SL g7311 ( 
.A(n_5489),
.Y(n_7311)
);

CKINVDCx20_ASAP7_75t_R g7312 ( 
.A(n_193),
.Y(n_7312)
);

CKINVDCx20_ASAP7_75t_R g7313 ( 
.A(n_4425),
.Y(n_7313)
);

INVx1_ASAP7_75t_SL g7314 ( 
.A(n_4732),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_4805),
.Y(n_7315)
);

CKINVDCx5p33_ASAP7_75t_R g7316 ( 
.A(n_2533),
.Y(n_7316)
);

CKINVDCx16_ASAP7_75t_R g7317 ( 
.A(n_2425),
.Y(n_7317)
);

CKINVDCx5p33_ASAP7_75t_R g7318 ( 
.A(n_1558),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_1620),
.Y(n_7319)
);

CKINVDCx5p33_ASAP7_75t_R g7320 ( 
.A(n_5183),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_4421),
.Y(n_7321)
);

BUFx6f_ASAP7_75t_L g7322 ( 
.A(n_5850),
.Y(n_7322)
);

CKINVDCx5p33_ASAP7_75t_R g7323 ( 
.A(n_221),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_2678),
.Y(n_7324)
);

CKINVDCx20_ASAP7_75t_R g7325 ( 
.A(n_3421),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_614),
.Y(n_7326)
);

BUFx5_ASAP7_75t_L g7327 ( 
.A(n_2659),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_3588),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_4401),
.Y(n_7329)
);

CKINVDCx5p33_ASAP7_75t_R g7330 ( 
.A(n_5836),
.Y(n_7330)
);

CKINVDCx5p33_ASAP7_75t_R g7331 ( 
.A(n_6036),
.Y(n_7331)
);

CKINVDCx5p33_ASAP7_75t_R g7332 ( 
.A(n_5759),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_1865),
.Y(n_7333)
);

CKINVDCx5p33_ASAP7_75t_R g7334 ( 
.A(n_439),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_191),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_4348),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_5650),
.Y(n_7337)
);

CKINVDCx5p33_ASAP7_75t_R g7338 ( 
.A(n_1810),
.Y(n_7338)
);

CKINVDCx5p33_ASAP7_75t_R g7339 ( 
.A(n_258),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_2617),
.Y(n_7340)
);

CKINVDCx5p33_ASAP7_75t_R g7341 ( 
.A(n_1857),
.Y(n_7341)
);

INVx2_ASAP7_75t_L g7342 ( 
.A(n_2367),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_1624),
.Y(n_7343)
);

CKINVDCx20_ASAP7_75t_R g7344 ( 
.A(n_4559),
.Y(n_7344)
);

CKINVDCx5p33_ASAP7_75t_R g7345 ( 
.A(n_4968),
.Y(n_7345)
);

INVx1_ASAP7_75t_L g7346 ( 
.A(n_6041),
.Y(n_7346)
);

INVx2_ASAP7_75t_L g7347 ( 
.A(n_4441),
.Y(n_7347)
);

CKINVDCx5p33_ASAP7_75t_R g7348 ( 
.A(n_1915),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_5142),
.Y(n_7349)
);

CKINVDCx5p33_ASAP7_75t_R g7350 ( 
.A(n_5877),
.Y(n_7350)
);

CKINVDCx5p33_ASAP7_75t_R g7351 ( 
.A(n_565),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_3562),
.Y(n_7352)
);

INVx2_ASAP7_75t_L g7353 ( 
.A(n_2067),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_520),
.Y(n_7354)
);

CKINVDCx5p33_ASAP7_75t_R g7355 ( 
.A(n_4092),
.Y(n_7355)
);

CKINVDCx5p33_ASAP7_75t_R g7356 ( 
.A(n_1698),
.Y(n_7356)
);

BUFx3_ASAP7_75t_L g7357 ( 
.A(n_4368),
.Y(n_7357)
);

CKINVDCx5p33_ASAP7_75t_R g7358 ( 
.A(n_79),
.Y(n_7358)
);

BUFx5_ASAP7_75t_L g7359 ( 
.A(n_627),
.Y(n_7359)
);

CKINVDCx5p33_ASAP7_75t_R g7360 ( 
.A(n_1923),
.Y(n_7360)
);

CKINVDCx16_ASAP7_75t_R g7361 ( 
.A(n_5922),
.Y(n_7361)
);

CKINVDCx5p33_ASAP7_75t_R g7362 ( 
.A(n_4352),
.Y(n_7362)
);

INVx1_ASAP7_75t_L g7363 ( 
.A(n_1921),
.Y(n_7363)
);

CKINVDCx5p33_ASAP7_75t_R g7364 ( 
.A(n_2876),
.Y(n_7364)
);

INVxp33_ASAP7_75t_L g7365 ( 
.A(n_2162),
.Y(n_7365)
);

INVxp67_ASAP7_75t_L g7366 ( 
.A(n_2242),
.Y(n_7366)
);

CKINVDCx16_ASAP7_75t_R g7367 ( 
.A(n_5311),
.Y(n_7367)
);

INVx1_ASAP7_75t_L g7368 ( 
.A(n_4532),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_956),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_1524),
.Y(n_7370)
);

BUFx2_ASAP7_75t_L g7371 ( 
.A(n_3061),
.Y(n_7371)
);

INVx1_ASAP7_75t_L g7372 ( 
.A(n_4869),
.Y(n_7372)
);

CKINVDCx5p33_ASAP7_75t_R g7373 ( 
.A(n_3104),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_2607),
.Y(n_7374)
);

CKINVDCx5p33_ASAP7_75t_R g7375 ( 
.A(n_4007),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_305),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_2949),
.Y(n_7377)
);

CKINVDCx20_ASAP7_75t_R g7378 ( 
.A(n_5278),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_4388),
.Y(n_7379)
);

CKINVDCx5p33_ASAP7_75t_R g7380 ( 
.A(n_174),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_390),
.Y(n_7381)
);

CKINVDCx5p33_ASAP7_75t_R g7382 ( 
.A(n_5743),
.Y(n_7382)
);

CKINVDCx5p33_ASAP7_75t_R g7383 ( 
.A(n_1096),
.Y(n_7383)
);

CKINVDCx5p33_ASAP7_75t_R g7384 ( 
.A(n_4949),
.Y(n_7384)
);

CKINVDCx20_ASAP7_75t_R g7385 ( 
.A(n_3957),
.Y(n_7385)
);

CKINVDCx5p33_ASAP7_75t_R g7386 ( 
.A(n_5021),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_739),
.Y(n_7387)
);

CKINVDCx5p33_ASAP7_75t_R g7388 ( 
.A(n_5891),
.Y(n_7388)
);

CKINVDCx5p33_ASAP7_75t_R g7389 ( 
.A(n_1591),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_4384),
.Y(n_7390)
);

BUFx6f_ASAP7_75t_L g7391 ( 
.A(n_2667),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_4376),
.Y(n_7392)
);

CKINVDCx20_ASAP7_75t_R g7393 ( 
.A(n_4408),
.Y(n_7393)
);

CKINVDCx5p33_ASAP7_75t_R g7394 ( 
.A(n_1669),
.Y(n_7394)
);

CKINVDCx5p33_ASAP7_75t_R g7395 ( 
.A(n_2006),
.Y(n_7395)
);

CKINVDCx5p33_ASAP7_75t_R g7396 ( 
.A(n_1556),
.Y(n_7396)
);

CKINVDCx5p33_ASAP7_75t_R g7397 ( 
.A(n_818),
.Y(n_7397)
);

CKINVDCx5p33_ASAP7_75t_R g7398 ( 
.A(n_4528),
.Y(n_7398)
);

CKINVDCx20_ASAP7_75t_R g7399 ( 
.A(n_729),
.Y(n_7399)
);

CKINVDCx5p33_ASAP7_75t_R g7400 ( 
.A(n_6053),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_4349),
.Y(n_7401)
);

INVx1_ASAP7_75t_L g7402 ( 
.A(n_3853),
.Y(n_7402)
);

CKINVDCx5p33_ASAP7_75t_R g7403 ( 
.A(n_4776),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_991),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_2520),
.Y(n_7405)
);

CKINVDCx5p33_ASAP7_75t_R g7406 ( 
.A(n_1395),
.Y(n_7406)
);

CKINVDCx5p33_ASAP7_75t_R g7407 ( 
.A(n_1600),
.Y(n_7407)
);

INVx2_ASAP7_75t_SL g7408 ( 
.A(n_4383),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_4646),
.Y(n_7409)
);

CKINVDCx5p33_ASAP7_75t_R g7410 ( 
.A(n_1128),
.Y(n_7410)
);

CKINVDCx5p33_ASAP7_75t_R g7411 ( 
.A(n_3229),
.Y(n_7411)
);

CKINVDCx5p33_ASAP7_75t_R g7412 ( 
.A(n_4350),
.Y(n_7412)
);

CKINVDCx5p33_ASAP7_75t_R g7413 ( 
.A(n_2654),
.Y(n_7413)
);

INVx1_ASAP7_75t_L g7414 ( 
.A(n_2592),
.Y(n_7414)
);

BUFx6f_ASAP7_75t_L g7415 ( 
.A(n_4873),
.Y(n_7415)
);

CKINVDCx20_ASAP7_75t_R g7416 ( 
.A(n_5645),
.Y(n_7416)
);

CKINVDCx5p33_ASAP7_75t_R g7417 ( 
.A(n_4491),
.Y(n_7417)
);

CKINVDCx5p33_ASAP7_75t_R g7418 ( 
.A(n_330),
.Y(n_7418)
);

CKINVDCx20_ASAP7_75t_R g7419 ( 
.A(n_1877),
.Y(n_7419)
);

CKINVDCx5p33_ASAP7_75t_R g7420 ( 
.A(n_4245),
.Y(n_7420)
);

CKINVDCx5p33_ASAP7_75t_R g7421 ( 
.A(n_4514),
.Y(n_7421)
);

CKINVDCx5p33_ASAP7_75t_R g7422 ( 
.A(n_2247),
.Y(n_7422)
);

CKINVDCx5p33_ASAP7_75t_R g7423 ( 
.A(n_163),
.Y(n_7423)
);

INVx1_ASAP7_75t_L g7424 ( 
.A(n_2174),
.Y(n_7424)
);

CKINVDCx5p33_ASAP7_75t_R g7425 ( 
.A(n_5708),
.Y(n_7425)
);

CKINVDCx5p33_ASAP7_75t_R g7426 ( 
.A(n_870),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_4377),
.Y(n_7427)
);

CKINVDCx5p33_ASAP7_75t_R g7428 ( 
.A(n_1637),
.Y(n_7428)
);

BUFx8_ASAP7_75t_SL g7429 ( 
.A(n_3824),
.Y(n_7429)
);

CKINVDCx16_ASAP7_75t_R g7430 ( 
.A(n_350),
.Y(n_7430)
);

CKINVDCx5p33_ASAP7_75t_R g7431 ( 
.A(n_4515),
.Y(n_7431)
);

BUFx3_ASAP7_75t_L g7432 ( 
.A(n_5988),
.Y(n_7432)
);

CKINVDCx5p33_ASAP7_75t_R g7433 ( 
.A(n_4354),
.Y(n_7433)
);

CKINVDCx5p33_ASAP7_75t_R g7434 ( 
.A(n_1660),
.Y(n_7434)
);

CKINVDCx5p33_ASAP7_75t_R g7435 ( 
.A(n_73),
.Y(n_7435)
);

CKINVDCx16_ASAP7_75t_R g7436 ( 
.A(n_4790),
.Y(n_7436)
);

CKINVDCx5p33_ASAP7_75t_R g7437 ( 
.A(n_5103),
.Y(n_7437)
);

INVx2_ASAP7_75t_L g7438 ( 
.A(n_4271),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_3252),
.Y(n_7439)
);

INVx1_ASAP7_75t_SL g7440 ( 
.A(n_3249),
.Y(n_7440)
);

CKINVDCx5p33_ASAP7_75t_R g7441 ( 
.A(n_4386),
.Y(n_7441)
);

CKINVDCx5p33_ASAP7_75t_R g7442 ( 
.A(n_2409),
.Y(n_7442)
);

CKINVDCx5p33_ASAP7_75t_R g7443 ( 
.A(n_541),
.Y(n_7443)
);

CKINVDCx5p33_ASAP7_75t_R g7444 ( 
.A(n_2966),
.Y(n_7444)
);

BUFx8_ASAP7_75t_SL g7445 ( 
.A(n_4027),
.Y(n_7445)
);

CKINVDCx5p33_ASAP7_75t_R g7446 ( 
.A(n_4346),
.Y(n_7446)
);

CKINVDCx5p33_ASAP7_75t_R g7447 ( 
.A(n_4541),
.Y(n_7447)
);

CKINVDCx5p33_ASAP7_75t_R g7448 ( 
.A(n_575),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_729),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_2979),
.Y(n_7450)
);

BUFx6f_ASAP7_75t_L g7451 ( 
.A(n_4550),
.Y(n_7451)
);

CKINVDCx5p33_ASAP7_75t_R g7452 ( 
.A(n_3579),
.Y(n_7452)
);

CKINVDCx5p33_ASAP7_75t_R g7453 ( 
.A(n_4177),
.Y(n_7453)
);

CKINVDCx5p33_ASAP7_75t_R g7454 ( 
.A(n_4118),
.Y(n_7454)
);

BUFx2_ASAP7_75t_L g7455 ( 
.A(n_3144),
.Y(n_7455)
);

CKINVDCx20_ASAP7_75t_R g7456 ( 
.A(n_5205),
.Y(n_7456)
);

CKINVDCx5p33_ASAP7_75t_R g7457 ( 
.A(n_3546),
.Y(n_7457)
);

INVx2_ASAP7_75t_SL g7458 ( 
.A(n_4526),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_76),
.Y(n_7459)
);

BUFx10_ASAP7_75t_L g7460 ( 
.A(n_5228),
.Y(n_7460)
);

INVx1_ASAP7_75t_SL g7461 ( 
.A(n_5546),
.Y(n_7461)
);

CKINVDCx5p33_ASAP7_75t_R g7462 ( 
.A(n_6052),
.Y(n_7462)
);

BUFx3_ASAP7_75t_L g7463 ( 
.A(n_5927),
.Y(n_7463)
);

INVx1_ASAP7_75t_SL g7464 ( 
.A(n_4299),
.Y(n_7464)
);

CKINVDCx5p33_ASAP7_75t_R g7465 ( 
.A(n_3960),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_2799),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_3011),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_3143),
.Y(n_7468)
);

BUFx3_ASAP7_75t_L g7469 ( 
.A(n_4423),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_3046),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_3243),
.Y(n_7471)
);

CKINVDCx5p33_ASAP7_75t_R g7472 ( 
.A(n_4194),
.Y(n_7472)
);

CKINVDCx5p33_ASAP7_75t_R g7473 ( 
.A(n_5532),
.Y(n_7473)
);

CKINVDCx5p33_ASAP7_75t_R g7474 ( 
.A(n_3261),
.Y(n_7474)
);

CKINVDCx5p33_ASAP7_75t_R g7475 ( 
.A(n_4035),
.Y(n_7475)
);

BUFx3_ASAP7_75t_L g7476 ( 
.A(n_4166),
.Y(n_7476)
);

INVxp33_ASAP7_75t_R g7477 ( 
.A(n_4529),
.Y(n_7477)
);

CKINVDCx5p33_ASAP7_75t_R g7478 ( 
.A(n_4631),
.Y(n_7478)
);

CKINVDCx20_ASAP7_75t_R g7479 ( 
.A(n_6061),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_2647),
.Y(n_7480)
);

CKINVDCx20_ASAP7_75t_R g7481 ( 
.A(n_2653),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_1927),
.Y(n_7482)
);

CKINVDCx5p33_ASAP7_75t_R g7483 ( 
.A(n_4519),
.Y(n_7483)
);

CKINVDCx5p33_ASAP7_75t_R g7484 ( 
.A(n_2433),
.Y(n_7484)
);

INVx1_ASAP7_75t_L g7485 ( 
.A(n_2611),
.Y(n_7485)
);

BUFx2_ASAP7_75t_L g7486 ( 
.A(n_3696),
.Y(n_7486)
);

INVx1_ASAP7_75t_SL g7487 ( 
.A(n_5305),
.Y(n_7487)
);

CKINVDCx5p33_ASAP7_75t_R g7488 ( 
.A(n_211),
.Y(n_7488)
);

CKINVDCx5p33_ASAP7_75t_R g7489 ( 
.A(n_1630),
.Y(n_7489)
);

BUFx3_ASAP7_75t_L g7490 ( 
.A(n_453),
.Y(n_7490)
);

BUFx3_ASAP7_75t_L g7491 ( 
.A(n_5819),
.Y(n_7491)
);

CKINVDCx5p33_ASAP7_75t_R g7492 ( 
.A(n_2124),
.Y(n_7492)
);

CKINVDCx5p33_ASAP7_75t_R g7493 ( 
.A(n_5786),
.Y(n_7493)
);

INVx1_ASAP7_75t_SL g7494 ( 
.A(n_1803),
.Y(n_7494)
);

BUFx5_ASAP7_75t_L g7495 ( 
.A(n_5615),
.Y(n_7495)
);

INVx2_ASAP7_75t_SL g7496 ( 
.A(n_2337),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_3157),
.Y(n_7497)
);

CKINVDCx5p33_ASAP7_75t_R g7498 ( 
.A(n_4420),
.Y(n_7498)
);

CKINVDCx5p33_ASAP7_75t_R g7499 ( 
.A(n_5661),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_2375),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_1575),
.Y(n_7501)
);

INVx2_ASAP7_75t_L g7502 ( 
.A(n_4176),
.Y(n_7502)
);

CKINVDCx5p33_ASAP7_75t_R g7503 ( 
.A(n_4528),
.Y(n_7503)
);

CKINVDCx5p33_ASAP7_75t_R g7504 ( 
.A(n_4432),
.Y(n_7504)
);

BUFx8_ASAP7_75t_SL g7505 ( 
.A(n_4235),
.Y(n_7505)
);

CKINVDCx5p33_ASAP7_75t_R g7506 ( 
.A(n_5865),
.Y(n_7506)
);

CKINVDCx5p33_ASAP7_75t_R g7507 ( 
.A(n_5686),
.Y(n_7507)
);

CKINVDCx5p33_ASAP7_75t_R g7508 ( 
.A(n_4002),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_4427),
.Y(n_7509)
);

INVx1_ASAP7_75t_L g7510 ( 
.A(n_3021),
.Y(n_7510)
);

CKINVDCx5p33_ASAP7_75t_R g7511 ( 
.A(n_2804),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_1856),
.Y(n_7512)
);

BUFx3_ASAP7_75t_L g7513 ( 
.A(n_3144),
.Y(n_7513)
);

INVx2_ASAP7_75t_L g7514 ( 
.A(n_4264),
.Y(n_7514)
);

CKINVDCx5p33_ASAP7_75t_R g7515 ( 
.A(n_4347),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_2306),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_4447),
.Y(n_7517)
);

CKINVDCx20_ASAP7_75t_R g7518 ( 
.A(n_3305),
.Y(n_7518)
);

CKINVDCx5p33_ASAP7_75t_R g7519 ( 
.A(n_411),
.Y(n_7519)
);

CKINVDCx16_ASAP7_75t_R g7520 ( 
.A(n_2282),
.Y(n_7520)
);

BUFx6f_ASAP7_75t_L g7521 ( 
.A(n_3456),
.Y(n_7521)
);

CKINVDCx5p33_ASAP7_75t_R g7522 ( 
.A(n_2207),
.Y(n_7522)
);

CKINVDCx5p33_ASAP7_75t_R g7523 ( 
.A(n_4412),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_2532),
.Y(n_7524)
);

CKINVDCx5p33_ASAP7_75t_R g7525 ( 
.A(n_4063),
.Y(n_7525)
);

INVx1_ASAP7_75t_L g7526 ( 
.A(n_3691),
.Y(n_7526)
);

CKINVDCx5p33_ASAP7_75t_R g7527 ( 
.A(n_4158),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_727),
.Y(n_7528)
);

CKINVDCx20_ASAP7_75t_R g7529 ( 
.A(n_6035),
.Y(n_7529)
);

INVx2_ASAP7_75t_L g7530 ( 
.A(n_4397),
.Y(n_7530)
);

CKINVDCx5p33_ASAP7_75t_R g7531 ( 
.A(n_5374),
.Y(n_7531)
);

INVx1_ASAP7_75t_L g7532 ( 
.A(n_5659),
.Y(n_7532)
);

CKINVDCx5p33_ASAP7_75t_R g7533 ( 
.A(n_2890),
.Y(n_7533)
);

CKINVDCx16_ASAP7_75t_R g7534 ( 
.A(n_4505),
.Y(n_7534)
);

HB1xp67_ASAP7_75t_L g7535 ( 
.A(n_1501),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_172),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_4315),
.Y(n_7537)
);

INVx1_ASAP7_75t_L g7538 ( 
.A(n_1486),
.Y(n_7538)
);

CKINVDCx5p33_ASAP7_75t_R g7539 ( 
.A(n_3951),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_3963),
.Y(n_7540)
);

BUFx3_ASAP7_75t_L g7541 ( 
.A(n_348),
.Y(n_7541)
);

CKINVDCx5p33_ASAP7_75t_R g7542 ( 
.A(n_1595),
.Y(n_7542)
);

CKINVDCx5p33_ASAP7_75t_R g7543 ( 
.A(n_1985),
.Y(n_7543)
);

BUFx2_ASAP7_75t_L g7544 ( 
.A(n_4153),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_3735),
.Y(n_7545)
);

CKINVDCx5p33_ASAP7_75t_R g7546 ( 
.A(n_6333),
.Y(n_7546)
);

CKINVDCx20_ASAP7_75t_R g7547 ( 
.A(n_6116),
.Y(n_7547)
);

CKINVDCx5p33_ASAP7_75t_R g7548 ( 
.A(n_6251),
.Y(n_7548)
);

CKINVDCx5p33_ASAP7_75t_R g7549 ( 
.A(n_6449),
.Y(n_7549)
);

CKINVDCx20_ASAP7_75t_R g7550 ( 
.A(n_6203),
.Y(n_7550)
);

CKINVDCx5p33_ASAP7_75t_R g7551 ( 
.A(n_6484),
.Y(n_7551)
);

CKINVDCx5p33_ASAP7_75t_R g7552 ( 
.A(n_7429),
.Y(n_7552)
);

BUFx6f_ASAP7_75t_L g7553 ( 
.A(n_6193),
.Y(n_7553)
);

NOR2xp67_ASAP7_75t_L g7554 ( 
.A(n_6227),
.B(n_0),
.Y(n_7554)
);

CKINVDCx5p33_ASAP7_75t_R g7555 ( 
.A(n_7445),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_6130),
.Y(n_7556)
);

CKINVDCx5p33_ASAP7_75t_R g7557 ( 
.A(n_7505),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_6130),
.Y(n_7558)
);

CKINVDCx5p33_ASAP7_75t_R g7559 ( 
.A(n_6649),
.Y(n_7559)
);

HB1xp67_ASAP7_75t_L g7560 ( 
.A(n_6126),
.Y(n_7560)
);

INVx2_ASAP7_75t_L g7561 ( 
.A(n_6130),
.Y(n_7561)
);

CKINVDCx5p33_ASAP7_75t_R g7562 ( 
.A(n_6082),
.Y(n_7562)
);

CKINVDCx5p33_ASAP7_75t_R g7563 ( 
.A(n_6086),
.Y(n_7563)
);

CKINVDCx5p33_ASAP7_75t_R g7564 ( 
.A(n_6102),
.Y(n_7564)
);

CKINVDCx20_ASAP7_75t_R g7565 ( 
.A(n_6205),
.Y(n_7565)
);

INVx1_ASAP7_75t_L g7566 ( 
.A(n_6130),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_6130),
.Y(n_7567)
);

INVx2_ASAP7_75t_L g7568 ( 
.A(n_6177),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_6177),
.Y(n_7569)
);

CKINVDCx5p33_ASAP7_75t_R g7570 ( 
.A(n_6105),
.Y(n_7570)
);

NOR2xp67_ASAP7_75t_L g7571 ( 
.A(n_6423),
.B(n_0),
.Y(n_7571)
);

CKINVDCx5p33_ASAP7_75t_R g7572 ( 
.A(n_6115),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_6177),
.Y(n_7573)
);

CKINVDCx5p33_ASAP7_75t_R g7574 ( 
.A(n_6119),
.Y(n_7574)
);

CKINVDCx20_ASAP7_75t_R g7575 ( 
.A(n_6234),
.Y(n_7575)
);

INVx2_ASAP7_75t_L g7576 ( 
.A(n_6177),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_6177),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_6241),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_6241),
.Y(n_7579)
);

CKINVDCx5p33_ASAP7_75t_R g7580 ( 
.A(n_6120),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_6241),
.Y(n_7581)
);

NOR2xp67_ASAP7_75t_L g7582 ( 
.A(n_6445),
.B(n_1),
.Y(n_7582)
);

CKINVDCx5p33_ASAP7_75t_R g7583 ( 
.A(n_6123),
.Y(n_7583)
);

CKINVDCx5p33_ASAP7_75t_R g7584 ( 
.A(n_6128),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_6241),
.Y(n_7585)
);

CKINVDCx5p33_ASAP7_75t_R g7586 ( 
.A(n_6131),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_6241),
.Y(n_7587)
);

CKINVDCx5p33_ASAP7_75t_R g7588 ( 
.A(n_6132),
.Y(n_7588)
);

CKINVDCx5p33_ASAP7_75t_R g7589 ( 
.A(n_6138),
.Y(n_7589)
);

INVx1_ASAP7_75t_L g7590 ( 
.A(n_6270),
.Y(n_7590)
);

CKINVDCx16_ASAP7_75t_R g7591 ( 
.A(n_6415),
.Y(n_7591)
);

CKINVDCx14_ASAP7_75t_R g7592 ( 
.A(n_6402),
.Y(n_7592)
);

CKINVDCx5p33_ASAP7_75t_R g7593 ( 
.A(n_6149),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_6270),
.Y(n_7594)
);

CKINVDCx5p33_ASAP7_75t_R g7595 ( 
.A(n_6153),
.Y(n_7595)
);

INVx2_ASAP7_75t_L g7596 ( 
.A(n_6270),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_6270),
.Y(n_7597)
);

CKINVDCx5p33_ASAP7_75t_R g7598 ( 
.A(n_6154),
.Y(n_7598)
);

CKINVDCx5p33_ASAP7_75t_R g7599 ( 
.A(n_6155),
.Y(n_7599)
);

INVx1_ASAP7_75t_L g7600 ( 
.A(n_6270),
.Y(n_7600)
);

CKINVDCx5p33_ASAP7_75t_R g7601 ( 
.A(n_6163),
.Y(n_7601)
);

INVx1_ASAP7_75t_L g7602 ( 
.A(n_6309),
.Y(n_7602)
);

INVx1_ASAP7_75t_L g7603 ( 
.A(n_6309),
.Y(n_7603)
);

INVx2_ASAP7_75t_L g7604 ( 
.A(n_6309),
.Y(n_7604)
);

INVx2_ASAP7_75t_L g7605 ( 
.A(n_6309),
.Y(n_7605)
);

CKINVDCx20_ASAP7_75t_R g7606 ( 
.A(n_6319),
.Y(n_7606)
);

CKINVDCx5p33_ASAP7_75t_R g7607 ( 
.A(n_6174),
.Y(n_7607)
);

INVx1_ASAP7_75t_L g7608 ( 
.A(n_6309),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_6381),
.Y(n_7609)
);

CKINVDCx14_ASAP7_75t_R g7610 ( 
.A(n_6490),
.Y(n_7610)
);

INVx1_ASAP7_75t_L g7611 ( 
.A(n_6381),
.Y(n_7611)
);

CKINVDCx5p33_ASAP7_75t_R g7612 ( 
.A(n_6182),
.Y(n_7612)
);

INVxp67_ASAP7_75t_SL g7613 ( 
.A(n_6676),
.Y(n_7613)
);

INVx2_ASAP7_75t_L g7614 ( 
.A(n_6381),
.Y(n_7614)
);

CKINVDCx5p33_ASAP7_75t_R g7615 ( 
.A(n_6184),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_6381),
.Y(n_7616)
);

INVx2_ASAP7_75t_L g7617 ( 
.A(n_6381),
.Y(n_7617)
);

BUFx6f_ASAP7_75t_L g7618 ( 
.A(n_6193),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_6699),
.Y(n_7619)
);

CKINVDCx5p33_ASAP7_75t_R g7620 ( 
.A(n_6188),
.Y(n_7620)
);

CKINVDCx5p33_ASAP7_75t_R g7621 ( 
.A(n_6207),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_6699),
.Y(n_7622)
);

CKINVDCx20_ASAP7_75t_R g7623 ( 
.A(n_6466),
.Y(n_7623)
);

CKINVDCx20_ASAP7_75t_R g7624 ( 
.A(n_6502),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_6699),
.Y(n_7625)
);

OR2x2_ASAP7_75t_L g7626 ( 
.A(n_6093),
.B(n_1),
.Y(n_7626)
);

INVxp67_ASAP7_75t_L g7627 ( 
.A(n_6121),
.Y(n_7627)
);

CKINVDCx20_ASAP7_75t_R g7628 ( 
.A(n_6583),
.Y(n_7628)
);

BUFx3_ASAP7_75t_L g7629 ( 
.A(n_6312),
.Y(n_7629)
);

CKINVDCx5p33_ASAP7_75t_R g7630 ( 
.A(n_6214),
.Y(n_7630)
);

NOR2xp67_ASAP7_75t_L g7631 ( 
.A(n_6511),
.B(n_2),
.Y(n_7631)
);

CKINVDCx5p33_ASAP7_75t_R g7632 ( 
.A(n_6216),
.Y(n_7632)
);

CKINVDCx5p33_ASAP7_75t_R g7633 ( 
.A(n_6218),
.Y(n_7633)
);

CKINVDCx5p33_ASAP7_75t_R g7634 ( 
.A(n_6220),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_6699),
.Y(n_7635)
);

CKINVDCx5p33_ASAP7_75t_R g7636 ( 
.A(n_6223),
.Y(n_7636)
);

CKINVDCx5p33_ASAP7_75t_R g7637 ( 
.A(n_6235),
.Y(n_7637)
);

CKINVDCx5p33_ASAP7_75t_R g7638 ( 
.A(n_6236),
.Y(n_7638)
);

BUFx6f_ASAP7_75t_L g7639 ( 
.A(n_6193),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_6699),
.Y(n_7640)
);

CKINVDCx5p33_ASAP7_75t_R g7641 ( 
.A(n_6249),
.Y(n_7641)
);

CKINVDCx20_ASAP7_75t_R g7642 ( 
.A(n_6632),
.Y(n_7642)
);

CKINVDCx5p33_ASAP7_75t_R g7643 ( 
.A(n_6255),
.Y(n_7643)
);

CKINVDCx5p33_ASAP7_75t_R g7644 ( 
.A(n_6265),
.Y(n_7644)
);

INVx1_ASAP7_75t_L g7645 ( 
.A(n_7327),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7327),
.Y(n_7646)
);

CKINVDCx5p33_ASAP7_75t_R g7647 ( 
.A(n_6286),
.Y(n_7647)
);

CKINVDCx5p33_ASAP7_75t_R g7648 ( 
.A(n_6298),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7327),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7327),
.Y(n_7650)
);

CKINVDCx5p33_ASAP7_75t_R g7651 ( 
.A(n_6311),
.Y(n_7651)
);

NOR2xp67_ASAP7_75t_L g7652 ( 
.A(n_6541),
.B(n_2),
.Y(n_7652)
);

CKINVDCx5p33_ASAP7_75t_R g7653 ( 
.A(n_6315),
.Y(n_7653)
);

INVx1_ASAP7_75t_L g7654 ( 
.A(n_7327),
.Y(n_7654)
);

CKINVDCx5p33_ASAP7_75t_R g7655 ( 
.A(n_6317),
.Y(n_7655)
);

CKINVDCx5p33_ASAP7_75t_R g7656 ( 
.A(n_6321),
.Y(n_7656)
);

CKINVDCx5p33_ASAP7_75t_R g7657 ( 
.A(n_6327),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7359),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_7359),
.Y(n_7659)
);

BUFx5_ASAP7_75t_L g7660 ( 
.A(n_6085),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_7359),
.Y(n_7661)
);

INVx2_ASAP7_75t_L g7662 ( 
.A(n_7359),
.Y(n_7662)
);

INVx1_ASAP7_75t_L g7663 ( 
.A(n_7359),
.Y(n_7663)
);

CKINVDCx5p33_ASAP7_75t_R g7664 ( 
.A(n_6350),
.Y(n_7664)
);

CKINVDCx5p33_ASAP7_75t_R g7665 ( 
.A(n_6353),
.Y(n_7665)
);

CKINVDCx5p33_ASAP7_75t_R g7666 ( 
.A(n_6356),
.Y(n_7666)
);

CKINVDCx5p33_ASAP7_75t_R g7667 ( 
.A(n_6362),
.Y(n_7667)
);

BUFx10_ASAP7_75t_L g7668 ( 
.A(n_7535),
.Y(n_7668)
);

INVx1_ASAP7_75t_L g7669 ( 
.A(n_6087),
.Y(n_7669)
);

CKINVDCx5p33_ASAP7_75t_R g7670 ( 
.A(n_6366),
.Y(n_7670)
);

CKINVDCx5p33_ASAP7_75t_R g7671 ( 
.A(n_6368),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_6087),
.Y(n_7672)
);

CKINVDCx5p33_ASAP7_75t_R g7673 ( 
.A(n_6385),
.Y(n_7673)
);

CKINVDCx5p33_ASAP7_75t_R g7674 ( 
.A(n_6391),
.Y(n_7674)
);

INVx1_ASAP7_75t_L g7675 ( 
.A(n_6087),
.Y(n_7675)
);

CKINVDCx5p33_ASAP7_75t_R g7676 ( 
.A(n_6407),
.Y(n_7676)
);

CKINVDCx5p33_ASAP7_75t_R g7677 ( 
.A(n_6434),
.Y(n_7677)
);

INVx1_ASAP7_75t_L g7678 ( 
.A(n_6090),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_6090),
.Y(n_7679)
);

CKINVDCx16_ASAP7_75t_R g7680 ( 
.A(n_6438),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_6090),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_6108),
.Y(n_7682)
);

CKINVDCx14_ASAP7_75t_R g7683 ( 
.A(n_7104),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_6108),
.Y(n_7684)
);

CKINVDCx5p33_ASAP7_75t_R g7685 ( 
.A(n_6436),
.Y(n_7685)
);

INVx1_ASAP7_75t_L g7686 ( 
.A(n_6108),
.Y(n_7686)
);

INVx1_ASAP7_75t_L g7687 ( 
.A(n_6113),
.Y(n_7687)
);

CKINVDCx5p33_ASAP7_75t_R g7688 ( 
.A(n_6442),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_6113),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_6113),
.Y(n_7690)
);

HB1xp67_ASAP7_75t_L g7691 ( 
.A(n_7534),
.Y(n_7691)
);

INVx1_ASAP7_75t_L g7692 ( 
.A(n_6151),
.Y(n_7692)
);

BUFx3_ASAP7_75t_L g7693 ( 
.A(n_6312),
.Y(n_7693)
);

CKINVDCx16_ASAP7_75t_R g7694 ( 
.A(n_6473),
.Y(n_7694)
);

CKINVDCx20_ASAP7_75t_R g7695 ( 
.A(n_6694),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_6151),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_6151),
.Y(n_7697)
);

CKINVDCx5p33_ASAP7_75t_R g7698 ( 
.A(n_6448),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_6167),
.Y(n_7699)
);

NOR2xp67_ASAP7_75t_L g7700 ( 
.A(n_6666),
.B(n_3),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_6167),
.Y(n_7701)
);

INVx1_ASAP7_75t_L g7702 ( 
.A(n_6167),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_6267),
.Y(n_7703)
);

CKINVDCx5p33_ASAP7_75t_R g7704 ( 
.A(n_6453),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_6267),
.Y(n_7705)
);

INVxp67_ASAP7_75t_L g7706 ( 
.A(n_6324),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_6267),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_6330),
.Y(n_7708)
);

CKINVDCx20_ASAP7_75t_R g7709 ( 
.A(n_6862),
.Y(n_7709)
);

CKINVDCx14_ASAP7_75t_R g7710 ( 
.A(n_6477),
.Y(n_7710)
);

CKINVDCx5p33_ASAP7_75t_R g7711 ( 
.A(n_6460),
.Y(n_7711)
);

CKINVDCx20_ASAP7_75t_R g7712 ( 
.A(n_6999),
.Y(n_7712)
);

CKINVDCx5p33_ASAP7_75t_R g7713 ( 
.A(n_6468),
.Y(n_7713)
);

CKINVDCx5p33_ASAP7_75t_R g7714 ( 
.A(n_6483),
.Y(n_7714)
);

INVxp67_ASAP7_75t_SL g7715 ( 
.A(n_7048),
.Y(n_7715)
);

CKINVDCx5p33_ASAP7_75t_R g7716 ( 
.A(n_6489),
.Y(n_7716)
);

OR2x2_ASAP7_75t_L g7717 ( 
.A(n_6667),
.B(n_4),
.Y(n_7717)
);

CKINVDCx5p33_ASAP7_75t_R g7718 ( 
.A(n_6522),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_6330),
.Y(n_7719)
);

CKINVDCx5p33_ASAP7_75t_R g7720 ( 
.A(n_6534),
.Y(n_7720)
);

CKINVDCx5p33_ASAP7_75t_R g7721 ( 
.A(n_6542),
.Y(n_7721)
);

CKINVDCx5p33_ASAP7_75t_R g7722 ( 
.A(n_6560),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_6330),
.Y(n_7723)
);

CKINVDCx5p33_ASAP7_75t_R g7724 ( 
.A(n_6564),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_6357),
.Y(n_7725)
);

XNOR2xp5_ASAP7_75t_L g7726 ( 
.A(n_6076),
.B(n_4),
.Y(n_7726)
);

BUFx3_ASAP7_75t_L g7727 ( 
.A(n_6517),
.Y(n_7727)
);

INVx1_ASAP7_75t_SL g7728 ( 
.A(n_6731),
.Y(n_7728)
);

NOR2xp67_ASAP7_75t_L g7729 ( 
.A(n_6735),
.B(n_5),
.Y(n_7729)
);

NOR2xp67_ASAP7_75t_L g7730 ( 
.A(n_6781),
.B(n_5),
.Y(n_7730)
);

CKINVDCx5p33_ASAP7_75t_R g7731 ( 
.A(n_6570),
.Y(n_7731)
);

CKINVDCx5p33_ASAP7_75t_R g7732 ( 
.A(n_6572),
.Y(n_7732)
);

INVxp67_ASAP7_75t_L g7733 ( 
.A(n_6945),
.Y(n_7733)
);

CKINVDCx14_ASAP7_75t_R g7734 ( 
.A(n_6498),
.Y(n_7734)
);

CKINVDCx16_ASAP7_75t_R g7735 ( 
.A(n_6549),
.Y(n_7735)
);

INVx1_ASAP7_75t_L g7736 ( 
.A(n_6357),
.Y(n_7736)
);

CKINVDCx5p33_ASAP7_75t_R g7737 ( 
.A(n_6593),
.Y(n_7737)
);

CKINVDCx5p33_ASAP7_75t_R g7738 ( 
.A(n_6597),
.Y(n_7738)
);

CKINVDCx5p33_ASAP7_75t_R g7739 ( 
.A(n_6605),
.Y(n_7739)
);

CKINVDCx20_ASAP7_75t_R g7740 ( 
.A(n_7049),
.Y(n_7740)
);

INVx1_ASAP7_75t_L g7741 ( 
.A(n_6357),
.Y(n_7741)
);

INVx1_ASAP7_75t_L g7742 ( 
.A(n_6535),
.Y(n_7742)
);

CKINVDCx5p33_ASAP7_75t_R g7743 ( 
.A(n_6609),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_6535),
.Y(n_7744)
);

CKINVDCx5p33_ASAP7_75t_R g7745 ( 
.A(n_6613),
.Y(n_7745)
);

BUFx6f_ASAP7_75t_L g7746 ( 
.A(n_6334),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_6535),
.Y(n_7747)
);

CKINVDCx5p33_ASAP7_75t_R g7748 ( 
.A(n_6614),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_6594),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_6594),
.Y(n_7750)
);

INVx1_ASAP7_75t_L g7751 ( 
.A(n_6594),
.Y(n_7751)
);

CKINVDCx20_ASAP7_75t_R g7752 ( 
.A(n_7529),
.Y(n_7752)
);

CKINVDCx5p33_ASAP7_75t_R g7753 ( 
.A(n_6622),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_6638),
.Y(n_7754)
);

BUFx2_ASAP7_75t_L g7755 ( 
.A(n_7079),
.Y(n_7755)
);

INVx1_ASAP7_75t_SL g7756 ( 
.A(n_7089),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_6638),
.Y(n_7757)
);

INVx1_ASAP7_75t_L g7758 ( 
.A(n_6638),
.Y(n_7758)
);

CKINVDCx5p33_ASAP7_75t_R g7759 ( 
.A(n_6631),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_6692),
.Y(n_7760)
);

CKINVDCx5p33_ASAP7_75t_R g7761 ( 
.A(n_6633),
.Y(n_7761)
);

BUFx6f_ASAP7_75t_L g7762 ( 
.A(n_6334),
.Y(n_7762)
);

CKINVDCx5p33_ASAP7_75t_R g7763 ( 
.A(n_6637),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_6692),
.Y(n_7764)
);

CKINVDCx5p33_ASAP7_75t_R g7765 ( 
.A(n_6643),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_6692),
.Y(n_7766)
);

INVx2_ASAP7_75t_L g7767 ( 
.A(n_6807),
.Y(n_7767)
);

CKINVDCx5p33_ASAP7_75t_R g7768 ( 
.A(n_6652),
.Y(n_7768)
);

CKINVDCx5p33_ASAP7_75t_R g7769 ( 
.A(n_6661),
.Y(n_7769)
);

CKINVDCx5p33_ASAP7_75t_R g7770 ( 
.A(n_6662),
.Y(n_7770)
);

CKINVDCx5p33_ASAP7_75t_R g7771 ( 
.A(n_6670),
.Y(n_7771)
);

CKINVDCx16_ASAP7_75t_R g7772 ( 
.A(n_6552),
.Y(n_7772)
);

CKINVDCx16_ASAP7_75t_R g7773 ( 
.A(n_6634),
.Y(n_7773)
);

CKINVDCx5p33_ASAP7_75t_R g7774 ( 
.A(n_6677),
.Y(n_7774)
);

CKINVDCx20_ASAP7_75t_R g7775 ( 
.A(n_7143),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_6807),
.Y(n_7776)
);

CKINVDCx5p33_ASAP7_75t_R g7777 ( 
.A(n_6683),
.Y(n_7777)
);

NOR2xp67_ASAP7_75t_L g7778 ( 
.A(n_7018),
.B(n_6),
.Y(n_7778)
);

CKINVDCx5p33_ASAP7_75t_R g7779 ( 
.A(n_6693),
.Y(n_7779)
);

CKINVDCx5p33_ASAP7_75t_R g7780 ( 
.A(n_6698),
.Y(n_7780)
);

BUFx10_ASAP7_75t_L g7781 ( 
.A(n_6495),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_6807),
.Y(n_7782)
);

CKINVDCx5p33_ASAP7_75t_R g7783 ( 
.A(n_6712),
.Y(n_7783)
);

HB1xp67_ASAP7_75t_L g7784 ( 
.A(n_6758),
.Y(n_7784)
);

BUFx6f_ASAP7_75t_L g7785 ( 
.A(n_6334),
.Y(n_7785)
);

CKINVDCx5p33_ASAP7_75t_R g7786 ( 
.A(n_6718),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_6912),
.Y(n_7787)
);

BUFx8_ASAP7_75t_SL g7788 ( 
.A(n_7254),
.Y(n_7788)
);

CKINVDCx5p33_ASAP7_75t_R g7789 ( 
.A(n_6743),
.Y(n_7789)
);

OR2x2_ASAP7_75t_L g7790 ( 
.A(n_7266),
.B(n_6),
.Y(n_7790)
);

CKINVDCx5p33_ASAP7_75t_R g7791 ( 
.A(n_6745),
.Y(n_7791)
);

CKINVDCx5p33_ASAP7_75t_R g7792 ( 
.A(n_6752),
.Y(n_7792)
);

CKINVDCx5p33_ASAP7_75t_R g7793 ( 
.A(n_6754),
.Y(n_7793)
);

CKINVDCx5p33_ASAP7_75t_R g7794 ( 
.A(n_6757),
.Y(n_7794)
);

CKINVDCx5p33_ASAP7_75t_R g7795 ( 
.A(n_6764),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_6912),
.Y(n_7796)
);

CKINVDCx5p33_ASAP7_75t_R g7797 ( 
.A(n_6770),
.Y(n_7797)
);

CKINVDCx11_ASAP7_75t_R g7798 ( 
.A(n_6103),
.Y(n_7798)
);

CKINVDCx5p33_ASAP7_75t_R g7799 ( 
.A(n_6780),
.Y(n_7799)
);

BUFx5_ASAP7_75t_L g7800 ( 
.A(n_6095),
.Y(n_7800)
);

INVx1_ASAP7_75t_L g7801 ( 
.A(n_6912),
.Y(n_7801)
);

CKINVDCx5p33_ASAP7_75t_R g7802 ( 
.A(n_6796),
.Y(n_7802)
);

INVx1_ASAP7_75t_L g7803 ( 
.A(n_7062),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7062),
.Y(n_7804)
);

INVx1_ASAP7_75t_L g7805 ( 
.A(n_7062),
.Y(n_7805)
);

CKINVDCx5p33_ASAP7_75t_R g7806 ( 
.A(n_6802),
.Y(n_7806)
);

INVx1_ASAP7_75t_L g7807 ( 
.A(n_7215),
.Y(n_7807)
);

CKINVDCx5p33_ASAP7_75t_R g7808 ( 
.A(n_6805),
.Y(n_7808)
);

CKINVDCx5p33_ASAP7_75t_R g7809 ( 
.A(n_6812),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7215),
.Y(n_7810)
);

CKINVDCx5p33_ASAP7_75t_R g7811 ( 
.A(n_6833),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_7215),
.Y(n_7812)
);

BUFx6f_ASAP7_75t_L g7813 ( 
.A(n_6373),
.Y(n_7813)
);

INVx2_ASAP7_75t_SL g7814 ( 
.A(n_6103),
.Y(n_7814)
);

CKINVDCx5p33_ASAP7_75t_R g7815 ( 
.A(n_6836),
.Y(n_7815)
);

BUFx10_ASAP7_75t_L g7816 ( 
.A(n_6322),
.Y(n_7816)
);

CKINVDCx5p33_ASAP7_75t_R g7817 ( 
.A(n_6852),
.Y(n_7817)
);

BUFx8_ASAP7_75t_SL g7818 ( 
.A(n_7288),
.Y(n_7818)
);

CKINVDCx5p33_ASAP7_75t_R g7819 ( 
.A(n_6858),
.Y(n_7819)
);

NOR2xp67_ASAP7_75t_L g7820 ( 
.A(n_7019),
.B(n_7),
.Y(n_7820)
);

INVx1_ASAP7_75t_SL g7821 ( 
.A(n_7371),
.Y(n_7821)
);

CKINVDCx5p33_ASAP7_75t_R g7822 ( 
.A(n_6860),
.Y(n_7822)
);

INVx1_ASAP7_75t_L g7823 ( 
.A(n_7253),
.Y(n_7823)
);

INVx1_ASAP7_75t_SL g7824 ( 
.A(n_7455),
.Y(n_7824)
);

CKINVDCx5p33_ASAP7_75t_R g7825 ( 
.A(n_6877),
.Y(n_7825)
);

CKINVDCx5p33_ASAP7_75t_R g7826 ( 
.A(n_6880),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7253),
.Y(n_7827)
);

INVx1_ASAP7_75t_L g7828 ( 
.A(n_7253),
.Y(n_7828)
);

CKINVDCx5p33_ASAP7_75t_R g7829 ( 
.A(n_6893),
.Y(n_7829)
);

CKINVDCx5p33_ASAP7_75t_R g7830 ( 
.A(n_6897),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_7256),
.Y(n_7831)
);

CKINVDCx5p33_ASAP7_75t_R g7832 ( 
.A(n_6900),
.Y(n_7832)
);

CKINVDCx5p33_ASAP7_75t_R g7833 ( 
.A(n_6920),
.Y(n_7833)
);

INVx1_ASAP7_75t_L g7834 ( 
.A(n_7256),
.Y(n_7834)
);

CKINVDCx5p33_ASAP7_75t_R g7835 ( 
.A(n_6921),
.Y(n_7835)
);

CKINVDCx5p33_ASAP7_75t_R g7836 ( 
.A(n_6923),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7256),
.Y(n_7837)
);

INVx1_ASAP7_75t_L g7838 ( 
.A(n_7391),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7391),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7391),
.Y(n_7840)
);

CKINVDCx5p33_ASAP7_75t_R g7841 ( 
.A(n_6925),
.Y(n_7841)
);

CKINVDCx20_ASAP7_75t_R g7842 ( 
.A(n_7205),
.Y(n_7842)
);

CKINVDCx20_ASAP7_75t_R g7843 ( 
.A(n_7344),
.Y(n_7843)
);

CKINVDCx5p33_ASAP7_75t_R g7844 ( 
.A(n_6931),
.Y(n_7844)
);

CKINVDCx5p33_ASAP7_75t_R g7845 ( 
.A(n_6941),
.Y(n_7845)
);

INVx2_ASAP7_75t_SL g7846 ( 
.A(n_6211),
.Y(n_7846)
);

CKINVDCx5p33_ASAP7_75t_R g7847 ( 
.A(n_6943),
.Y(n_7847)
);

INVx1_ASAP7_75t_SL g7848 ( 
.A(n_7486),
.Y(n_7848)
);

CKINVDCx20_ASAP7_75t_R g7849 ( 
.A(n_7378),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_7521),
.Y(n_7850)
);

INVx2_ASAP7_75t_L g7851 ( 
.A(n_7521),
.Y(n_7851)
);

BUFx2_ASAP7_75t_L g7852 ( 
.A(n_7544),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_7521),
.Y(n_7853)
);

BUFx3_ASAP7_75t_L g7854 ( 
.A(n_6517),
.Y(n_7854)
);

CKINVDCx5p33_ASAP7_75t_R g7855 ( 
.A(n_6950),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_6246),
.Y(n_7856)
);

BUFx2_ASAP7_75t_L g7857 ( 
.A(n_7541),
.Y(n_7857)
);

CKINVDCx5p33_ASAP7_75t_R g7858 ( 
.A(n_6966),
.Y(n_7858)
);

CKINVDCx5p33_ASAP7_75t_R g7859 ( 
.A(n_6979),
.Y(n_7859)
);

INVx3_ASAP7_75t_L g7860 ( 
.A(n_6347),
.Y(n_7860)
);

CKINVDCx5p33_ASAP7_75t_R g7861 ( 
.A(n_6995),
.Y(n_7861)
);

INVxp67_ASAP7_75t_L g7862 ( 
.A(n_6400),
.Y(n_7862)
);

HB1xp67_ASAP7_75t_L g7863 ( 
.A(n_6788),
.Y(n_7863)
);

CKINVDCx5p33_ASAP7_75t_R g7864 ( 
.A(n_6998),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_6382),
.Y(n_7865)
);

INVx1_ASAP7_75t_L g7866 ( 
.A(n_6383),
.Y(n_7866)
);

CKINVDCx5p33_ASAP7_75t_R g7867 ( 
.A(n_7011),
.Y(n_7867)
);

CKINVDCx5p33_ASAP7_75t_R g7868 ( 
.A(n_7016),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_6470),
.Y(n_7869)
);

HB1xp67_ASAP7_75t_L g7870 ( 
.A(n_6795),
.Y(n_7870)
);

INVxp67_ASAP7_75t_L g7871 ( 
.A(n_6424),
.Y(n_7871)
);

INVx1_ASAP7_75t_L g7872 ( 
.A(n_6568),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_6573),
.Y(n_7873)
);

INVx1_ASAP7_75t_SL g7874 ( 
.A(n_6089),
.Y(n_7874)
);

CKINVDCx5p33_ASAP7_75t_R g7875 ( 
.A(n_7032),
.Y(n_7875)
);

CKINVDCx16_ASAP7_75t_R g7876 ( 
.A(n_6809),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_6596),
.Y(n_7877)
);

CKINVDCx5p33_ASAP7_75t_R g7878 ( 
.A(n_7038),
.Y(n_7878)
);

CKINVDCx5p33_ASAP7_75t_R g7879 ( 
.A(n_7041),
.Y(n_7879)
);

CKINVDCx5p33_ASAP7_75t_R g7880 ( 
.A(n_7042),
.Y(n_7880)
);

CKINVDCx5p33_ASAP7_75t_R g7881 ( 
.A(n_7053),
.Y(n_7881)
);

INVx1_ASAP7_75t_L g7882 ( 
.A(n_6791),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_6838),
.Y(n_7883)
);

NOR2xp67_ASAP7_75t_L g7884 ( 
.A(n_7366),
.B(n_7),
.Y(n_7884)
);

BUFx6f_ASAP7_75t_L g7885 ( 
.A(n_6373),
.Y(n_7885)
);

CKINVDCx5p33_ASAP7_75t_R g7886 ( 
.A(n_7054),
.Y(n_7886)
);

INVxp67_ASAP7_75t_L g7887 ( 
.A(n_6707),
.Y(n_7887)
);

CKINVDCx5p33_ASAP7_75t_R g7888 ( 
.A(n_7073),
.Y(n_7888)
);

CKINVDCx5p33_ASAP7_75t_R g7889 ( 
.A(n_7106),
.Y(n_7889)
);

CKINVDCx5p33_ASAP7_75t_R g7890 ( 
.A(n_7109),
.Y(n_7890)
);

CKINVDCx5p33_ASAP7_75t_R g7891 ( 
.A(n_7112),
.Y(n_7891)
);

INVx1_ASAP7_75t_L g7892 ( 
.A(n_6874),
.Y(n_7892)
);

INVx2_ASAP7_75t_L g7893 ( 
.A(n_6185),
.Y(n_7893)
);

INVx1_ASAP7_75t_L g7894 ( 
.A(n_6949),
.Y(n_7894)
);

INVx3_ASAP7_75t_L g7895 ( 
.A(n_6959),
.Y(n_7895)
);

CKINVDCx5p33_ASAP7_75t_R g7896 ( 
.A(n_7117),
.Y(n_7896)
);

INVx1_ASAP7_75t_L g7897 ( 
.A(n_6975),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_7021),
.Y(n_7898)
);

CKINVDCx5p33_ASAP7_75t_R g7899 ( 
.A(n_7120),
.Y(n_7899)
);

CKINVDCx5p33_ASAP7_75t_R g7900 ( 
.A(n_7130),
.Y(n_7900)
);

CKINVDCx5p33_ASAP7_75t_R g7901 ( 
.A(n_7150),
.Y(n_7901)
);

BUFx3_ASAP7_75t_L g7902 ( 
.A(n_6963),
.Y(n_7902)
);

INVx1_ASAP7_75t_L g7903 ( 
.A(n_7357),
.Y(n_7903)
);

CKINVDCx5p33_ASAP7_75t_R g7904 ( 
.A(n_7153),
.Y(n_7904)
);

INVx1_ASAP7_75t_L g7905 ( 
.A(n_7469),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7476),
.Y(n_7906)
);

CKINVDCx5p33_ASAP7_75t_R g7907 ( 
.A(n_7192),
.Y(n_7907)
);

CKINVDCx5p33_ASAP7_75t_R g7908 ( 
.A(n_7199),
.Y(n_7908)
);

NOR2xp67_ASAP7_75t_L g7909 ( 
.A(n_7233),
.B(n_8),
.Y(n_7909)
);

CKINVDCx5p33_ASAP7_75t_R g7910 ( 
.A(n_7207),
.Y(n_7910)
);

CKINVDCx5p33_ASAP7_75t_R g7911 ( 
.A(n_7218),
.Y(n_7911)
);

CKINVDCx5p33_ASAP7_75t_R g7912 ( 
.A(n_7221),
.Y(n_7912)
);

CKINVDCx16_ASAP7_75t_R g7913 ( 
.A(n_6821),
.Y(n_7913)
);

INVxp33_ASAP7_75t_L g7914 ( 
.A(n_7287),
.Y(n_7914)
);

INVx1_ASAP7_75t_L g7915 ( 
.A(n_7490),
.Y(n_7915)
);

CKINVDCx5p33_ASAP7_75t_R g7916 ( 
.A(n_7231),
.Y(n_7916)
);

INVx1_ASAP7_75t_L g7917 ( 
.A(n_7513),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7540),
.Y(n_7918)
);

INVx1_ASAP7_75t_L g7919 ( 
.A(n_7545),
.Y(n_7919)
);

INVx1_ASAP7_75t_L g7920 ( 
.A(n_6088),
.Y(n_7920)
);

CKINVDCx5p33_ASAP7_75t_R g7921 ( 
.A(n_7290),
.Y(n_7921)
);

CKINVDCx5p33_ASAP7_75t_R g7922 ( 
.A(n_7292),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_7524),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7526),
.Y(n_7924)
);

INVx1_ASAP7_75t_L g7925 ( 
.A(n_7528),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_7536),
.Y(n_7926)
);

CKINVDCx5p33_ASAP7_75t_R g7927 ( 
.A(n_7294),
.Y(n_7927)
);

BUFx2_ASAP7_75t_L g7928 ( 
.A(n_6853),
.Y(n_7928)
);

CKINVDCx5p33_ASAP7_75t_R g7929 ( 
.A(n_7320),
.Y(n_7929)
);

INVx1_ASAP7_75t_L g7930 ( 
.A(n_7537),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_7538),
.Y(n_7931)
);

INVx2_ASAP7_75t_SL g7932 ( 
.A(n_6211),
.Y(n_7932)
);

INVx1_ASAP7_75t_L g7933 ( 
.A(n_6092),
.Y(n_7933)
);

INVx2_ASAP7_75t_L g7934 ( 
.A(n_6185),
.Y(n_7934)
);

NOR2xp33_ASAP7_75t_L g7935 ( 
.A(n_7280),
.B(n_8),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_6094),
.Y(n_7936)
);

CKINVDCx5p33_ASAP7_75t_R g7937 ( 
.A(n_7330),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_6104),
.Y(n_7938)
);

INVx1_ASAP7_75t_L g7939 ( 
.A(n_6112),
.Y(n_7939)
);

CKINVDCx5p33_ASAP7_75t_R g7940 ( 
.A(n_7331),
.Y(n_7940)
);

INVx1_ASAP7_75t_L g7941 ( 
.A(n_6124),
.Y(n_7941)
);

HB1xp67_ASAP7_75t_L g7942 ( 
.A(n_7520),
.Y(n_7942)
);

CKINVDCx5p33_ASAP7_75t_R g7943 ( 
.A(n_7332),
.Y(n_7943)
);

INVx1_ASAP7_75t_SL g7944 ( 
.A(n_6287),
.Y(n_7944)
);

CKINVDCx5p33_ASAP7_75t_R g7945 ( 
.A(n_7345),
.Y(n_7945)
);

INVx1_ASAP7_75t_L g7946 ( 
.A(n_6125),
.Y(n_7946)
);

INVx1_ASAP7_75t_SL g7947 ( 
.A(n_6228),
.Y(n_7947)
);

CKINVDCx5p33_ASAP7_75t_R g7948 ( 
.A(n_7350),
.Y(n_7948)
);

CKINVDCx5p33_ASAP7_75t_R g7949 ( 
.A(n_7382),
.Y(n_7949)
);

INVx1_ASAP7_75t_L g7950 ( 
.A(n_6129),
.Y(n_7950)
);

CKINVDCx5p33_ASAP7_75t_R g7951 ( 
.A(n_7384),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_6133),
.Y(n_7952)
);

INVx1_ASAP7_75t_L g7953 ( 
.A(n_6134),
.Y(n_7953)
);

CKINVDCx5p33_ASAP7_75t_R g7954 ( 
.A(n_7386),
.Y(n_7954)
);

CKINVDCx20_ASAP7_75t_R g7955 ( 
.A(n_7416),
.Y(n_7955)
);

INVx2_ASAP7_75t_L g7956 ( 
.A(n_6185),
.Y(n_7956)
);

INVx1_ASAP7_75t_L g7957 ( 
.A(n_7516),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7517),
.Y(n_7958)
);

INVx1_ASAP7_75t_L g7959 ( 
.A(n_6139),
.Y(n_7959)
);

OR2x2_ASAP7_75t_L g7960 ( 
.A(n_6172),
.B(n_10),
.Y(n_7960)
);

INVx1_ASAP7_75t_L g7961 ( 
.A(n_6142),
.Y(n_7961)
);

INVx1_ASAP7_75t_L g7962 ( 
.A(n_6143),
.Y(n_7962)
);

CKINVDCx5p33_ASAP7_75t_R g7963 ( 
.A(n_7388),
.Y(n_7963)
);

CKINVDCx5p33_ASAP7_75t_R g7964 ( 
.A(n_7400),
.Y(n_7964)
);

CKINVDCx5p33_ASAP7_75t_R g7965 ( 
.A(n_7403),
.Y(n_7965)
);

CKINVDCx5p33_ASAP7_75t_R g7966 ( 
.A(n_7425),
.Y(n_7966)
);

CKINVDCx5p33_ASAP7_75t_R g7967 ( 
.A(n_7437),
.Y(n_7967)
);

INVx1_ASAP7_75t_L g7968 ( 
.A(n_6162),
.Y(n_7968)
);

INVx2_ASAP7_75t_L g7969 ( 
.A(n_6185),
.Y(n_7969)
);

CKINVDCx5p33_ASAP7_75t_R g7970 ( 
.A(n_7462),
.Y(n_7970)
);

CKINVDCx5p33_ASAP7_75t_R g7971 ( 
.A(n_7473),
.Y(n_7971)
);

BUFx3_ASAP7_75t_L g7972 ( 
.A(n_6963),
.Y(n_7972)
);

CKINVDCx5p33_ASAP7_75t_R g7973 ( 
.A(n_7478),
.Y(n_7973)
);

CKINVDCx5p33_ASAP7_75t_R g7974 ( 
.A(n_7493),
.Y(n_7974)
);

BUFx2_ASAP7_75t_L g7975 ( 
.A(n_6957),
.Y(n_7975)
);

INVx2_ASAP7_75t_L g7976 ( 
.A(n_6185),
.Y(n_7976)
);

INVx1_ASAP7_75t_L g7977 ( 
.A(n_6180),
.Y(n_7977)
);

CKINVDCx5p33_ASAP7_75t_R g7978 ( 
.A(n_7499),
.Y(n_7978)
);

CKINVDCx5p33_ASAP7_75t_R g7979 ( 
.A(n_7506),
.Y(n_7979)
);

CKINVDCx16_ASAP7_75t_R g7980 ( 
.A(n_7064),
.Y(n_7980)
);

CKINVDCx5p33_ASAP7_75t_R g7981 ( 
.A(n_7507),
.Y(n_7981)
);

CKINVDCx5p33_ASAP7_75t_R g7982 ( 
.A(n_7531),
.Y(n_7982)
);

CKINVDCx5p33_ASAP7_75t_R g7983 ( 
.A(n_7456),
.Y(n_7983)
);

CKINVDCx5p33_ASAP7_75t_R g7984 ( 
.A(n_7479),
.Y(n_7984)
);

CKINVDCx20_ASAP7_75t_R g7985 ( 
.A(n_6264),
.Y(n_7985)
);

CKINVDCx5p33_ASAP7_75t_R g7986 ( 
.A(n_7076),
.Y(n_7986)
);

INVx1_ASAP7_75t_L g7987 ( 
.A(n_6186),
.Y(n_7987)
);

BUFx3_ASAP7_75t_L g7988 ( 
.A(n_7198),
.Y(n_7988)
);

INVx1_ASAP7_75t_L g7989 ( 
.A(n_6190),
.Y(n_7989)
);

INVx2_ASAP7_75t_L g7990 ( 
.A(n_7022),
.Y(n_7990)
);

CKINVDCx5p33_ASAP7_75t_R g7991 ( 
.A(n_7100),
.Y(n_7991)
);

CKINVDCx5p33_ASAP7_75t_R g7992 ( 
.A(n_7149),
.Y(n_7992)
);

CKINVDCx5p33_ASAP7_75t_R g7993 ( 
.A(n_7151),
.Y(n_7993)
);

INVx1_ASAP7_75t_L g7994 ( 
.A(n_6192),
.Y(n_7994)
);

BUFx10_ASAP7_75t_L g7995 ( 
.A(n_6078),
.Y(n_7995)
);

NOR2xp67_ASAP7_75t_L g7996 ( 
.A(n_6452),
.B(n_11),
.Y(n_7996)
);

CKINVDCx5p33_ASAP7_75t_R g7997 ( 
.A(n_7164),
.Y(n_7997)
);

INVx1_ASAP7_75t_L g7998 ( 
.A(n_6199),
.Y(n_7998)
);

BUFx3_ASAP7_75t_L g7999 ( 
.A(n_7198),
.Y(n_7999)
);

INVx1_ASAP7_75t_SL g8000 ( 
.A(n_6189),
.Y(n_8000)
);

CKINVDCx20_ASAP7_75t_R g8001 ( 
.A(n_7046),
.Y(n_8001)
);

INVx2_ASAP7_75t_L g8002 ( 
.A(n_7022),
.Y(n_8002)
);

CKINVDCx16_ASAP7_75t_R g8003 ( 
.A(n_7317),
.Y(n_8003)
);

INVx2_ASAP7_75t_L g8004 ( 
.A(n_7022),
.Y(n_8004)
);

CKINVDCx20_ASAP7_75t_R g8005 ( 
.A(n_7235),
.Y(n_8005)
);

CKINVDCx20_ASAP7_75t_R g8006 ( 
.A(n_7361),
.Y(n_8006)
);

BUFx6f_ASAP7_75t_L g8007 ( 
.A(n_6373),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_6212),
.Y(n_8008)
);

INVx1_ASAP7_75t_L g8009 ( 
.A(n_6239),
.Y(n_8009)
);

CKINVDCx5p33_ASAP7_75t_R g8010 ( 
.A(n_7430),
.Y(n_8010)
);

INVx1_ASAP7_75t_L g8011 ( 
.A(n_6242),
.Y(n_8011)
);

BUFx6f_ASAP7_75t_L g8012 ( 
.A(n_6655),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_6253),
.Y(n_8013)
);

INVx1_ASAP7_75t_L g8014 ( 
.A(n_6258),
.Y(n_8014)
);

CKINVDCx5p33_ASAP7_75t_R g8015 ( 
.A(n_6746),
.Y(n_8015)
);

INVx1_ASAP7_75t_L g8016 ( 
.A(n_7767),
.Y(n_8016)
);

CKINVDCx5p33_ASAP7_75t_R g8017 ( 
.A(n_7562),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7851),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7669),
.Y(n_8019)
);

INVx1_ASAP7_75t_L g8020 ( 
.A(n_7672),
.Y(n_8020)
);

CKINVDCx5p33_ASAP7_75t_R g8021 ( 
.A(n_7563),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7675),
.Y(n_8022)
);

INVx1_ASAP7_75t_L g8023 ( 
.A(n_7678),
.Y(n_8023)
);

INVx1_ASAP7_75t_L g8024 ( 
.A(n_7679),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7681),
.Y(n_8025)
);

INVx1_ASAP7_75t_L g8026 ( 
.A(n_7682),
.Y(n_8026)
);

HB1xp67_ASAP7_75t_L g8027 ( 
.A(n_7986),
.Y(n_8027)
);

INVx1_ASAP7_75t_L g8028 ( 
.A(n_7684),
.Y(n_8028)
);

INVx1_ASAP7_75t_L g8029 ( 
.A(n_7686),
.Y(n_8029)
);

INVx1_ASAP7_75t_L g8030 ( 
.A(n_7687),
.Y(n_8030)
);

BUFx2_ASAP7_75t_L g8031 ( 
.A(n_7991),
.Y(n_8031)
);

BUFx5_ASAP7_75t_L g8032 ( 
.A(n_7556),
.Y(n_8032)
);

INVx1_ASAP7_75t_L g8033 ( 
.A(n_7689),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_7690),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_7692),
.Y(n_8035)
);

INVxp67_ASAP7_75t_L g8036 ( 
.A(n_7560),
.Y(n_8036)
);

INVx1_ASAP7_75t_L g8037 ( 
.A(n_7696),
.Y(n_8037)
);

INVxp67_ASAP7_75t_SL g8038 ( 
.A(n_7553),
.Y(n_8038)
);

INVx1_ASAP7_75t_L g8039 ( 
.A(n_7697),
.Y(n_8039)
);

INVxp33_ASAP7_75t_SL g8040 ( 
.A(n_7559),
.Y(n_8040)
);

INVx1_ASAP7_75t_L g8041 ( 
.A(n_7699),
.Y(n_8041)
);

INVx1_ASAP7_75t_L g8042 ( 
.A(n_7701),
.Y(n_8042)
);

INVxp33_ASAP7_75t_SL g8043 ( 
.A(n_7549),
.Y(n_8043)
);

INVx3_ASAP7_75t_L g8044 ( 
.A(n_7553),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_7702),
.Y(n_8045)
);

INVx1_ASAP7_75t_L g8046 ( 
.A(n_7703),
.Y(n_8046)
);

BUFx2_ASAP7_75t_L g8047 ( 
.A(n_7992),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7705),
.Y(n_8048)
);

CKINVDCx5p33_ASAP7_75t_R g8049 ( 
.A(n_7564),
.Y(n_8049)
);

INVx1_ASAP7_75t_L g8050 ( 
.A(n_7707),
.Y(n_8050)
);

INVx1_ASAP7_75t_L g8051 ( 
.A(n_7708),
.Y(n_8051)
);

INVx1_ASAP7_75t_L g8052 ( 
.A(n_7719),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_7723),
.Y(n_8053)
);

INVx1_ASAP7_75t_L g8054 ( 
.A(n_7725),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_7736),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_7741),
.Y(n_8056)
);

INVx1_ASAP7_75t_L g8057 ( 
.A(n_7742),
.Y(n_8057)
);

INVx1_ASAP7_75t_L g8058 ( 
.A(n_7744),
.Y(n_8058)
);

CKINVDCx5p33_ASAP7_75t_R g8059 ( 
.A(n_7570),
.Y(n_8059)
);

INVx1_ASAP7_75t_L g8060 ( 
.A(n_7747),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_7749),
.Y(n_8061)
);

INVx1_ASAP7_75t_L g8062 ( 
.A(n_7750),
.Y(n_8062)
);

CKINVDCx20_ASAP7_75t_R g8063 ( 
.A(n_7547),
.Y(n_8063)
);

INVxp67_ASAP7_75t_SL g8064 ( 
.A(n_7553),
.Y(n_8064)
);

INVx1_ASAP7_75t_L g8065 ( 
.A(n_7751),
.Y(n_8065)
);

CKINVDCx5p33_ASAP7_75t_R g8066 ( 
.A(n_7572),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7754),
.Y(n_8067)
);

CKINVDCx20_ASAP7_75t_R g8068 ( 
.A(n_7550),
.Y(n_8068)
);

CKINVDCx5p33_ASAP7_75t_R g8069 ( 
.A(n_7574),
.Y(n_8069)
);

INVx1_ASAP7_75t_L g8070 ( 
.A(n_7757),
.Y(n_8070)
);

INVxp67_ASAP7_75t_SL g8071 ( 
.A(n_7618),
.Y(n_8071)
);

INVxp33_ASAP7_75t_SL g8072 ( 
.A(n_7551),
.Y(n_8072)
);

INVxp67_ASAP7_75t_SL g8073 ( 
.A(n_7618),
.Y(n_8073)
);

INVx1_ASAP7_75t_L g8074 ( 
.A(n_7758),
.Y(n_8074)
);

CKINVDCx16_ASAP7_75t_R g8075 ( 
.A(n_7591),
.Y(n_8075)
);

INVx1_ASAP7_75t_L g8076 ( 
.A(n_7760),
.Y(n_8076)
);

INVx1_ASAP7_75t_L g8077 ( 
.A(n_7764),
.Y(n_8077)
);

BUFx3_ASAP7_75t_L g8078 ( 
.A(n_7860),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7766),
.Y(n_8079)
);

INVxp33_ASAP7_75t_SL g8080 ( 
.A(n_7552),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_7776),
.Y(n_8081)
);

CKINVDCx5p33_ASAP7_75t_R g8082 ( 
.A(n_7580),
.Y(n_8082)
);

INVx1_ASAP7_75t_L g8083 ( 
.A(n_7782),
.Y(n_8083)
);

BUFx3_ASAP7_75t_L g8084 ( 
.A(n_7860),
.Y(n_8084)
);

CKINVDCx5p33_ASAP7_75t_R g8085 ( 
.A(n_7583),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_7787),
.Y(n_8086)
);

CKINVDCx5p33_ASAP7_75t_R g8087 ( 
.A(n_7584),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_7796),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_7801),
.Y(n_8089)
);

CKINVDCx20_ASAP7_75t_R g8090 ( 
.A(n_7565),
.Y(n_8090)
);

INVx1_ASAP7_75t_L g8091 ( 
.A(n_7803),
.Y(n_8091)
);

INVxp67_ASAP7_75t_SL g8092 ( 
.A(n_7618),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_7804),
.Y(n_8093)
);

CKINVDCx20_ASAP7_75t_R g8094 ( 
.A(n_7575),
.Y(n_8094)
);

CKINVDCx5p33_ASAP7_75t_R g8095 ( 
.A(n_7586),
.Y(n_8095)
);

INVx1_ASAP7_75t_L g8096 ( 
.A(n_7805),
.Y(n_8096)
);

INVxp33_ASAP7_75t_SL g8097 ( 
.A(n_7555),
.Y(n_8097)
);

INVx3_ASAP7_75t_L g8098 ( 
.A(n_7639),
.Y(n_8098)
);

INVx1_ASAP7_75t_L g8099 ( 
.A(n_7807),
.Y(n_8099)
);

INVx2_ASAP7_75t_L g8100 ( 
.A(n_7639),
.Y(n_8100)
);

INVxp67_ASAP7_75t_L g8101 ( 
.A(n_7691),
.Y(n_8101)
);

INVxp67_ASAP7_75t_SL g8102 ( 
.A(n_7639),
.Y(n_8102)
);

INVx1_ASAP7_75t_L g8103 ( 
.A(n_7810),
.Y(n_8103)
);

CKINVDCx5p33_ASAP7_75t_R g8104 ( 
.A(n_7588),
.Y(n_8104)
);

INVx1_ASAP7_75t_L g8105 ( 
.A(n_7812),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_7823),
.Y(n_8106)
);

INVx1_ASAP7_75t_L g8107 ( 
.A(n_7827),
.Y(n_8107)
);

INVx1_ASAP7_75t_L g8108 ( 
.A(n_7828),
.Y(n_8108)
);

INVx1_ASAP7_75t_L g8109 ( 
.A(n_7831),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_7834),
.Y(n_8110)
);

INVxp67_ASAP7_75t_L g8111 ( 
.A(n_7784),
.Y(n_8111)
);

INVx1_ASAP7_75t_L g8112 ( 
.A(n_7837),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7838),
.Y(n_8113)
);

CKINVDCx5p33_ASAP7_75t_R g8114 ( 
.A(n_7589),
.Y(n_8114)
);

CKINVDCx5p33_ASAP7_75t_R g8115 ( 
.A(n_7593),
.Y(n_8115)
);

CKINVDCx20_ASAP7_75t_R g8116 ( 
.A(n_7606),
.Y(n_8116)
);

INVx1_ASAP7_75t_L g8117 ( 
.A(n_7839),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_7840),
.Y(n_8118)
);

INVxp67_ASAP7_75t_L g8119 ( 
.A(n_7863),
.Y(n_8119)
);

INVx1_ASAP7_75t_L g8120 ( 
.A(n_7850),
.Y(n_8120)
);

INVx1_ASAP7_75t_L g8121 ( 
.A(n_7853),
.Y(n_8121)
);

INVx1_ASAP7_75t_L g8122 ( 
.A(n_7746),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_7746),
.Y(n_8123)
);

INVx1_ASAP7_75t_L g8124 ( 
.A(n_7746),
.Y(n_8124)
);

INVx1_ASAP7_75t_L g8125 ( 
.A(n_7762),
.Y(n_8125)
);

INVxp67_ASAP7_75t_SL g8126 ( 
.A(n_7762),
.Y(n_8126)
);

INVxp67_ASAP7_75t_SL g8127 ( 
.A(n_7762),
.Y(n_8127)
);

BUFx3_ASAP7_75t_L g8128 ( 
.A(n_7895),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_7785),
.Y(n_8129)
);

HB1xp67_ASAP7_75t_L g8130 ( 
.A(n_7993),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_7785),
.Y(n_8131)
);

INVx1_ASAP7_75t_L g8132 ( 
.A(n_7785),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_7813),
.Y(n_8133)
);

CKINVDCx14_ASAP7_75t_R g8134 ( 
.A(n_7592),
.Y(n_8134)
);

INVxp33_ASAP7_75t_SL g8135 ( 
.A(n_7557),
.Y(n_8135)
);

INVx1_ASAP7_75t_L g8136 ( 
.A(n_7813),
.Y(n_8136)
);

INVx1_ASAP7_75t_L g8137 ( 
.A(n_7813),
.Y(n_8137)
);

CKINVDCx20_ASAP7_75t_R g8138 ( 
.A(n_7623),
.Y(n_8138)
);

CKINVDCx5p33_ASAP7_75t_R g8139 ( 
.A(n_7595),
.Y(n_8139)
);

INVx1_ASAP7_75t_L g8140 ( 
.A(n_7885),
.Y(n_8140)
);

INVx1_ASAP7_75t_L g8141 ( 
.A(n_7885),
.Y(n_8141)
);

INVxp67_ASAP7_75t_SL g8142 ( 
.A(n_7885),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_8007),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_8007),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_8007),
.Y(n_8145)
);

CKINVDCx5p33_ASAP7_75t_R g8146 ( 
.A(n_7598),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_8012),
.Y(n_8147)
);

CKINVDCx5p33_ASAP7_75t_R g8148 ( 
.A(n_7599),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_8012),
.Y(n_8149)
);

INVx1_ASAP7_75t_L g8150 ( 
.A(n_8012),
.Y(n_8150)
);

INVx1_ASAP7_75t_L g8151 ( 
.A(n_7558),
.Y(n_8151)
);

INVxp67_ASAP7_75t_SL g8152 ( 
.A(n_7895),
.Y(n_8152)
);

BUFx6f_ASAP7_75t_L g8153 ( 
.A(n_7561),
.Y(n_8153)
);

INVx1_ASAP7_75t_L g8154 ( 
.A(n_7566),
.Y(n_8154)
);

INVx1_ASAP7_75t_L g8155 ( 
.A(n_7567),
.Y(n_8155)
);

INVxp67_ASAP7_75t_SL g8156 ( 
.A(n_7935),
.Y(n_8156)
);

HB1xp67_ASAP7_75t_L g8157 ( 
.A(n_7997),
.Y(n_8157)
);

INVx2_ASAP7_75t_L g8158 ( 
.A(n_7568),
.Y(n_8158)
);

CKINVDCx5p33_ASAP7_75t_R g8159 ( 
.A(n_7601),
.Y(n_8159)
);

INVx1_ASAP7_75t_L g8160 ( 
.A(n_7569),
.Y(n_8160)
);

INVx2_ASAP7_75t_L g8161 ( 
.A(n_7576),
.Y(n_8161)
);

INVxp67_ASAP7_75t_SL g8162 ( 
.A(n_7909),
.Y(n_8162)
);

CKINVDCx20_ASAP7_75t_R g8163 ( 
.A(n_7624),
.Y(n_8163)
);

INVx2_ASAP7_75t_L g8164 ( 
.A(n_7596),
.Y(n_8164)
);

INVxp67_ASAP7_75t_SL g8165 ( 
.A(n_7856),
.Y(n_8165)
);

INVxp33_ASAP7_75t_SL g8166 ( 
.A(n_7983),
.Y(n_8166)
);

CKINVDCx5p33_ASAP7_75t_R g8167 ( 
.A(n_7607),
.Y(n_8167)
);

CKINVDCx5p33_ASAP7_75t_R g8168 ( 
.A(n_7612),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7573),
.Y(n_8169)
);

INVxp67_ASAP7_75t_SL g8170 ( 
.A(n_7865),
.Y(n_8170)
);

INVxp33_ASAP7_75t_L g8171 ( 
.A(n_7870),
.Y(n_8171)
);

INVx1_ASAP7_75t_L g8172 ( 
.A(n_7577),
.Y(n_8172)
);

INVxp67_ASAP7_75t_L g8173 ( 
.A(n_7942),
.Y(n_8173)
);

INVxp67_ASAP7_75t_SL g8174 ( 
.A(n_7866),
.Y(n_8174)
);

INVx1_ASAP7_75t_L g8175 ( 
.A(n_7578),
.Y(n_8175)
);

INVxp67_ASAP7_75t_SL g8176 ( 
.A(n_7869),
.Y(n_8176)
);

INVx1_ASAP7_75t_L g8177 ( 
.A(n_7579),
.Y(n_8177)
);

INVx1_ASAP7_75t_L g8178 ( 
.A(n_7581),
.Y(n_8178)
);

CKINVDCx5p33_ASAP7_75t_R g8179 ( 
.A(n_7615),
.Y(n_8179)
);

INVx1_ASAP7_75t_L g8180 ( 
.A(n_7585),
.Y(n_8180)
);

INVx1_ASAP7_75t_L g8181 ( 
.A(n_7587),
.Y(n_8181)
);

INVx1_ASAP7_75t_L g8182 ( 
.A(n_7590),
.Y(n_8182)
);

CKINVDCx20_ASAP7_75t_R g8183 ( 
.A(n_7628),
.Y(n_8183)
);

HB1xp67_ASAP7_75t_L g8184 ( 
.A(n_8010),
.Y(n_8184)
);

CKINVDCx5p33_ASAP7_75t_R g8185 ( 
.A(n_7620),
.Y(n_8185)
);

INVxp67_ASAP7_75t_SL g8186 ( 
.A(n_7872),
.Y(n_8186)
);

HB1xp67_ASAP7_75t_L g8187 ( 
.A(n_7928),
.Y(n_8187)
);

BUFx2_ASAP7_75t_L g8188 ( 
.A(n_7985),
.Y(n_8188)
);

CKINVDCx20_ASAP7_75t_R g8189 ( 
.A(n_7642),
.Y(n_8189)
);

INVxp33_ASAP7_75t_SL g8190 ( 
.A(n_7984),
.Y(n_8190)
);

CKINVDCx5p33_ASAP7_75t_R g8191 ( 
.A(n_7621),
.Y(n_8191)
);

CKINVDCx20_ASAP7_75t_R g8192 ( 
.A(n_7695),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7594),
.Y(n_8193)
);

INVx1_ASAP7_75t_L g8194 ( 
.A(n_7597),
.Y(n_8194)
);

CKINVDCx20_ASAP7_75t_R g8195 ( 
.A(n_7709),
.Y(n_8195)
);

INVxp67_ASAP7_75t_SL g8196 ( 
.A(n_7873),
.Y(n_8196)
);

INVx1_ASAP7_75t_L g8197 ( 
.A(n_7600),
.Y(n_8197)
);

INVx2_ASAP7_75t_L g8198 ( 
.A(n_7604),
.Y(n_8198)
);

INVx1_ASAP7_75t_SL g8199 ( 
.A(n_7874),
.Y(n_8199)
);

INVx1_ASAP7_75t_L g8200 ( 
.A(n_7602),
.Y(n_8200)
);

CKINVDCx5p33_ASAP7_75t_R g8201 ( 
.A(n_7630),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_7603),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_7608),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_7609),
.Y(n_8204)
);

INVx2_ASAP7_75t_L g8205 ( 
.A(n_7605),
.Y(n_8205)
);

INVx1_ASAP7_75t_SL g8206 ( 
.A(n_7944),
.Y(n_8206)
);

INVx2_ASAP7_75t_L g8207 ( 
.A(n_7614),
.Y(n_8207)
);

INVxp67_ASAP7_75t_SL g8208 ( 
.A(n_7877),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_7611),
.Y(n_8209)
);

INVx1_ASAP7_75t_L g8210 ( 
.A(n_7616),
.Y(n_8210)
);

INVxp67_ASAP7_75t_SL g8211 ( 
.A(n_7882),
.Y(n_8211)
);

CKINVDCx5p33_ASAP7_75t_R g8212 ( 
.A(n_7632),
.Y(n_8212)
);

INVx1_ASAP7_75t_L g8213 ( 
.A(n_7619),
.Y(n_8213)
);

BUFx2_ASAP7_75t_L g8214 ( 
.A(n_8001),
.Y(n_8214)
);

INVxp33_ASAP7_75t_SL g8215 ( 
.A(n_7548),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_7625),
.Y(n_8216)
);

INVx1_ASAP7_75t_L g8217 ( 
.A(n_7635),
.Y(n_8217)
);

INVx1_ASAP7_75t_L g8218 ( 
.A(n_7640),
.Y(n_8218)
);

CKINVDCx16_ASAP7_75t_R g8219 ( 
.A(n_7680),
.Y(n_8219)
);

INVx1_ASAP7_75t_L g8220 ( 
.A(n_7645),
.Y(n_8220)
);

CKINVDCx20_ASAP7_75t_R g8221 ( 
.A(n_7712),
.Y(n_8221)
);

INVxp33_ASAP7_75t_L g8222 ( 
.A(n_7914),
.Y(n_8222)
);

CKINVDCx5p33_ASAP7_75t_R g8223 ( 
.A(n_7633),
.Y(n_8223)
);

INVx1_ASAP7_75t_L g8224 ( 
.A(n_7646),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_7649),
.Y(n_8225)
);

INVxp67_ASAP7_75t_SL g8226 ( 
.A(n_7883),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7650),
.Y(n_8227)
);

INVx1_ASAP7_75t_L g8228 ( 
.A(n_7654),
.Y(n_8228)
);

INVx1_ASAP7_75t_L g8229 ( 
.A(n_7658),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_7659),
.Y(n_8230)
);

CKINVDCx5p33_ASAP7_75t_R g8231 ( 
.A(n_7634),
.Y(n_8231)
);

INVx1_ASAP7_75t_L g8232 ( 
.A(n_7661),
.Y(n_8232)
);

CKINVDCx16_ASAP7_75t_R g8233 ( 
.A(n_7694),
.Y(n_8233)
);

INVxp67_ASAP7_75t_SL g8234 ( 
.A(n_7892),
.Y(n_8234)
);

INVxp33_ASAP7_75t_SL g8235 ( 
.A(n_7546),
.Y(n_8235)
);

INVx1_ASAP7_75t_L g8236 ( 
.A(n_7663),
.Y(n_8236)
);

BUFx3_ASAP7_75t_L g8237 ( 
.A(n_7857),
.Y(n_8237)
);

INVx1_ASAP7_75t_L g8238 ( 
.A(n_7918),
.Y(n_8238)
);

INVx1_ASAP7_75t_L g8239 ( 
.A(n_7919),
.Y(n_8239)
);

INVx1_ASAP7_75t_L g8240 ( 
.A(n_7920),
.Y(n_8240)
);

INVx1_ASAP7_75t_L g8241 ( 
.A(n_7923),
.Y(n_8241)
);

INVxp67_ASAP7_75t_SL g8242 ( 
.A(n_7894),
.Y(n_8242)
);

INVx1_ASAP7_75t_L g8243 ( 
.A(n_7924),
.Y(n_8243)
);

INVxp33_ASAP7_75t_L g8244 ( 
.A(n_7975),
.Y(n_8244)
);

CKINVDCx16_ASAP7_75t_R g8245 ( 
.A(n_7735),
.Y(n_8245)
);

CKINVDCx20_ASAP7_75t_R g8246 ( 
.A(n_7740),
.Y(n_8246)
);

INVx1_ASAP7_75t_L g8247 ( 
.A(n_7925),
.Y(n_8247)
);

INVxp67_ASAP7_75t_SL g8248 ( 
.A(n_7897),
.Y(n_8248)
);

BUFx3_ASAP7_75t_L g8249 ( 
.A(n_7898),
.Y(n_8249)
);

INVx1_ASAP7_75t_SL g8250 ( 
.A(n_7947),
.Y(n_8250)
);

INVxp67_ASAP7_75t_SL g8251 ( 
.A(n_7903),
.Y(n_8251)
);

INVx1_ASAP7_75t_L g8252 ( 
.A(n_7926),
.Y(n_8252)
);

INVx1_ASAP7_75t_L g8253 ( 
.A(n_7930),
.Y(n_8253)
);

INVx2_ASAP7_75t_L g8254 ( 
.A(n_7617),
.Y(n_8254)
);

CKINVDCx20_ASAP7_75t_R g8255 ( 
.A(n_7752),
.Y(n_8255)
);

CKINVDCx20_ASAP7_75t_R g8256 ( 
.A(n_7775),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7931),
.Y(n_8257)
);

CKINVDCx5p33_ASAP7_75t_R g8258 ( 
.A(n_7636),
.Y(n_8258)
);

INVxp67_ASAP7_75t_SL g8259 ( 
.A(n_7905),
.Y(n_8259)
);

CKINVDCx5p33_ASAP7_75t_R g8260 ( 
.A(n_7637),
.Y(n_8260)
);

CKINVDCx5p33_ASAP7_75t_R g8261 ( 
.A(n_7638),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_7933),
.Y(n_8262)
);

INVx1_ASAP7_75t_L g8263 ( 
.A(n_7936),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_7938),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_7939),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_7941),
.Y(n_8266)
);

INVx1_ASAP7_75t_L g8267 ( 
.A(n_7946),
.Y(n_8267)
);

CKINVDCx5p33_ASAP7_75t_R g8268 ( 
.A(n_7641),
.Y(n_8268)
);

INVxp67_ASAP7_75t_L g8269 ( 
.A(n_7629),
.Y(n_8269)
);

CKINVDCx16_ASAP7_75t_R g8270 ( 
.A(n_7772),
.Y(n_8270)
);

INVxp67_ASAP7_75t_SL g8271 ( 
.A(n_7906),
.Y(n_8271)
);

INVx2_ASAP7_75t_L g8272 ( 
.A(n_7622),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_7950),
.Y(n_8273)
);

INVx1_ASAP7_75t_L g8274 ( 
.A(n_7952),
.Y(n_8274)
);

INVx1_ASAP7_75t_L g8275 ( 
.A(n_7953),
.Y(n_8275)
);

INVx1_ASAP7_75t_L g8276 ( 
.A(n_7957),
.Y(n_8276)
);

INVx1_ASAP7_75t_L g8277 ( 
.A(n_7958),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_7959),
.Y(n_8278)
);

CKINVDCx5p33_ASAP7_75t_R g8279 ( 
.A(n_7643),
.Y(n_8279)
);

CKINVDCx5p33_ASAP7_75t_R g8280 ( 
.A(n_7644),
.Y(n_8280)
);

INVx1_ASAP7_75t_L g8281 ( 
.A(n_7961),
.Y(n_8281)
);

INVx1_ASAP7_75t_L g8282 ( 
.A(n_7962),
.Y(n_8282)
);

CKINVDCx5p33_ASAP7_75t_R g8283 ( 
.A(n_7647),
.Y(n_8283)
);

INVx1_ASAP7_75t_L g8284 ( 
.A(n_7968),
.Y(n_8284)
);

INVxp33_ASAP7_75t_L g8285 ( 
.A(n_7755),
.Y(n_8285)
);

BUFx3_ASAP7_75t_L g8286 ( 
.A(n_7915),
.Y(n_8286)
);

HB1xp67_ASAP7_75t_L g8287 ( 
.A(n_7773),
.Y(n_8287)
);

INVx1_ASAP7_75t_L g8288 ( 
.A(n_7977),
.Y(n_8288)
);

INVx1_ASAP7_75t_L g8289 ( 
.A(n_7987),
.Y(n_8289)
);

CKINVDCx5p33_ASAP7_75t_R g8290 ( 
.A(n_7648),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_7989),
.Y(n_8291)
);

INVx1_ASAP7_75t_L g8292 ( 
.A(n_7994),
.Y(n_8292)
);

INVx1_ASAP7_75t_L g8293 ( 
.A(n_7998),
.Y(n_8293)
);

INVx1_ASAP7_75t_L g8294 ( 
.A(n_8008),
.Y(n_8294)
);

CKINVDCx5p33_ASAP7_75t_R g8295 ( 
.A(n_7651),
.Y(n_8295)
);

INVxp67_ASAP7_75t_SL g8296 ( 
.A(n_7917),
.Y(n_8296)
);

CKINVDCx5p33_ASAP7_75t_R g8297 ( 
.A(n_7653),
.Y(n_8297)
);

NOR2xp33_ASAP7_75t_L g8298 ( 
.A(n_7655),
.B(n_7080),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_8009),
.Y(n_8299)
);

INVx2_ASAP7_75t_L g8300 ( 
.A(n_7662),
.Y(n_8300)
);

INVxp33_ASAP7_75t_SL g8301 ( 
.A(n_7656),
.Y(n_8301)
);

CKINVDCx5p33_ASAP7_75t_R g8302 ( 
.A(n_7657),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_8011),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_8013),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_8014),
.Y(n_8305)
);

CKINVDCx5p33_ASAP7_75t_R g8306 ( 
.A(n_7664),
.Y(n_8306)
);

INVxp67_ASAP7_75t_SL g8307 ( 
.A(n_7862),
.Y(n_8307)
);

INVxp33_ASAP7_75t_SL g8308 ( 
.A(n_7665),
.Y(n_8308)
);

CKINVDCx5p33_ASAP7_75t_R g8309 ( 
.A(n_7666),
.Y(n_8309)
);

CKINVDCx16_ASAP7_75t_R g8310 ( 
.A(n_7876),
.Y(n_8310)
);

CKINVDCx5p33_ASAP7_75t_R g8311 ( 
.A(n_7667),
.Y(n_8311)
);

INVx1_ASAP7_75t_L g8312 ( 
.A(n_7893),
.Y(n_8312)
);

INVxp67_ASAP7_75t_SL g8313 ( 
.A(n_7871),
.Y(n_8313)
);

HB1xp67_ASAP7_75t_L g8314 ( 
.A(n_7913),
.Y(n_8314)
);

INVx1_ASAP7_75t_L g8315 ( 
.A(n_7934),
.Y(n_8315)
);

INVx1_ASAP7_75t_L g8316 ( 
.A(n_7956),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_7969),
.Y(n_8317)
);

INVx1_ASAP7_75t_L g8318 ( 
.A(n_7976),
.Y(n_8318)
);

CKINVDCx5p33_ASAP7_75t_R g8319 ( 
.A(n_7670),
.Y(n_8319)
);

BUFx2_ASAP7_75t_L g8320 ( 
.A(n_8005),
.Y(n_8320)
);

CKINVDCx5p33_ASAP7_75t_R g8321 ( 
.A(n_7671),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_7990),
.Y(n_8322)
);

INVx2_ASAP7_75t_SL g8323 ( 
.A(n_7995),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_8002),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_8004),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7660),
.Y(n_8326)
);

INVx1_ASAP7_75t_L g8327 ( 
.A(n_7660),
.Y(n_8327)
);

INVx1_ASAP7_75t_L g8328 ( 
.A(n_7660),
.Y(n_8328)
);

BUFx6f_ASAP7_75t_L g8329 ( 
.A(n_7960),
.Y(n_8329)
);

INVx2_ASAP7_75t_L g8330 ( 
.A(n_7660),
.Y(n_8330)
);

CKINVDCx5p33_ASAP7_75t_R g8331 ( 
.A(n_7673),
.Y(n_8331)
);

INVxp67_ASAP7_75t_L g8332 ( 
.A(n_7693),
.Y(n_8332)
);

INVx1_ASAP7_75t_L g8333 ( 
.A(n_7660),
.Y(n_8333)
);

INVx1_ASAP7_75t_L g8334 ( 
.A(n_7800),
.Y(n_8334)
);

INVx2_ASAP7_75t_L g8335 ( 
.A(n_7800),
.Y(n_8335)
);

NOR2xp33_ASAP7_75t_L g8336 ( 
.A(n_7674),
.B(n_7098),
.Y(n_8336)
);

CKINVDCx20_ASAP7_75t_R g8337 ( 
.A(n_7842),
.Y(n_8337)
);

INVx1_ASAP7_75t_L g8338 ( 
.A(n_7800),
.Y(n_8338)
);

CKINVDCx5p33_ASAP7_75t_R g8339 ( 
.A(n_7676),
.Y(n_8339)
);

INVx1_ASAP7_75t_L g8340 ( 
.A(n_7800),
.Y(n_8340)
);

INVxp67_ASAP7_75t_SL g8341 ( 
.A(n_7887),
.Y(n_8341)
);

INVx1_ASAP7_75t_SL g8342 ( 
.A(n_8000),
.Y(n_8342)
);

INVx2_ASAP7_75t_L g8343 ( 
.A(n_7800),
.Y(n_8343)
);

INVxp67_ASAP7_75t_SL g8344 ( 
.A(n_7613),
.Y(n_8344)
);

HB1xp67_ASAP7_75t_L g8345 ( 
.A(n_7980),
.Y(n_8345)
);

CKINVDCx16_ASAP7_75t_R g8346 ( 
.A(n_8003),
.Y(n_8346)
);

INVx3_ASAP7_75t_L g8347 ( 
.A(n_7626),
.Y(n_8347)
);

INVxp67_ASAP7_75t_SL g8348 ( 
.A(n_7715),
.Y(n_8348)
);

INVx1_ASAP7_75t_L g8349 ( 
.A(n_7996),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_7554),
.Y(n_8350)
);

CKINVDCx5p33_ASAP7_75t_R g8351 ( 
.A(n_7677),
.Y(n_8351)
);

CKINVDCx5p33_ASAP7_75t_R g8352 ( 
.A(n_7685),
.Y(n_8352)
);

INVx1_ASAP7_75t_L g8353 ( 
.A(n_7571),
.Y(n_8353)
);

INVx1_ASAP7_75t_L g8354 ( 
.A(n_7582),
.Y(n_8354)
);

INVx1_ASAP7_75t_L g8355 ( 
.A(n_7631),
.Y(n_8355)
);

INVxp33_ASAP7_75t_SL g8356 ( 
.A(n_7688),
.Y(n_8356)
);

INVx1_ASAP7_75t_L g8357 ( 
.A(n_7652),
.Y(n_8357)
);

INVx1_ASAP7_75t_L g8358 ( 
.A(n_7700),
.Y(n_8358)
);

CKINVDCx5p33_ASAP7_75t_R g8359 ( 
.A(n_7698),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7729),
.Y(n_8360)
);

INVx1_ASAP7_75t_L g8361 ( 
.A(n_7730),
.Y(n_8361)
);

INVxp33_ASAP7_75t_L g8362 ( 
.A(n_7852),
.Y(n_8362)
);

HB1xp67_ASAP7_75t_L g8363 ( 
.A(n_7727),
.Y(n_8363)
);

INVx1_ASAP7_75t_L g8364 ( 
.A(n_7778),
.Y(n_8364)
);

INVxp33_ASAP7_75t_L g8365 ( 
.A(n_7788),
.Y(n_8365)
);

INVx1_ASAP7_75t_L g8366 ( 
.A(n_7820),
.Y(n_8366)
);

INVxp67_ASAP7_75t_SL g8367 ( 
.A(n_7627),
.Y(n_8367)
);

INVx1_ASAP7_75t_L g8368 ( 
.A(n_7884),
.Y(n_8368)
);

CKINVDCx5p33_ASAP7_75t_R g8369 ( 
.A(n_7704),
.Y(n_8369)
);

INVx1_ASAP7_75t_L g8370 ( 
.A(n_7854),
.Y(n_8370)
);

BUFx3_ASAP7_75t_L g8371 ( 
.A(n_7711),
.Y(n_8371)
);

BUFx2_ASAP7_75t_SL g8372 ( 
.A(n_8006),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7902),
.Y(n_8373)
);

CKINVDCx5p33_ASAP7_75t_R g8374 ( 
.A(n_7713),
.Y(n_8374)
);

INVxp33_ASAP7_75t_L g8375 ( 
.A(n_7818),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7972),
.Y(n_8376)
);

CKINVDCx5p33_ASAP7_75t_R g8377 ( 
.A(n_7714),
.Y(n_8377)
);

INVxp67_ASAP7_75t_SL g8378 ( 
.A(n_7706),
.Y(n_8378)
);

INVx1_ASAP7_75t_L g8379 ( 
.A(n_7988),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7999),
.Y(n_8380)
);

INVxp67_ASAP7_75t_L g8381 ( 
.A(n_7814),
.Y(n_8381)
);

CKINVDCx5p33_ASAP7_75t_R g8382 ( 
.A(n_7716),
.Y(n_8382)
);

INVx1_ASAP7_75t_L g8383 ( 
.A(n_7718),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_7720),
.Y(n_8384)
);

INVx1_ASAP7_75t_L g8385 ( 
.A(n_7721),
.Y(n_8385)
);

INVx1_ASAP7_75t_L g8386 ( 
.A(n_7722),
.Y(n_8386)
);

CKINVDCx16_ASAP7_75t_R g8387 ( 
.A(n_7610),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_7724),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7731),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7732),
.Y(n_8390)
);

CKINVDCx5p33_ASAP7_75t_R g8391 ( 
.A(n_7737),
.Y(n_8391)
);

HB1xp67_ASAP7_75t_L g8392 ( 
.A(n_7728),
.Y(n_8392)
);

CKINVDCx5p33_ASAP7_75t_R g8393 ( 
.A(n_7738),
.Y(n_8393)
);

INVx2_ASAP7_75t_L g8394 ( 
.A(n_7717),
.Y(n_8394)
);

INVxp33_ASAP7_75t_SL g8395 ( 
.A(n_7739),
.Y(n_8395)
);

INVx1_ASAP7_75t_L g8396 ( 
.A(n_7743),
.Y(n_8396)
);

CKINVDCx20_ASAP7_75t_R g8397 ( 
.A(n_7843),
.Y(n_8397)
);

INVx1_ASAP7_75t_L g8398 ( 
.A(n_7745),
.Y(n_8398)
);

CKINVDCx5p33_ASAP7_75t_R g8399 ( 
.A(n_7748),
.Y(n_8399)
);

INVx1_ASAP7_75t_L g8400 ( 
.A(n_7753),
.Y(n_8400)
);

CKINVDCx5p33_ASAP7_75t_R g8401 ( 
.A(n_7759),
.Y(n_8401)
);

INVx1_ASAP7_75t_L g8402 ( 
.A(n_7761),
.Y(n_8402)
);

CKINVDCx5p33_ASAP7_75t_R g8403 ( 
.A(n_7763),
.Y(n_8403)
);

INVx1_ASAP7_75t_SL g8404 ( 
.A(n_7849),
.Y(n_8404)
);

CKINVDCx20_ASAP7_75t_R g8405 ( 
.A(n_7955),
.Y(n_8405)
);

INVx1_ASAP7_75t_L g8406 ( 
.A(n_7765),
.Y(n_8406)
);

HB1xp67_ASAP7_75t_L g8407 ( 
.A(n_7756),
.Y(n_8407)
);

INVx1_ASAP7_75t_L g8408 ( 
.A(n_7768),
.Y(n_8408)
);

CKINVDCx5p33_ASAP7_75t_R g8409 ( 
.A(n_7769),
.Y(n_8409)
);

INVxp67_ASAP7_75t_L g8410 ( 
.A(n_7846),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_7770),
.Y(n_8411)
);

CKINVDCx20_ASAP7_75t_R g8412 ( 
.A(n_7771),
.Y(n_8412)
);

BUFx3_ASAP7_75t_L g8413 ( 
.A(n_7774),
.Y(n_8413)
);

INVx1_ASAP7_75t_L g8414 ( 
.A(n_7777),
.Y(n_8414)
);

INVx1_ASAP7_75t_L g8415 ( 
.A(n_7779),
.Y(n_8415)
);

INVx1_ASAP7_75t_L g8416 ( 
.A(n_7780),
.Y(n_8416)
);

INVxp67_ASAP7_75t_SL g8417 ( 
.A(n_7733),
.Y(n_8417)
);

CKINVDCx20_ASAP7_75t_R g8418 ( 
.A(n_7783),
.Y(n_8418)
);

INVx1_ASAP7_75t_L g8419 ( 
.A(n_7786),
.Y(n_8419)
);

CKINVDCx20_ASAP7_75t_R g8420 ( 
.A(n_7789),
.Y(n_8420)
);

INVxp67_ASAP7_75t_SL g8421 ( 
.A(n_7790),
.Y(n_8421)
);

INVxp67_ASAP7_75t_SL g8422 ( 
.A(n_7932),
.Y(n_8422)
);

INVx1_ASAP7_75t_L g8423 ( 
.A(n_7791),
.Y(n_8423)
);

CKINVDCx5p33_ASAP7_75t_R g8424 ( 
.A(n_7792),
.Y(n_8424)
);

INVxp67_ASAP7_75t_L g8425 ( 
.A(n_7821),
.Y(n_8425)
);

INVx1_ASAP7_75t_L g8426 ( 
.A(n_7793),
.Y(n_8426)
);

CKINVDCx20_ASAP7_75t_R g8427 ( 
.A(n_7794),
.Y(n_8427)
);

INVx1_ASAP7_75t_L g8428 ( 
.A(n_7795),
.Y(n_8428)
);

CKINVDCx5p33_ASAP7_75t_R g8429 ( 
.A(n_7797),
.Y(n_8429)
);

INVxp67_ASAP7_75t_SL g8430 ( 
.A(n_7824),
.Y(n_8430)
);

CKINVDCx5p33_ASAP7_75t_R g8431 ( 
.A(n_7799),
.Y(n_8431)
);

CKINVDCx5p33_ASAP7_75t_R g8432 ( 
.A(n_7802),
.Y(n_8432)
);

INVx1_ASAP7_75t_L g8433 ( 
.A(n_7806),
.Y(n_8433)
);

CKINVDCx5p33_ASAP7_75t_R g8434 ( 
.A(n_7808),
.Y(n_8434)
);

CKINVDCx5p33_ASAP7_75t_R g8435 ( 
.A(n_7809),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_7811),
.Y(n_8436)
);

INVx1_ASAP7_75t_L g8437 ( 
.A(n_7815),
.Y(n_8437)
);

HB1xp67_ASAP7_75t_L g8438 ( 
.A(n_7848),
.Y(n_8438)
);

CKINVDCx16_ASAP7_75t_R g8439 ( 
.A(n_7683),
.Y(n_8439)
);

INVx1_ASAP7_75t_L g8440 ( 
.A(n_7817),
.Y(n_8440)
);

CKINVDCx20_ASAP7_75t_R g8441 ( 
.A(n_7819),
.Y(n_8441)
);

CKINVDCx5p33_ASAP7_75t_R g8442 ( 
.A(n_7822),
.Y(n_8442)
);

CKINVDCx5p33_ASAP7_75t_R g8443 ( 
.A(n_7825),
.Y(n_8443)
);

INVxp67_ASAP7_75t_L g8444 ( 
.A(n_7995),
.Y(n_8444)
);

CKINVDCx20_ASAP7_75t_R g8445 ( 
.A(n_7826),
.Y(n_8445)
);

HB1xp67_ASAP7_75t_L g8446 ( 
.A(n_7829),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_7830),
.Y(n_8447)
);

CKINVDCx14_ASAP7_75t_R g8448 ( 
.A(n_7710),
.Y(n_8448)
);

HB1xp67_ASAP7_75t_L g8449 ( 
.A(n_7832),
.Y(n_8449)
);

CKINVDCx5p33_ASAP7_75t_R g8450 ( 
.A(n_7833),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_7835),
.Y(n_8451)
);

CKINVDCx5p33_ASAP7_75t_R g8452 ( 
.A(n_7836),
.Y(n_8452)
);

INVxp67_ASAP7_75t_L g8453 ( 
.A(n_7668),
.Y(n_8453)
);

CKINVDCx5p33_ASAP7_75t_R g8454 ( 
.A(n_7841),
.Y(n_8454)
);

HB1xp67_ASAP7_75t_L g8455 ( 
.A(n_7844),
.Y(n_8455)
);

CKINVDCx16_ASAP7_75t_R g8456 ( 
.A(n_7734),
.Y(n_8456)
);

INVx1_ASAP7_75t_L g8457 ( 
.A(n_7845),
.Y(n_8457)
);

NOR2xp67_ASAP7_75t_L g8458 ( 
.A(n_8015),
.B(n_6824),
.Y(n_8458)
);

INVx1_ASAP7_75t_L g8459 ( 
.A(n_7847),
.Y(n_8459)
);

INVx1_ASAP7_75t_L g8460 ( 
.A(n_7855),
.Y(n_8460)
);

INVx1_ASAP7_75t_L g8461 ( 
.A(n_7858),
.Y(n_8461)
);

INVx1_ASAP7_75t_L g8462 ( 
.A(n_7859),
.Y(n_8462)
);

CKINVDCx20_ASAP7_75t_R g8463 ( 
.A(n_7861),
.Y(n_8463)
);

CKINVDCx5p33_ASAP7_75t_R g8464 ( 
.A(n_7864),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_7867),
.Y(n_8465)
);

INVx1_ASAP7_75t_L g8466 ( 
.A(n_7868),
.Y(n_8466)
);

INVx1_ASAP7_75t_L g8467 ( 
.A(n_7875),
.Y(n_8467)
);

INVx1_ASAP7_75t_L g8468 ( 
.A(n_7878),
.Y(n_8468)
);

INVx2_ASAP7_75t_L g8469 ( 
.A(n_7879),
.Y(n_8469)
);

CKINVDCx20_ASAP7_75t_R g8470 ( 
.A(n_7880),
.Y(n_8470)
);

INVx1_ASAP7_75t_L g8471 ( 
.A(n_7881),
.Y(n_8471)
);

CKINVDCx5p33_ASAP7_75t_R g8472 ( 
.A(n_7886),
.Y(n_8472)
);

INVxp67_ASAP7_75t_L g8473 ( 
.A(n_7668),
.Y(n_8473)
);

INVxp67_ASAP7_75t_SL g8474 ( 
.A(n_7726),
.Y(n_8474)
);

CKINVDCx5p33_ASAP7_75t_R g8475 ( 
.A(n_7888),
.Y(n_8475)
);

INVx1_ASAP7_75t_L g8476 ( 
.A(n_7889),
.Y(n_8476)
);

INVx1_ASAP7_75t_L g8477 ( 
.A(n_7890),
.Y(n_8477)
);

INVx1_ASAP7_75t_L g8478 ( 
.A(n_7891),
.Y(n_8478)
);

INVx1_ASAP7_75t_L g8479 ( 
.A(n_7896),
.Y(n_8479)
);

INVx1_ASAP7_75t_L g8480 ( 
.A(n_7899),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_7900),
.Y(n_8481)
);

CKINVDCx16_ASAP7_75t_R g8482 ( 
.A(n_7781),
.Y(n_8482)
);

BUFx2_ASAP7_75t_L g8483 ( 
.A(n_7901),
.Y(n_8483)
);

INVx1_ASAP7_75t_L g8484 ( 
.A(n_7904),
.Y(n_8484)
);

BUFx6f_ASAP7_75t_L g8485 ( 
.A(n_7781),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_7907),
.Y(n_8486)
);

INVx1_ASAP7_75t_L g8487 ( 
.A(n_7908),
.Y(n_8487)
);

CKINVDCx5p33_ASAP7_75t_R g8488 ( 
.A(n_7910),
.Y(n_8488)
);

HB1xp67_ASAP7_75t_L g8489 ( 
.A(n_7911),
.Y(n_8489)
);

CKINVDCx5p33_ASAP7_75t_R g8490 ( 
.A(n_7912),
.Y(n_8490)
);

INVxp67_ASAP7_75t_SL g8491 ( 
.A(n_7916),
.Y(n_8491)
);

INVx1_ASAP7_75t_L g8492 ( 
.A(n_7921),
.Y(n_8492)
);

INVxp67_ASAP7_75t_L g8493 ( 
.A(n_7816),
.Y(n_8493)
);

INVx1_ASAP7_75t_L g8494 ( 
.A(n_7922),
.Y(n_8494)
);

CKINVDCx20_ASAP7_75t_R g8495 ( 
.A(n_7927),
.Y(n_8495)
);

CKINVDCx20_ASAP7_75t_R g8496 ( 
.A(n_7929),
.Y(n_8496)
);

INVxp67_ASAP7_75t_L g8497 ( 
.A(n_7816),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_7937),
.Y(n_8498)
);

INVx2_ASAP7_75t_L g8499 ( 
.A(n_7940),
.Y(n_8499)
);

INVx1_ASAP7_75t_L g8500 ( 
.A(n_7943),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7945),
.Y(n_8501)
);

CKINVDCx5p33_ASAP7_75t_R g8502 ( 
.A(n_7948),
.Y(n_8502)
);

CKINVDCx5p33_ASAP7_75t_R g8503 ( 
.A(n_7949),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_7951),
.Y(n_8504)
);

INVx1_ASAP7_75t_L g8505 ( 
.A(n_7954),
.Y(n_8505)
);

CKINVDCx20_ASAP7_75t_R g8506 ( 
.A(n_7963),
.Y(n_8506)
);

INVxp33_ASAP7_75t_L g8507 ( 
.A(n_7798),
.Y(n_8507)
);

HB1xp67_ASAP7_75t_L g8508 ( 
.A(n_7964),
.Y(n_8508)
);

BUFx3_ASAP7_75t_L g8509 ( 
.A(n_7965),
.Y(n_8509)
);

INVx1_ASAP7_75t_L g8510 ( 
.A(n_7966),
.Y(n_8510)
);

INVx1_ASAP7_75t_SL g8511 ( 
.A(n_7967),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_7970),
.Y(n_8512)
);

INVxp67_ASAP7_75t_L g8513 ( 
.A(n_7971),
.Y(n_8513)
);

INVxp33_ASAP7_75t_L g8514 ( 
.A(n_7973),
.Y(n_8514)
);

CKINVDCx20_ASAP7_75t_R g8515 ( 
.A(n_7974),
.Y(n_8515)
);

CKINVDCx5p33_ASAP7_75t_R g8516 ( 
.A(n_7978),
.Y(n_8516)
);

INVx1_ASAP7_75t_L g8517 ( 
.A(n_7979),
.Y(n_8517)
);

INVx1_ASAP7_75t_L g8518 ( 
.A(n_7981),
.Y(n_8518)
);

INVx1_ASAP7_75t_L g8519 ( 
.A(n_7982),
.Y(n_8519)
);

INVx1_ASAP7_75t_L g8520 ( 
.A(n_7767),
.Y(n_8520)
);

NOR2xp67_ASAP7_75t_L g8521 ( 
.A(n_8015),
.B(n_6201),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_7767),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_7767),
.Y(n_8523)
);

INVx1_ASAP7_75t_L g8524 ( 
.A(n_7767),
.Y(n_8524)
);

INVxp67_ASAP7_75t_SL g8525 ( 
.A(n_7553),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_7767),
.Y(n_8526)
);

INVxp67_ASAP7_75t_L g8527 ( 
.A(n_7560),
.Y(n_8527)
);

INVx1_ASAP7_75t_L g8528 ( 
.A(n_7767),
.Y(n_8528)
);

BUFx3_ASAP7_75t_L g8529 ( 
.A(n_7860),
.Y(n_8529)
);

INVx1_ASAP7_75t_L g8530 ( 
.A(n_7767),
.Y(n_8530)
);

INVxp67_ASAP7_75t_SL g8531 ( 
.A(n_7553),
.Y(n_8531)
);

CKINVDCx14_ASAP7_75t_R g8532 ( 
.A(n_7592),
.Y(n_8532)
);

INVx1_ASAP7_75t_L g8533 ( 
.A(n_7767),
.Y(n_8533)
);

INVx2_ASAP7_75t_L g8534 ( 
.A(n_7767),
.Y(n_8534)
);

NAND2xp5_ASAP7_75t_L g8535 ( 
.A(n_7562),
.B(n_7044),
.Y(n_8535)
);

INVx1_ASAP7_75t_L g8536 ( 
.A(n_7767),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_7767),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_7767),
.Y(n_8538)
);

CKINVDCx20_ASAP7_75t_R g8539 ( 
.A(n_7547),
.Y(n_8539)
);

CKINVDCx5p33_ASAP7_75t_R g8540 ( 
.A(n_7562),
.Y(n_8540)
);

INVx1_ASAP7_75t_L g8541 ( 
.A(n_7767),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_7767),
.Y(n_8542)
);

BUFx3_ASAP7_75t_L g8543 ( 
.A(n_7860),
.Y(n_8543)
);

INVx2_ASAP7_75t_L g8544 ( 
.A(n_7767),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_7767),
.Y(n_8545)
);

INVx1_ASAP7_75t_L g8546 ( 
.A(n_7767),
.Y(n_8546)
);

INVxp67_ASAP7_75t_SL g8547 ( 
.A(n_7553),
.Y(n_8547)
);

INVxp67_ASAP7_75t_SL g8548 ( 
.A(n_7553),
.Y(n_8548)
);

CKINVDCx5p33_ASAP7_75t_R g8549 ( 
.A(n_8017),
.Y(n_8549)
);

INVx2_ASAP7_75t_L g8550 ( 
.A(n_8153),
.Y(n_8550)
);

INVx1_ASAP7_75t_L g8551 ( 
.A(n_8238),
.Y(n_8551)
);

OAI22xp5_ASAP7_75t_L g8552 ( 
.A1(n_8156),
.A2(n_7436),
.B1(n_7367),
.B2(n_6891),
.Y(n_8552)
);

INVx2_ASAP7_75t_L g8553 ( 
.A(n_8153),
.Y(n_8553)
);

OAI22x1_ASAP7_75t_SL g8554 ( 
.A1(n_8199),
.A2(n_6100),
.B1(n_6137),
.B2(n_6091),
.Y(n_8554)
);

BUFx6f_ASAP7_75t_L g8555 ( 
.A(n_8044),
.Y(n_8555)
);

NAND2xp5_ASAP7_75t_L g8556 ( 
.A(n_8162),
.B(n_6500),
.Y(n_8556)
);

INVx2_ASAP7_75t_L g8557 ( 
.A(n_8153),
.Y(n_8557)
);

NOR2xp33_ASAP7_75t_SL g8558 ( 
.A(n_8425),
.B(n_7208),
.Y(n_8558)
);

HB1xp67_ASAP7_75t_L g8559 ( 
.A(n_8392),
.Y(n_8559)
);

INVx2_ASAP7_75t_L g8560 ( 
.A(n_8100),
.Y(n_8560)
);

BUFx6f_ASAP7_75t_L g8561 ( 
.A(n_8044),
.Y(n_8561)
);

INVx6_ASAP7_75t_L g8562 ( 
.A(n_8485),
.Y(n_8562)
);

OAI21x1_ASAP7_75t_L g8563 ( 
.A1(n_8326),
.A2(n_6195),
.B(n_6165),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_8239),
.Y(n_8564)
);

INVx1_ASAP7_75t_L g8565 ( 
.A(n_8240),
.Y(n_8565)
);

BUFx6f_ASAP7_75t_L g8566 ( 
.A(n_8098),
.Y(n_8566)
);

AND2x4_ASAP7_75t_L g8567 ( 
.A(n_8237),
.B(n_8152),
.Y(n_8567)
);

AND2x4_ASAP7_75t_L g8568 ( 
.A(n_8078),
.B(n_6196),
.Y(n_8568)
);

INVx1_ASAP7_75t_L g8569 ( 
.A(n_8241),
.Y(n_8569)
);

INVx1_ASAP7_75t_L g8570 ( 
.A(n_8243),
.Y(n_8570)
);

AND2x4_ASAP7_75t_L g8571 ( 
.A(n_8084),
.B(n_8128),
.Y(n_8571)
);

CKINVDCx16_ASAP7_75t_R g8572 ( 
.A(n_8075),
.Y(n_8572)
);

AND2x2_ASAP7_75t_L g8573 ( 
.A(n_8430),
.B(n_7365),
.Y(n_8573)
);

AND2x4_ASAP7_75t_L g8574 ( 
.A(n_8529),
.B(n_8543),
.Y(n_8574)
);

INVx3_ASAP7_75t_L g8575 ( 
.A(n_8098),
.Y(n_8575)
);

INVx2_ASAP7_75t_L g8576 ( 
.A(n_8534),
.Y(n_8576)
);

INVx1_ASAP7_75t_L g8577 ( 
.A(n_8247),
.Y(n_8577)
);

NAND2xp5_ASAP7_75t_L g8578 ( 
.A(n_8535),
.B(n_6587),
.Y(n_8578)
);

CKINVDCx6p67_ASAP7_75t_R g8579 ( 
.A(n_8387),
.Y(n_8579)
);

INVx4_ASAP7_75t_L g8580 ( 
.A(n_8021),
.Y(n_8580)
);

INVx1_ASAP7_75t_L g8581 ( 
.A(n_8252),
.Y(n_8581)
);

NAND2xp5_ASAP7_75t_L g8582 ( 
.A(n_8344),
.B(n_6803),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_8253),
.Y(n_8583)
);

INVx2_ASAP7_75t_SL g8584 ( 
.A(n_8407),
.Y(n_8584)
);

BUFx6f_ASAP7_75t_L g8585 ( 
.A(n_8249),
.Y(n_8585)
);

INVx1_ASAP7_75t_L g8586 ( 
.A(n_8257),
.Y(n_8586)
);

BUFx6f_ASAP7_75t_L g8587 ( 
.A(n_8286),
.Y(n_8587)
);

INVx3_ASAP7_75t_L g8588 ( 
.A(n_8158),
.Y(n_8588)
);

BUFx6f_ASAP7_75t_L g8589 ( 
.A(n_8122),
.Y(n_8589)
);

INVx6_ASAP7_75t_L g8590 ( 
.A(n_8485),
.Y(n_8590)
);

NAND2xp5_ASAP7_75t_L g8591 ( 
.A(n_8348),
.B(n_6902),
.Y(n_8591)
);

INVx2_ASAP7_75t_L g8592 ( 
.A(n_8544),
.Y(n_8592)
);

BUFx8_ASAP7_75t_L g8593 ( 
.A(n_8485),
.Y(n_8593)
);

INVx2_ASAP7_75t_L g8594 ( 
.A(n_8161),
.Y(n_8594)
);

INVx1_ASAP7_75t_L g8595 ( 
.A(n_8262),
.Y(n_8595)
);

AND2x4_ASAP7_75t_L g8596 ( 
.A(n_8370),
.B(n_6469),
.Y(n_8596)
);

OA21x2_ASAP7_75t_L g8597 ( 
.A1(n_8327),
.A2(n_6615),
.B(n_6567),
.Y(n_8597)
);

HB1xp67_ASAP7_75t_L g8598 ( 
.A(n_8438),
.Y(n_8598)
);

NAND2xp5_ASAP7_75t_L g8599 ( 
.A(n_8038),
.B(n_7136),
.Y(n_8599)
);

INVx2_ASAP7_75t_L g8600 ( 
.A(n_8164),
.Y(n_8600)
);

INVx2_ASAP7_75t_L g8601 ( 
.A(n_8198),
.Y(n_8601)
);

BUFx2_ASAP7_75t_L g8602 ( 
.A(n_8206),
.Y(n_8602)
);

HB1xp67_ASAP7_75t_L g8603 ( 
.A(n_8250),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_8263),
.Y(n_8604)
);

CKINVDCx6p67_ASAP7_75t_R g8605 ( 
.A(n_8439),
.Y(n_8605)
);

BUFx6f_ASAP7_75t_L g8606 ( 
.A(n_8123),
.Y(n_8606)
);

AOI22xp5_ASAP7_75t_L g8607 ( 
.A1(n_8298),
.A2(n_6257),
.B1(n_6471),
.B2(n_6176),
.Y(n_8607)
);

INVx2_ASAP7_75t_L g8608 ( 
.A(n_8205),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8264),
.Y(n_8609)
);

INVx1_ASAP7_75t_L g8610 ( 
.A(n_8265),
.Y(n_8610)
);

INVx2_ASAP7_75t_L g8611 ( 
.A(n_8207),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_8266),
.Y(n_8612)
);

INVx2_ASAP7_75t_L g8613 ( 
.A(n_8254),
.Y(n_8613)
);

INVx2_ASAP7_75t_L g8614 ( 
.A(n_8272),
.Y(n_8614)
);

CKINVDCx20_ASAP7_75t_R g8615 ( 
.A(n_8063),
.Y(n_8615)
);

BUFx6f_ASAP7_75t_L g8616 ( 
.A(n_8124),
.Y(n_8616)
);

BUFx3_ASAP7_75t_L g8617 ( 
.A(n_8371),
.Y(n_8617)
);

AOI22xp33_ASAP7_75t_L g8618 ( 
.A1(n_8347),
.A2(n_6080),
.B1(n_6173),
.B2(n_6110),
.Y(n_8618)
);

NAND2xp5_ASAP7_75t_L g8619 ( 
.A(n_8064),
.B(n_8071),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_8300),
.Y(n_8620)
);

CKINVDCx5p33_ASAP7_75t_R g8621 ( 
.A(n_8049),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_8267),
.Y(n_8622)
);

BUFx3_ASAP7_75t_L g8623 ( 
.A(n_8413),
.Y(n_8623)
);

INVx2_ASAP7_75t_L g8624 ( 
.A(n_8125),
.Y(n_8624)
);

NAND2xp5_ASAP7_75t_L g8625 ( 
.A(n_8073),
.B(n_6538),
.Y(n_8625)
);

BUFx6f_ASAP7_75t_L g8626 ( 
.A(n_8129),
.Y(n_8626)
);

BUFx12f_ASAP7_75t_L g8627 ( 
.A(n_8059),
.Y(n_8627)
);

BUFx6f_ASAP7_75t_L g8628 ( 
.A(n_8131),
.Y(n_8628)
);

AND2x4_ASAP7_75t_L g8629 ( 
.A(n_8373),
.B(n_6546),
.Y(n_8629)
);

INVxp67_ASAP7_75t_L g8630 ( 
.A(n_8342),
.Y(n_8630)
);

AND2x4_ASAP7_75t_L g8631 ( 
.A(n_8376),
.B(n_6639),
.Y(n_8631)
);

INVx2_ASAP7_75t_L g8632 ( 
.A(n_8132),
.Y(n_8632)
);

AND2x4_ASAP7_75t_L g8633 ( 
.A(n_8379),
.B(n_6642),
.Y(n_8633)
);

BUFx3_ASAP7_75t_L g8634 ( 
.A(n_8509),
.Y(n_8634)
);

INVx1_ASAP7_75t_L g8635 ( 
.A(n_8273),
.Y(n_8635)
);

INVx2_ASAP7_75t_L g8636 ( 
.A(n_8133),
.Y(n_8636)
);

INVx2_ASAP7_75t_L g8637 ( 
.A(n_8136),
.Y(n_8637)
);

INVx2_ASAP7_75t_L g8638 ( 
.A(n_8137),
.Y(n_8638)
);

INVx2_ASAP7_75t_SL g8639 ( 
.A(n_8329),
.Y(n_8639)
);

NAND2xp5_ASAP7_75t_L g8640 ( 
.A(n_8092),
.B(n_6645),
.Y(n_8640)
);

NOR2xp33_ASAP7_75t_L g8641 ( 
.A(n_8383),
.B(n_6765),
.Y(n_8641)
);

NAND2xp5_ASAP7_75t_L g8642 ( 
.A(n_8102),
.B(n_6786),
.Y(n_8642)
);

INVx1_ASAP7_75t_L g8643 ( 
.A(n_8274),
.Y(n_8643)
);

INVxp67_ASAP7_75t_L g8644 ( 
.A(n_8187),
.Y(n_8644)
);

AND2x4_ASAP7_75t_L g8645 ( 
.A(n_8380),
.B(n_6928),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_8275),
.Y(n_8646)
);

INVx2_ASAP7_75t_L g8647 ( 
.A(n_8140),
.Y(n_8647)
);

NOR2x1_ASAP7_75t_L g8648 ( 
.A(n_8384),
.B(n_6117),
.Y(n_8648)
);

INVx3_ASAP7_75t_L g8649 ( 
.A(n_8141),
.Y(n_8649)
);

BUFx6f_ASAP7_75t_L g8650 ( 
.A(n_8143),
.Y(n_8650)
);

BUFx6f_ASAP7_75t_L g8651 ( 
.A(n_8144),
.Y(n_8651)
);

NAND2xp5_ASAP7_75t_L g8652 ( 
.A(n_8126),
.B(n_6859),
.Y(n_8652)
);

INVx2_ASAP7_75t_L g8653 ( 
.A(n_8145),
.Y(n_8653)
);

AOI22xp5_ASAP7_75t_L g8654 ( 
.A1(n_8336),
.A2(n_7108),
.B1(n_7311),
.B2(n_6952),
.Y(n_8654)
);

INVx3_ASAP7_75t_L g8655 ( 
.A(n_8147),
.Y(n_8655)
);

NOR2xp33_ASAP7_75t_L g8656 ( 
.A(n_8385),
.B(n_7314),
.Y(n_8656)
);

INVx2_ASAP7_75t_L g8657 ( 
.A(n_8149),
.Y(n_8657)
);

INVx1_ASAP7_75t_L g8658 ( 
.A(n_8276),
.Y(n_8658)
);

CKINVDCx5p33_ASAP7_75t_R g8659 ( 
.A(n_8066),
.Y(n_8659)
);

INVx2_ASAP7_75t_SL g8660 ( 
.A(n_8329),
.Y(n_8660)
);

INVx1_ASAP7_75t_L g8661 ( 
.A(n_8277),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_8278),
.Y(n_8662)
);

NOR2xp33_ASAP7_75t_L g8663 ( 
.A(n_8386),
.B(n_8388),
.Y(n_8663)
);

BUFx6f_ASAP7_75t_L g8664 ( 
.A(n_8150),
.Y(n_8664)
);

INVx2_ASAP7_75t_L g8665 ( 
.A(n_8019),
.Y(n_8665)
);

INVx3_ASAP7_75t_L g8666 ( 
.A(n_8329),
.Y(n_8666)
);

OAI21x1_ASAP7_75t_L g8667 ( 
.A1(n_8328),
.A2(n_6857),
.B(n_6847),
.Y(n_8667)
);

OA21x2_ASAP7_75t_L g8668 ( 
.A1(n_8333),
.A2(n_7004),
.B(n_6868),
.Y(n_8668)
);

INVx1_ASAP7_75t_L g8669 ( 
.A(n_8281),
.Y(n_8669)
);

INVx2_ASAP7_75t_L g8670 ( 
.A(n_8020),
.Y(n_8670)
);

BUFx12f_ASAP7_75t_L g8671 ( 
.A(n_8069),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_8022),
.Y(n_8672)
);

INVx3_ASAP7_75t_L g8673 ( 
.A(n_8282),
.Y(n_8673)
);

AOI22x1_ASAP7_75t_SL g8674 ( 
.A1(n_8474),
.A2(n_6250),
.B1(n_6279),
.B2(n_6204),
.Y(n_8674)
);

OA21x2_ASAP7_75t_L g8675 ( 
.A1(n_8334),
.A2(n_7110),
.B(n_7034),
.Y(n_8675)
);

INVxp33_ASAP7_75t_SL g8676 ( 
.A(n_8287),
.Y(n_8676)
);

NAND2xp5_ASAP7_75t_L g8677 ( 
.A(n_8127),
.B(n_7461),
.Y(n_8677)
);

INVx3_ASAP7_75t_L g8678 ( 
.A(n_8284),
.Y(n_8678)
);

BUFx6f_ASAP7_75t_L g8679 ( 
.A(n_8288),
.Y(n_8679)
);

OA21x2_ASAP7_75t_L g8680 ( 
.A1(n_8338),
.A2(n_7309),
.B(n_7144),
.Y(n_8680)
);

CKINVDCx5p33_ASAP7_75t_R g8681 ( 
.A(n_8082),
.Y(n_8681)
);

BUFx6f_ASAP7_75t_L g8682 ( 
.A(n_8289),
.Y(n_8682)
);

BUFx6f_ASAP7_75t_L g8683 ( 
.A(n_8291),
.Y(n_8683)
);

AND2x2_ASAP7_75t_L g8684 ( 
.A(n_8222),
.B(n_6285),
.Y(n_8684)
);

INVx5_ASAP7_75t_L g8685 ( 
.A(n_8219),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_8292),
.Y(n_8686)
);

INVx2_ASAP7_75t_L g8687 ( 
.A(n_8023),
.Y(n_8687)
);

INVx1_ASAP7_75t_L g8688 ( 
.A(n_8293),
.Y(n_8688)
);

INVx2_ASAP7_75t_L g8689 ( 
.A(n_8024),
.Y(n_8689)
);

AND2x2_ASAP7_75t_SL g8690 ( 
.A(n_8233),
.B(n_6225),
.Y(n_8690)
);

HB1xp67_ASAP7_75t_L g8691 ( 
.A(n_8314),
.Y(n_8691)
);

INVx2_ASAP7_75t_L g8692 ( 
.A(n_8025),
.Y(n_8692)
);

BUFx6f_ASAP7_75t_L g8693 ( 
.A(n_8294),
.Y(n_8693)
);

INVx2_ASAP7_75t_SL g8694 ( 
.A(n_8345),
.Y(n_8694)
);

BUFx6f_ASAP7_75t_L g8695 ( 
.A(n_8299),
.Y(n_8695)
);

INVx1_ASAP7_75t_L g8696 ( 
.A(n_8303),
.Y(n_8696)
);

AND2x6_ASAP7_75t_L g8697 ( 
.A(n_8389),
.B(n_6077),
.Y(n_8697)
);

BUFx2_ASAP7_75t_L g8698 ( 
.A(n_8381),
.Y(n_8698)
);

INVx2_ASAP7_75t_L g8699 ( 
.A(n_8026),
.Y(n_8699)
);

AND2x4_ASAP7_75t_L g8700 ( 
.A(n_8469),
.B(n_7015),
.Y(n_8700)
);

INVx1_ASAP7_75t_L g8701 ( 
.A(n_8304),
.Y(n_8701)
);

INVx2_ASAP7_75t_L g8702 ( 
.A(n_8028),
.Y(n_8702)
);

INVx2_ASAP7_75t_L g8703 ( 
.A(n_8029),
.Y(n_8703)
);

INVx1_ASAP7_75t_L g8704 ( 
.A(n_8305),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_8030),
.Y(n_8705)
);

NOR2xp33_ASAP7_75t_L g8706 ( 
.A(n_8390),
.B(n_7487),
.Y(n_8706)
);

INVx2_ASAP7_75t_SL g8707 ( 
.A(n_8363),
.Y(n_8707)
);

OA21x2_ASAP7_75t_L g8708 ( 
.A1(n_8340),
.A2(n_7409),
.B(n_6136),
.Y(n_8708)
);

BUFx12f_ASAP7_75t_L g8709 ( 
.A(n_8085),
.Y(n_8709)
);

BUFx6f_ASAP7_75t_L g8710 ( 
.A(n_8033),
.Y(n_8710)
);

INVx2_ASAP7_75t_L g8711 ( 
.A(n_8034),
.Y(n_8711)
);

BUFx12f_ASAP7_75t_L g8712 ( 
.A(n_8087),
.Y(n_8712)
);

OAI21x1_ASAP7_75t_L g8713 ( 
.A1(n_8330),
.A2(n_6157),
.B(n_6122),
.Y(n_8713)
);

INVx3_ASAP7_75t_L g8714 ( 
.A(n_8151),
.Y(n_8714)
);

INVxp67_ASAP7_75t_L g8715 ( 
.A(n_8349),
.Y(n_8715)
);

BUFx8_ASAP7_75t_L g8716 ( 
.A(n_8031),
.Y(n_8716)
);

BUFx6f_ASAP7_75t_L g8717 ( 
.A(n_8035),
.Y(n_8717)
);

INVx6_ASAP7_75t_L g8718 ( 
.A(n_8245),
.Y(n_8718)
);

BUFx8_ASAP7_75t_L g8719 ( 
.A(n_8047),
.Y(n_8719)
);

NAND2xp5_ASAP7_75t_L g8720 ( 
.A(n_8142),
.B(n_6313),
.Y(n_8720)
);

BUFx6f_ASAP7_75t_L g8721 ( 
.A(n_8037),
.Y(n_8721)
);

AND2x4_ASAP7_75t_L g8722 ( 
.A(n_8499),
.B(n_7244),
.Y(n_8722)
);

BUFx3_ASAP7_75t_L g8723 ( 
.A(n_8412),
.Y(n_8723)
);

CKINVDCx5p33_ASAP7_75t_R g8724 ( 
.A(n_8095),
.Y(n_8724)
);

NAND2xp5_ASAP7_75t_L g8725 ( 
.A(n_8525),
.B(n_6454),
.Y(n_8725)
);

NAND2xp5_ASAP7_75t_L g8726 ( 
.A(n_8531),
.B(n_8547),
.Y(n_8726)
);

OAI22xp5_ASAP7_75t_L g8727 ( 
.A1(n_8421),
.A2(n_6081),
.B1(n_6083),
.B2(n_6079),
.Y(n_8727)
);

INVx2_ASAP7_75t_L g8728 ( 
.A(n_8039),
.Y(n_8728)
);

BUFx2_ASAP7_75t_L g8729 ( 
.A(n_8410),
.Y(n_8729)
);

AND2x2_ASAP7_75t_L g8730 ( 
.A(n_8307),
.B(n_6285),
.Y(n_8730)
);

BUFx2_ASAP7_75t_L g8731 ( 
.A(n_8269),
.Y(n_8731)
);

AND2x4_ASAP7_75t_L g8732 ( 
.A(n_8347),
.B(n_7408),
.Y(n_8732)
);

OAI21x1_ASAP7_75t_L g8733 ( 
.A1(n_8335),
.A2(n_6209),
.B(n_6178),
.Y(n_8733)
);

INVx2_ASAP7_75t_L g8734 ( 
.A(n_8041),
.Y(n_8734)
);

INVx1_ASAP7_75t_L g8735 ( 
.A(n_8154),
.Y(n_8735)
);

AND2x4_ASAP7_75t_L g8736 ( 
.A(n_8332),
.B(n_7458),
.Y(n_8736)
);

OA21x2_ASAP7_75t_L g8737 ( 
.A1(n_8343),
.A2(n_6230),
.B(n_6221),
.Y(n_8737)
);

CKINVDCx5p33_ASAP7_75t_R g8738 ( 
.A(n_8104),
.Y(n_8738)
);

AND2x2_ASAP7_75t_L g8739 ( 
.A(n_8313),
.B(n_6413),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_8155),
.Y(n_8740)
);

INVx1_ASAP7_75t_L g8741 ( 
.A(n_8160),
.Y(n_8741)
);

INVx1_ASAP7_75t_L g8742 ( 
.A(n_8169),
.Y(n_8742)
);

INVx2_ASAP7_75t_L g8743 ( 
.A(n_8042),
.Y(n_8743)
);

BUFx6f_ASAP7_75t_L g8744 ( 
.A(n_8045),
.Y(n_8744)
);

BUFx6f_ASAP7_75t_L g8745 ( 
.A(n_8046),
.Y(n_8745)
);

INVx2_ASAP7_75t_L g8746 ( 
.A(n_8048),
.Y(n_8746)
);

INVx2_ASAP7_75t_L g8747 ( 
.A(n_8050),
.Y(n_8747)
);

INVx1_ASAP7_75t_L g8748 ( 
.A(n_8172),
.Y(n_8748)
);

INVx2_ASAP7_75t_L g8749 ( 
.A(n_8051),
.Y(n_8749)
);

NOR2xp33_ASAP7_75t_L g8750 ( 
.A(n_8396),
.B(n_7496),
.Y(n_8750)
);

INVx1_ASAP7_75t_L g8751 ( 
.A(n_8175),
.Y(n_8751)
);

BUFx6f_ASAP7_75t_L g8752 ( 
.A(n_8052),
.Y(n_8752)
);

INVx2_ASAP7_75t_L g8753 ( 
.A(n_8053),
.Y(n_8753)
);

INVx2_ASAP7_75t_L g8754 ( 
.A(n_8054),
.Y(n_8754)
);

CKINVDCx20_ASAP7_75t_R g8755 ( 
.A(n_8068),
.Y(n_8755)
);

INVx5_ASAP7_75t_L g8756 ( 
.A(n_8270),
.Y(n_8756)
);

OA21x2_ASAP7_75t_L g8757 ( 
.A1(n_8177),
.A2(n_6233),
.B(n_6231),
.Y(n_8757)
);

INVx4_ASAP7_75t_L g8758 ( 
.A(n_8114),
.Y(n_8758)
);

BUFx6f_ASAP7_75t_L g8759 ( 
.A(n_8055),
.Y(n_8759)
);

BUFx2_ASAP7_75t_L g8760 ( 
.A(n_8036),
.Y(n_8760)
);

INVx2_ASAP7_75t_L g8761 ( 
.A(n_8056),
.Y(n_8761)
);

INVx1_ASAP7_75t_L g8762 ( 
.A(n_8178),
.Y(n_8762)
);

OAI22xp5_ASAP7_75t_SL g8763 ( 
.A1(n_8310),
.A2(n_6331),
.B1(n_6343),
.B2(n_6299),
.Y(n_8763)
);

AND2x2_ASAP7_75t_L g8764 ( 
.A(n_8341),
.B(n_6413),
.Y(n_8764)
);

BUFx6f_ASAP7_75t_L g8765 ( 
.A(n_8057),
.Y(n_8765)
);

INVx3_ASAP7_75t_L g8766 ( 
.A(n_8180),
.Y(n_8766)
);

CKINVDCx11_ASAP7_75t_R g8767 ( 
.A(n_8090),
.Y(n_8767)
);

INVx3_ASAP7_75t_L g8768 ( 
.A(n_8181),
.Y(n_8768)
);

INVx1_ASAP7_75t_L g8769 ( 
.A(n_8182),
.Y(n_8769)
);

BUFx6f_ASAP7_75t_L g8770 ( 
.A(n_8058),
.Y(n_8770)
);

AND2x4_ASAP7_75t_L g8771 ( 
.A(n_8398),
.B(n_6977),
.Y(n_8771)
);

BUFx6f_ASAP7_75t_L g8772 ( 
.A(n_8060),
.Y(n_8772)
);

BUFx3_ASAP7_75t_L g8773 ( 
.A(n_8418),
.Y(n_8773)
);

OAI22x1_ASAP7_75t_SL g8774 ( 
.A1(n_8094),
.A2(n_6428),
.B1(n_6444),
.B2(n_6360),
.Y(n_8774)
);

INVx2_ASAP7_75t_L g8775 ( 
.A(n_8061),
.Y(n_8775)
);

INVx2_ASAP7_75t_SL g8776 ( 
.A(n_8394),
.Y(n_8776)
);

INVx1_ASAP7_75t_L g8777 ( 
.A(n_8193),
.Y(n_8777)
);

BUFx6f_ASAP7_75t_L g8778 ( 
.A(n_8062),
.Y(n_8778)
);

BUFx6f_ASAP7_75t_L g8779 ( 
.A(n_8065),
.Y(n_8779)
);

INVx1_ASAP7_75t_L g8780 ( 
.A(n_8194),
.Y(n_8780)
);

CKINVDCx20_ASAP7_75t_R g8781 ( 
.A(n_8116),
.Y(n_8781)
);

AND2x2_ASAP7_75t_L g8782 ( 
.A(n_8367),
.B(n_6558),
.Y(n_8782)
);

AND2x2_ASAP7_75t_L g8783 ( 
.A(n_8378),
.B(n_8417),
.Y(n_8783)
);

INVx1_ASAP7_75t_L g8784 ( 
.A(n_8197),
.Y(n_8784)
);

OA21x2_ASAP7_75t_L g8785 ( 
.A1(n_8200),
.A2(n_6269),
.B(n_6263),
.Y(n_8785)
);

INVx2_ASAP7_75t_L g8786 ( 
.A(n_8067),
.Y(n_8786)
);

INVx1_ASAP7_75t_L g8787 ( 
.A(n_8202),
.Y(n_8787)
);

INVx3_ASAP7_75t_L g8788 ( 
.A(n_8203),
.Y(n_8788)
);

NAND2xp5_ASAP7_75t_SL g8789 ( 
.A(n_8511),
.B(n_7460),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_8548),
.B(n_7001),
.Y(n_8790)
);

INVxp67_ASAP7_75t_L g8791 ( 
.A(n_8422),
.Y(n_8791)
);

INVx2_ASAP7_75t_L g8792 ( 
.A(n_8070),
.Y(n_8792)
);

BUFx6f_ASAP7_75t_L g8793 ( 
.A(n_8074),
.Y(n_8793)
);

AOI22xp5_ASAP7_75t_L g8794 ( 
.A1(n_8400),
.A2(n_8406),
.B1(n_8408),
.B2(n_8402),
.Y(n_8794)
);

INVx3_ASAP7_75t_L g8795 ( 
.A(n_8204),
.Y(n_8795)
);

INVx1_ASAP7_75t_L g8796 ( 
.A(n_8209),
.Y(n_8796)
);

AND2x4_ASAP7_75t_L g8797 ( 
.A(n_8411),
.B(n_7183),
.Y(n_8797)
);

BUFx2_ASAP7_75t_L g8798 ( 
.A(n_8101),
.Y(n_8798)
);

OAI21x1_ASAP7_75t_L g8799 ( 
.A1(n_8210),
.A2(n_6301),
.B(n_6283),
.Y(n_8799)
);

BUFx6f_ASAP7_75t_L g8800 ( 
.A(n_8076),
.Y(n_8800)
);

BUFx8_ASAP7_75t_L g8801 ( 
.A(n_8188),
.Y(n_8801)
);

BUFx6f_ASAP7_75t_L g8802 ( 
.A(n_8077),
.Y(n_8802)
);

AND2x2_ASAP7_75t_L g8803 ( 
.A(n_8285),
.B(n_6558),
.Y(n_8803)
);

NAND2xp5_ASAP7_75t_SL g8804 ( 
.A(n_8456),
.B(n_7460),
.Y(n_8804)
);

XNOR2x2_ASAP7_75t_L g8805 ( 
.A(n_8404),
.B(n_6437),
.Y(n_8805)
);

BUFx6f_ASAP7_75t_L g8806 ( 
.A(n_8079),
.Y(n_8806)
);

XOR2xp5_ASAP7_75t_L g8807 ( 
.A(n_8138),
.B(n_6457),
.Y(n_8807)
);

BUFx6f_ASAP7_75t_L g8808 ( 
.A(n_8081),
.Y(n_8808)
);

INVx3_ASAP7_75t_L g8809 ( 
.A(n_8213),
.Y(n_8809)
);

AND2x6_ASAP7_75t_L g8810 ( 
.A(n_8414),
.B(n_6107),
.Y(n_8810)
);

BUFx2_ASAP7_75t_L g8811 ( 
.A(n_8111),
.Y(n_8811)
);

BUFx6f_ASAP7_75t_L g8812 ( 
.A(n_8083),
.Y(n_8812)
);

INVx2_ASAP7_75t_L g8813 ( 
.A(n_8086),
.Y(n_8813)
);

INVx2_ASAP7_75t_L g8814 ( 
.A(n_8088),
.Y(n_8814)
);

AND2x2_ASAP7_75t_L g8815 ( 
.A(n_8362),
.B(n_8350),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_8216),
.Y(n_8816)
);

OAI21x1_ASAP7_75t_L g8817 ( 
.A1(n_8217),
.A2(n_6336),
.B(n_6303),
.Y(n_8817)
);

NAND2xp5_ASAP7_75t_L g8818 ( 
.A(n_8032),
.B(n_7265),
.Y(n_8818)
);

AND2x2_ASAP7_75t_L g8819 ( 
.A(n_8353),
.B(n_8354),
.Y(n_8819)
);

AOI22xp5_ASAP7_75t_L g8820 ( 
.A1(n_8415),
.A2(n_6146),
.B1(n_6160),
.B2(n_6127),
.Y(n_8820)
);

HB1xp67_ASAP7_75t_L g8821 ( 
.A(n_8119),
.Y(n_8821)
);

INVxp67_ASAP7_75t_L g8822 ( 
.A(n_8355),
.Y(n_8822)
);

OAI22xp5_ASAP7_75t_L g8823 ( 
.A1(n_8416),
.A2(n_6096),
.B1(n_6097),
.B2(n_6084),
.Y(n_8823)
);

BUFx6f_ASAP7_75t_L g8824 ( 
.A(n_8089),
.Y(n_8824)
);

INVx1_ASAP7_75t_L g8825 ( 
.A(n_8218),
.Y(n_8825)
);

AND2x4_ASAP7_75t_L g8826 ( 
.A(n_8419),
.B(n_7432),
.Y(n_8826)
);

BUFx2_ASAP7_75t_L g8827 ( 
.A(n_8173),
.Y(n_8827)
);

INVx1_ASAP7_75t_L g8828 ( 
.A(n_8220),
.Y(n_8828)
);

INVx2_ASAP7_75t_L g8829 ( 
.A(n_8091),
.Y(n_8829)
);

CKINVDCx20_ASAP7_75t_R g8830 ( 
.A(n_8163),
.Y(n_8830)
);

AND2x4_ASAP7_75t_L g8831 ( 
.A(n_8423),
.B(n_7463),
.Y(n_8831)
);

CKINVDCx5p33_ASAP7_75t_R g8832 ( 
.A(n_8115),
.Y(n_8832)
);

INVx2_ASAP7_75t_L g8833 ( 
.A(n_8093),
.Y(n_8833)
);

BUFx6f_ASAP7_75t_L g8834 ( 
.A(n_8096),
.Y(n_8834)
);

AOI22x1_ASAP7_75t_SL g8835 ( 
.A1(n_8183),
.A2(n_6521),
.B1(n_6545),
.B2(n_6479),
.Y(n_8835)
);

OA21x2_ASAP7_75t_L g8836 ( 
.A1(n_8224),
.A2(n_6388),
.B(n_6354),
.Y(n_8836)
);

INVx2_ASAP7_75t_L g8837 ( 
.A(n_8099),
.Y(n_8837)
);

NAND2xp5_ASAP7_75t_L g8838 ( 
.A(n_8032),
.B(n_7491),
.Y(n_8838)
);

BUFx2_ASAP7_75t_L g8839 ( 
.A(n_8527),
.Y(n_8839)
);

INVx3_ASAP7_75t_L g8840 ( 
.A(n_8225),
.Y(n_8840)
);

INVx1_ASAP7_75t_L g8841 ( 
.A(n_8227),
.Y(n_8841)
);

CKINVDCx20_ASAP7_75t_R g8842 ( 
.A(n_8189),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_8228),
.Y(n_8843)
);

AND2x4_ASAP7_75t_L g8844 ( 
.A(n_8426),
.B(n_6259),
.Y(n_8844)
);

INVx5_ASAP7_75t_L g8845 ( 
.A(n_8346),
.Y(n_8845)
);

AOI22xp5_ASAP7_75t_L g8846 ( 
.A1(n_8428),
.A2(n_6237),
.B1(n_6254),
.B2(n_6166),
.Y(n_8846)
);

AND2x4_ASAP7_75t_L g8847 ( 
.A(n_8433),
.B(n_6260),
.Y(n_8847)
);

INVx2_ASAP7_75t_L g8848 ( 
.A(n_8103),
.Y(n_8848)
);

INVx3_ASAP7_75t_L g8849 ( 
.A(n_8229),
.Y(n_8849)
);

BUFx6f_ASAP7_75t_L g8850 ( 
.A(n_8105),
.Y(n_8850)
);

INVx2_ASAP7_75t_L g8851 ( 
.A(n_8106),
.Y(n_8851)
);

AND2x4_ASAP7_75t_L g8852 ( 
.A(n_8436),
.B(n_6261),
.Y(n_8852)
);

INVxp33_ASAP7_75t_SL g8853 ( 
.A(n_8139),
.Y(n_8853)
);

INVx3_ASAP7_75t_L g8854 ( 
.A(n_8230),
.Y(n_8854)
);

BUFx2_ASAP7_75t_L g8855 ( 
.A(n_8214),
.Y(n_8855)
);

BUFx12f_ASAP7_75t_L g8856 ( 
.A(n_8146),
.Y(n_8856)
);

BUFx6f_ASAP7_75t_L g8857 ( 
.A(n_8107),
.Y(n_8857)
);

BUFx6f_ASAP7_75t_L g8858 ( 
.A(n_8108),
.Y(n_8858)
);

AOI22xp5_ASAP7_75t_L g8859 ( 
.A1(n_8437),
.A2(n_8447),
.B1(n_8451),
.B2(n_8440),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_8232),
.Y(n_8860)
);

AND2x4_ASAP7_75t_L g8861 ( 
.A(n_8457),
.B(n_6266),
.Y(n_8861)
);

INVx1_ASAP7_75t_L g8862 ( 
.A(n_8236),
.Y(n_8862)
);

INVx2_ASAP7_75t_L g8863 ( 
.A(n_8109),
.Y(n_8863)
);

INVx2_ASAP7_75t_L g8864 ( 
.A(n_8110),
.Y(n_8864)
);

AND2x6_ASAP7_75t_L g8865 ( 
.A(n_8459),
.B(n_8460),
.Y(n_8865)
);

NOR2xp33_ASAP7_75t_L g8866 ( 
.A(n_8461),
.B(n_8462),
.Y(n_8866)
);

OA21x2_ASAP7_75t_L g8867 ( 
.A1(n_8312),
.A2(n_6430),
.B(n_6411),
.Y(n_8867)
);

BUFx8_ASAP7_75t_SL g8868 ( 
.A(n_8192),
.Y(n_8868)
);

AND2x6_ASAP7_75t_L g8869 ( 
.A(n_8465),
.B(n_6397),
.Y(n_8869)
);

OAI21x1_ASAP7_75t_L g8870 ( 
.A1(n_8315),
.A2(n_6494),
.B(n_6464),
.Y(n_8870)
);

HB1xp67_ASAP7_75t_L g8871 ( 
.A(n_8171),
.Y(n_8871)
);

OA21x2_ASAP7_75t_L g8872 ( 
.A1(n_8316),
.A2(n_6509),
.B(n_6496),
.Y(n_8872)
);

CKINVDCx6p67_ASAP7_75t_R g8873 ( 
.A(n_8482),
.Y(n_8873)
);

NAND2xp5_ASAP7_75t_L g8874 ( 
.A(n_8032),
.B(n_6513),
.Y(n_8874)
);

INVx1_ASAP7_75t_L g8875 ( 
.A(n_8317),
.Y(n_8875)
);

BUFx6f_ASAP7_75t_L g8876 ( 
.A(n_8112),
.Y(n_8876)
);

NAND2xp5_ASAP7_75t_L g8877 ( 
.A(n_8032),
.B(n_8318),
.Y(n_8877)
);

INVx2_ASAP7_75t_L g8878 ( 
.A(n_8113),
.Y(n_8878)
);

INVx4_ASAP7_75t_L g8879 ( 
.A(n_8148),
.Y(n_8879)
);

INVx2_ASAP7_75t_L g8880 ( 
.A(n_8117),
.Y(n_8880)
);

AND2x2_ASAP7_75t_L g8881 ( 
.A(n_8357),
.B(n_6595),
.Y(n_8881)
);

NAND2xp5_ASAP7_75t_L g8882 ( 
.A(n_8032),
.B(n_6514),
.Y(n_8882)
);

INVx3_ASAP7_75t_L g8883 ( 
.A(n_8322),
.Y(n_8883)
);

INVx5_ASAP7_75t_L g8884 ( 
.A(n_8323),
.Y(n_8884)
);

BUFx2_ASAP7_75t_L g8885 ( 
.A(n_8320),
.Y(n_8885)
);

INVx2_ASAP7_75t_L g8886 ( 
.A(n_8118),
.Y(n_8886)
);

INVx2_ASAP7_75t_L g8887 ( 
.A(n_8120),
.Y(n_8887)
);

INVx1_ASAP7_75t_L g8888 ( 
.A(n_8324),
.Y(n_8888)
);

AND2x4_ASAP7_75t_L g8889 ( 
.A(n_8466),
.B(n_6271),
.Y(n_8889)
);

BUFx6f_ASAP7_75t_L g8890 ( 
.A(n_8121),
.Y(n_8890)
);

BUFx2_ASAP7_75t_L g8891 ( 
.A(n_8453),
.Y(n_8891)
);

BUFx6f_ASAP7_75t_L g8892 ( 
.A(n_8325),
.Y(n_8892)
);

BUFx6f_ASAP7_75t_L g8893 ( 
.A(n_8016),
.Y(n_8893)
);

BUFx6f_ASAP7_75t_L g8894 ( 
.A(n_8018),
.Y(n_8894)
);

INVx4_ASAP7_75t_L g8895 ( 
.A(n_8159),
.Y(n_8895)
);

BUFx6f_ASAP7_75t_L g8896 ( 
.A(n_8520),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8522),
.Y(n_8897)
);

INVx2_ASAP7_75t_L g8898 ( 
.A(n_8523),
.Y(n_8898)
);

INVx2_ASAP7_75t_L g8899 ( 
.A(n_8524),
.Y(n_8899)
);

INVx2_ASAP7_75t_L g8900 ( 
.A(n_8526),
.Y(n_8900)
);

INVx1_ASAP7_75t_L g8901 ( 
.A(n_8528),
.Y(n_8901)
);

INVx5_ASAP7_75t_L g8902 ( 
.A(n_8483),
.Y(n_8902)
);

HB1xp67_ASAP7_75t_L g8903 ( 
.A(n_8244),
.Y(n_8903)
);

INVx2_ASAP7_75t_L g8904 ( 
.A(n_8530),
.Y(n_8904)
);

INVx2_ASAP7_75t_L g8905 ( 
.A(n_8533),
.Y(n_8905)
);

INVx1_ASAP7_75t_L g8906 ( 
.A(n_8536),
.Y(n_8906)
);

INVx1_ASAP7_75t_L g8907 ( 
.A(n_8537),
.Y(n_8907)
);

INVx3_ASAP7_75t_L g8908 ( 
.A(n_8538),
.Y(n_8908)
);

BUFx6f_ASAP7_75t_L g8909 ( 
.A(n_8541),
.Y(n_8909)
);

CKINVDCx5p33_ASAP7_75t_R g8910 ( 
.A(n_8167),
.Y(n_8910)
);

INVx3_ASAP7_75t_L g8911 ( 
.A(n_8542),
.Y(n_8911)
);

INVx2_ASAP7_75t_L g8912 ( 
.A(n_8545),
.Y(n_8912)
);

HB1xp67_ASAP7_75t_L g8913 ( 
.A(n_8458),
.Y(n_8913)
);

CKINVDCx20_ASAP7_75t_R g8914 ( 
.A(n_8195),
.Y(n_8914)
);

BUFx6f_ASAP7_75t_L g8915 ( 
.A(n_8546),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_L g8916 ( 
.A(n_8521),
.B(n_8467),
.Y(n_8916)
);

INVx5_ASAP7_75t_L g8917 ( 
.A(n_8134),
.Y(n_8917)
);

INVx2_ASAP7_75t_SL g8918 ( 
.A(n_8027),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_8165),
.Y(n_8919)
);

BUFx3_ASAP7_75t_L g8920 ( 
.A(n_8420),
.Y(n_8920)
);

INVx3_ASAP7_75t_L g8921 ( 
.A(n_8358),
.Y(n_8921)
);

HB1xp67_ASAP7_75t_L g8922 ( 
.A(n_8130),
.Y(n_8922)
);

AND2x4_ASAP7_75t_L g8923 ( 
.A(n_8468),
.B(n_6276),
.Y(n_8923)
);

INVx1_ASAP7_75t_L g8924 ( 
.A(n_8170),
.Y(n_8924)
);

CKINVDCx6p67_ASAP7_75t_R g8925 ( 
.A(n_8372),
.Y(n_8925)
);

OAI22xp5_ASAP7_75t_L g8926 ( 
.A1(n_8471),
.A2(n_6099),
.B1(n_6101),
.B2(n_6098),
.Y(n_8926)
);

BUFx6f_ASAP7_75t_L g8927 ( 
.A(n_8360),
.Y(n_8927)
);

CKINVDCx5p33_ASAP7_75t_R g8928 ( 
.A(n_8168),
.Y(n_8928)
);

INVx2_ASAP7_75t_L g8929 ( 
.A(n_8361),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_8174),
.Y(n_8930)
);

INVx2_ASAP7_75t_L g8931 ( 
.A(n_8364),
.Y(n_8931)
);

INVx2_ASAP7_75t_SL g8932 ( 
.A(n_8157),
.Y(n_8932)
);

INVx2_ASAP7_75t_L g8933 ( 
.A(n_8366),
.Y(n_8933)
);

NOR2xp33_ASAP7_75t_L g8934 ( 
.A(n_8476),
.B(n_8477),
.Y(n_8934)
);

INVx3_ASAP7_75t_L g8935 ( 
.A(n_8368),
.Y(n_8935)
);

INVx3_ASAP7_75t_L g8936 ( 
.A(n_8478),
.Y(n_8936)
);

CKINVDCx5p33_ASAP7_75t_R g8937 ( 
.A(n_8179),
.Y(n_8937)
);

AND2x4_ASAP7_75t_L g8938 ( 
.A(n_8479),
.B(n_8480),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_8176),
.Y(n_8939)
);

INVx2_ASAP7_75t_L g8940 ( 
.A(n_8186),
.Y(n_8940)
);

BUFx6f_ASAP7_75t_L g8941 ( 
.A(n_8481),
.Y(n_8941)
);

CKINVDCx20_ASAP7_75t_R g8942 ( 
.A(n_8221),
.Y(n_8942)
);

INVx1_ASAP7_75t_L g8943 ( 
.A(n_8196),
.Y(n_8943)
);

INVx1_ASAP7_75t_L g8944 ( 
.A(n_8208),
.Y(n_8944)
);

BUFx2_ASAP7_75t_L g8945 ( 
.A(n_8473),
.Y(n_8945)
);

OAI22x1_ASAP7_75t_SL g8946 ( 
.A1(n_8246),
.A2(n_6580),
.B1(n_6584),
.B2(n_6551),
.Y(n_8946)
);

INVx2_ASAP7_75t_L g8947 ( 
.A(n_8211),
.Y(n_8947)
);

OAI22x1_ASAP7_75t_SL g8948 ( 
.A1(n_8255),
.A2(n_6653),
.B1(n_6656),
.B2(n_6599),
.Y(n_8948)
);

INVx2_ASAP7_75t_L g8949 ( 
.A(n_8226),
.Y(n_8949)
);

INVx2_ASAP7_75t_L g8950 ( 
.A(n_8234),
.Y(n_8950)
);

INVx2_ASAP7_75t_L g8951 ( 
.A(n_8242),
.Y(n_8951)
);

INVx1_ASAP7_75t_L g8952 ( 
.A(n_8248),
.Y(n_8952)
);

INVx1_ASAP7_75t_L g8953 ( 
.A(n_8251),
.Y(n_8953)
);

AOI22xp5_ASAP7_75t_L g8954 ( 
.A1(n_8484),
.A2(n_6431),
.B1(n_6439),
.B2(n_6414),
.Y(n_8954)
);

AND2x4_ASAP7_75t_L g8955 ( 
.A(n_8486),
.B(n_6277),
.Y(n_8955)
);

OAI22x1_ASAP7_75t_SL g8956 ( 
.A1(n_8256),
.A2(n_6702),
.B1(n_6734),
.B2(n_6659),
.Y(n_8956)
);

AND2x4_ASAP7_75t_L g8957 ( 
.A(n_8487),
.B(n_8492),
.Y(n_8957)
);

BUFx6f_ASAP7_75t_L g8958 ( 
.A(n_8494),
.Y(n_8958)
);

BUFx3_ASAP7_75t_L g8959 ( 
.A(n_8427),
.Y(n_8959)
);

INVx3_ASAP7_75t_L g8960 ( 
.A(n_8498),
.Y(n_8960)
);

BUFx12f_ASAP7_75t_L g8961 ( 
.A(n_8185),
.Y(n_8961)
);

BUFx6f_ASAP7_75t_L g8962 ( 
.A(n_8500),
.Y(n_8962)
);

BUFx8_ASAP7_75t_SL g8963 ( 
.A(n_8337),
.Y(n_8963)
);

BUFx6f_ASAP7_75t_L g8964 ( 
.A(n_8501),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_8259),
.Y(n_8965)
);

AND2x2_ASAP7_75t_L g8966 ( 
.A(n_8514),
.B(n_6595),
.Y(n_8966)
);

BUFx12f_ASAP7_75t_L g8967 ( 
.A(n_8191),
.Y(n_8967)
);

NAND2xp5_ASAP7_75t_L g8968 ( 
.A(n_8504),
.B(n_6550),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_L g8969 ( 
.A(n_8505),
.B(n_6553),
.Y(n_8969)
);

NOR2x1_ASAP7_75t_L g8970 ( 
.A(n_8510),
.B(n_6561),
.Y(n_8970)
);

INVx2_ASAP7_75t_L g8971 ( 
.A(n_8271),
.Y(n_8971)
);

INVx3_ASAP7_75t_L g8972 ( 
.A(n_8512),
.Y(n_8972)
);

HB1xp67_ASAP7_75t_L g8973 ( 
.A(n_8184),
.Y(n_8973)
);

BUFx12f_ASAP7_75t_L g8974 ( 
.A(n_8201),
.Y(n_8974)
);

OAI21x1_ASAP7_75t_L g8975 ( 
.A1(n_8517),
.A2(n_6641),
.B(n_6627),
.Y(n_8975)
);

INVx2_ASAP7_75t_SL g8976 ( 
.A(n_8446),
.Y(n_8976)
);

OAI21x1_ASAP7_75t_L g8977 ( 
.A1(n_8518),
.A2(n_6697),
.B(n_6648),
.Y(n_8977)
);

AOI22xp5_ASAP7_75t_L g8978 ( 
.A1(n_8519),
.A2(n_6598),
.B1(n_6665),
.B2(n_6507),
.Y(n_8978)
);

CKINVDCx5p33_ASAP7_75t_R g8979 ( 
.A(n_8212),
.Y(n_8979)
);

AOI22xp5_ASAP7_75t_L g8980 ( 
.A1(n_8301),
.A2(n_6856),
.B1(n_6899),
.B2(n_6794),
.Y(n_8980)
);

INVx2_ASAP7_75t_L g8981 ( 
.A(n_8296),
.Y(n_8981)
);

CKINVDCx16_ASAP7_75t_R g8982 ( 
.A(n_8397),
.Y(n_8982)
);

AND2x2_ASAP7_75t_L g8983 ( 
.A(n_8532),
.B(n_6620),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_8449),
.Y(n_8984)
);

OA21x2_ASAP7_75t_L g8985 ( 
.A1(n_8491),
.A2(n_6808),
.B(n_6800),
.Y(n_8985)
);

INVx2_ASAP7_75t_L g8986 ( 
.A(n_8513),
.Y(n_8986)
);

BUFx2_ASAP7_75t_L g8987 ( 
.A(n_8493),
.Y(n_8987)
);

INVx4_ASAP7_75t_L g8988 ( 
.A(n_8223),
.Y(n_8988)
);

INVx2_ASAP7_75t_L g8989 ( 
.A(n_8455),
.Y(n_8989)
);

INVx2_ASAP7_75t_L g8990 ( 
.A(n_8489),
.Y(n_8990)
);

AOI22xp5_ASAP7_75t_L g8991 ( 
.A1(n_8308),
.A2(n_8395),
.B1(n_8356),
.B2(n_8231),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_8508),
.Y(n_8992)
);

NOR2xp33_ASAP7_75t_L g8993 ( 
.A(n_8258),
.B(n_6106),
.Y(n_8993)
);

INVx2_ASAP7_75t_L g8994 ( 
.A(n_8260),
.Y(n_8994)
);

INVx6_ASAP7_75t_L g8995 ( 
.A(n_8043),
.Y(n_8995)
);

INVx2_ASAP7_75t_L g8996 ( 
.A(n_8261),
.Y(n_8996)
);

INVx5_ASAP7_75t_L g8997 ( 
.A(n_8072),
.Y(n_8997)
);

CKINVDCx5p33_ASAP7_75t_R g8998 ( 
.A(n_8268),
.Y(n_8998)
);

INVx2_ASAP7_75t_L g8999 ( 
.A(n_8279),
.Y(n_8999)
);

NOR2xp33_ASAP7_75t_L g9000 ( 
.A(n_8280),
.B(n_6109),
.Y(n_9000)
);

OA21x2_ASAP7_75t_L g9001 ( 
.A1(n_8283),
.A2(n_6861),
.B(n_6825),
.Y(n_9001)
);

INVx1_ASAP7_75t_L g9002 ( 
.A(n_8290),
.Y(n_9002)
);

AND2x4_ASAP7_75t_L g9003 ( 
.A(n_8497),
.B(n_8444),
.Y(n_9003)
);

OAI22xp5_ASAP7_75t_SL g9004 ( 
.A1(n_8441),
.A2(n_6769),
.B1(n_6778),
.B2(n_6750),
.Y(n_9004)
);

AND2x4_ASAP7_75t_L g9005 ( 
.A(n_8295),
.B(n_6278),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8297),
.Y(n_9006)
);

INVx1_ASAP7_75t_L g9007 ( 
.A(n_8302),
.Y(n_9007)
);

BUFx6f_ASAP7_75t_L g9008 ( 
.A(n_8306),
.Y(n_9008)
);

INVx1_ASAP7_75t_L g9009 ( 
.A(n_8309),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8311),
.Y(n_9010)
);

INVx4_ASAP7_75t_L g9011 ( 
.A(n_8319),
.Y(n_9011)
);

CKINVDCx16_ASAP7_75t_R g9012 ( 
.A(n_8405),
.Y(n_9012)
);

INVx1_ASAP7_75t_L g9013 ( 
.A(n_8321),
.Y(n_9013)
);

NAND2xp5_ASAP7_75t_L g9014 ( 
.A(n_8331),
.B(n_6864),
.Y(n_9014)
);

BUFx2_ASAP7_75t_L g9015 ( 
.A(n_8445),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_8339),
.Y(n_9016)
);

INVx3_ASAP7_75t_L g9017 ( 
.A(n_8351),
.Y(n_9017)
);

BUFx2_ASAP7_75t_L g9018 ( 
.A(n_8463),
.Y(n_9018)
);

BUFx12f_ASAP7_75t_L g9019 ( 
.A(n_8352),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_8359),
.Y(n_9020)
);

INVx1_ASAP7_75t_L g9021 ( 
.A(n_8369),
.Y(n_9021)
);

AND2x2_ASAP7_75t_L g9022 ( 
.A(n_8448),
.B(n_6620),
.Y(n_9022)
);

INVx1_ASAP7_75t_L g9023 ( 
.A(n_8374),
.Y(n_9023)
);

BUFx6f_ASAP7_75t_L g9024 ( 
.A(n_8377),
.Y(n_9024)
);

INVx2_ASAP7_75t_L g9025 ( 
.A(n_8382),
.Y(n_9025)
);

BUFx6f_ASAP7_75t_L g9026 ( 
.A(n_8391),
.Y(n_9026)
);

INVx2_ASAP7_75t_L g9027 ( 
.A(n_8393),
.Y(n_9027)
);

INVx2_ASAP7_75t_L g9028 ( 
.A(n_8399),
.Y(n_9028)
);

BUFx6f_ASAP7_75t_L g9029 ( 
.A(n_8401),
.Y(n_9029)
);

BUFx2_ASAP7_75t_L g9030 ( 
.A(n_8470),
.Y(n_9030)
);

AOI22x1_ASAP7_75t_SL g9031 ( 
.A1(n_8539),
.A2(n_6801),
.B1(n_6817),
.B2(n_6787),
.Y(n_9031)
);

NAND2xp5_ASAP7_75t_L g9032 ( 
.A(n_8403),
.B(n_6915),
.Y(n_9032)
);

INVx6_ASAP7_75t_L g9033 ( 
.A(n_8080),
.Y(n_9033)
);

BUFx3_ASAP7_75t_L g9034 ( 
.A(n_8495),
.Y(n_9034)
);

INVx1_ASAP7_75t_L g9035 ( 
.A(n_8409),
.Y(n_9035)
);

AOI22xp5_ASAP7_75t_L g9036 ( 
.A1(n_8424),
.A2(n_7012),
.B1(n_7027),
.B2(n_7008),
.Y(n_9036)
);

INVx3_ASAP7_75t_L g9037 ( 
.A(n_8429),
.Y(n_9037)
);

INVx1_ASAP7_75t_L g9038 ( 
.A(n_8431),
.Y(n_9038)
);

INVx4_ASAP7_75t_L g9039 ( 
.A(n_8432),
.Y(n_9039)
);

INVx1_ASAP7_75t_L g9040 ( 
.A(n_8434),
.Y(n_9040)
);

BUFx6f_ASAP7_75t_L g9041 ( 
.A(n_8435),
.Y(n_9041)
);

INVx6_ASAP7_75t_L g9042 ( 
.A(n_8097),
.Y(n_9042)
);

BUFx6f_ASAP7_75t_L g9043 ( 
.A(n_8442),
.Y(n_9043)
);

INVx2_ASAP7_75t_L g9044 ( 
.A(n_8443),
.Y(n_9044)
);

AOI22xp5_ASAP7_75t_L g9045 ( 
.A1(n_8450),
.A2(n_8454),
.B1(n_8464),
.B2(n_8452),
.Y(n_9045)
);

BUFx6f_ASAP7_75t_L g9046 ( 
.A(n_8472),
.Y(n_9046)
);

INVx2_ASAP7_75t_L g9047 ( 
.A(n_8475),
.Y(n_9047)
);

INVx2_ASAP7_75t_SL g9048 ( 
.A(n_8488),
.Y(n_9048)
);

OAI21x1_ASAP7_75t_L g9049 ( 
.A1(n_8490),
.A2(n_6953),
.B(n_6937),
.Y(n_9049)
);

CKINVDCx20_ASAP7_75t_R g9050 ( 
.A(n_8496),
.Y(n_9050)
);

INVx6_ASAP7_75t_L g9051 ( 
.A(n_8135),
.Y(n_9051)
);

CKINVDCx6p67_ASAP7_75t_R g9052 ( 
.A(n_8506),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_8502),
.Y(n_9053)
);

INVx2_ASAP7_75t_L g9054 ( 
.A(n_8503),
.Y(n_9054)
);

INVx1_ASAP7_75t_L g9055 ( 
.A(n_8516),
.Y(n_9055)
);

OAI22xp5_ASAP7_75t_L g9056 ( 
.A1(n_8540),
.A2(n_6114),
.B1(n_6118),
.B2(n_6111),
.Y(n_9056)
);

INVx2_ASAP7_75t_L g9057 ( 
.A(n_8515),
.Y(n_9057)
);

INVx2_ASAP7_75t_L g9058 ( 
.A(n_8166),
.Y(n_9058)
);

INVx1_ASAP7_75t_L g9059 ( 
.A(n_8040),
.Y(n_9059)
);

AND2x2_ASAP7_75t_L g9060 ( 
.A(n_8507),
.B(n_6629),
.Y(n_9060)
);

NAND2xp33_ASAP7_75t_L g9061 ( 
.A(n_8365),
.B(n_6655),
.Y(n_9061)
);

INVx5_ASAP7_75t_L g9062 ( 
.A(n_8235),
.Y(n_9062)
);

AND2x2_ASAP7_75t_L g9063 ( 
.A(n_8375),
.B(n_6629),
.Y(n_9063)
);

CKINVDCx5p33_ASAP7_75t_R g9064 ( 
.A(n_8190),
.Y(n_9064)
);

HB1xp67_ASAP7_75t_L g9065 ( 
.A(n_8215),
.Y(n_9065)
);

BUFx3_ASAP7_75t_L g9066 ( 
.A(n_8078),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8238),
.Y(n_9067)
);

OAI21x1_ASAP7_75t_L g9068 ( 
.A1(n_8326),
.A2(n_6965),
.B(n_6956),
.Y(n_9068)
);

INVx3_ASAP7_75t_L g9069 ( 
.A(n_8078),
.Y(n_9069)
);

XNOR2xp5_ASAP7_75t_L g9070 ( 
.A(n_8063),
.B(n_6818),
.Y(n_9070)
);

CKINVDCx5p33_ASAP7_75t_R g9071 ( 
.A(n_8017),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_8238),
.Y(n_9072)
);

INVx1_ASAP7_75t_L g9073 ( 
.A(n_8238),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_8238),
.Y(n_9074)
);

INVx1_ASAP7_75t_L g9075 ( 
.A(n_8238),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_8238),
.Y(n_9076)
);

BUFx2_ASAP7_75t_L g9077 ( 
.A(n_8425),
.Y(n_9077)
);

INVx2_ASAP7_75t_L g9078 ( 
.A(n_8153),
.Y(n_9078)
);

HB1xp67_ASAP7_75t_L g9079 ( 
.A(n_8425),
.Y(n_9079)
);

AND2x4_ASAP7_75t_L g9080 ( 
.A(n_8237),
.B(n_6281),
.Y(n_9080)
);

OAI21x1_ASAP7_75t_L g9081 ( 
.A1(n_8326),
.A2(n_7025),
.B(n_6990),
.Y(n_9081)
);

BUFx6f_ASAP7_75t_L g9082 ( 
.A(n_8044),
.Y(n_9082)
);

OA21x2_ASAP7_75t_L g9083 ( 
.A1(n_8326),
.A2(n_7029),
.B(n_7028),
.Y(n_9083)
);

BUFx12f_ASAP7_75t_L g9084 ( 
.A(n_8017),
.Y(n_9084)
);

AND2x4_ASAP7_75t_L g9085 ( 
.A(n_8237),
.B(n_6288),
.Y(n_9085)
);

BUFx8_ASAP7_75t_SL g9086 ( 
.A(n_8063),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_8238),
.Y(n_9087)
);

BUFx6f_ASAP7_75t_L g9088 ( 
.A(n_8044),
.Y(n_9088)
);

INVxp67_ASAP7_75t_L g9089 ( 
.A(n_8392),
.Y(n_9089)
);

INVx5_ASAP7_75t_L g9090 ( 
.A(n_8485),
.Y(n_9090)
);

HB1xp67_ASAP7_75t_L g9091 ( 
.A(n_8425),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_8238),
.Y(n_9092)
);

BUFx8_ASAP7_75t_L g9093 ( 
.A(n_8485),
.Y(n_9093)
);

OAI21x1_ASAP7_75t_L g9094 ( 
.A1(n_8326),
.A2(n_7160),
.B(n_7158),
.Y(n_9094)
);

BUFx6f_ASAP7_75t_L g9095 ( 
.A(n_8044),
.Y(n_9095)
);

INVx2_ASAP7_75t_L g9096 ( 
.A(n_8153),
.Y(n_9096)
);

HB1xp67_ASAP7_75t_L g9097 ( 
.A(n_8425),
.Y(n_9097)
);

BUFx3_ASAP7_75t_L g9098 ( 
.A(n_8078),
.Y(n_9098)
);

BUFx6f_ASAP7_75t_L g9099 ( 
.A(n_8044),
.Y(n_9099)
);

OA21x2_ASAP7_75t_L g9100 ( 
.A1(n_8326),
.A2(n_7162),
.B(n_7161),
.Y(n_9100)
);

BUFx12f_ASAP7_75t_L g9101 ( 
.A(n_8017),
.Y(n_9101)
);

OAI21x1_ASAP7_75t_L g9102 ( 
.A1(n_8326),
.A2(n_7234),
.B(n_7191),
.Y(n_9102)
);

AND2x2_ASAP7_75t_L g9103 ( 
.A(n_8430),
.B(n_6696),
.Y(n_9103)
);

CKINVDCx16_ASAP7_75t_R g9104 ( 
.A(n_8075),
.Y(n_9104)
);

BUFx6f_ASAP7_75t_L g9105 ( 
.A(n_8044),
.Y(n_9105)
);

AND2x2_ASAP7_75t_L g9106 ( 
.A(n_8430),
.B(n_6696),
.Y(n_9106)
);

INVx2_ASAP7_75t_L g9107 ( 
.A(n_8153),
.Y(n_9107)
);

INVx3_ASAP7_75t_L g9108 ( 
.A(n_8078),
.Y(n_9108)
);

INVx2_ASAP7_75t_L g9109 ( 
.A(n_8153),
.Y(n_9109)
);

BUFx6f_ASAP7_75t_L g9110 ( 
.A(n_8044),
.Y(n_9110)
);

NAND2xp5_ASAP7_75t_L g9111 ( 
.A(n_8162),
.B(n_7245),
.Y(n_9111)
);

HB1xp67_ASAP7_75t_L g9112 ( 
.A(n_8425),
.Y(n_9112)
);

BUFx2_ASAP7_75t_L g9113 ( 
.A(n_8425),
.Y(n_9113)
);

INVx3_ASAP7_75t_L g9114 ( 
.A(n_8078),
.Y(n_9114)
);

INVxp67_ASAP7_75t_L g9115 ( 
.A(n_8392),
.Y(n_9115)
);

CKINVDCx20_ASAP7_75t_R g9116 ( 
.A(n_8063),
.Y(n_9116)
);

NAND2x1_ASAP7_75t_L g9117 ( 
.A(n_8151),
.B(n_6537),
.Y(n_9117)
);

BUFx6f_ASAP7_75t_L g9118 ( 
.A(n_8044),
.Y(n_9118)
);

CKINVDCx5p33_ASAP7_75t_R g9119 ( 
.A(n_8017),
.Y(n_9119)
);

BUFx2_ASAP7_75t_L g9120 ( 
.A(n_8425),
.Y(n_9120)
);

BUFx6f_ASAP7_75t_L g9121 ( 
.A(n_8044),
.Y(n_9121)
);

XNOR2x2_ASAP7_75t_L g9122 ( 
.A(n_8199),
.B(n_7477),
.Y(n_9122)
);

AOI22xp5_ASAP7_75t_L g9123 ( 
.A1(n_8156),
.A2(n_7045),
.B1(n_7063),
.B2(n_7043),
.Y(n_9123)
);

BUFx3_ASAP7_75t_L g9124 ( 
.A(n_8078),
.Y(n_9124)
);

BUFx8_ASAP7_75t_L g9125 ( 
.A(n_8485),
.Y(n_9125)
);

BUFx6f_ASAP7_75t_L g9126 ( 
.A(n_8044),
.Y(n_9126)
);

INVx2_ASAP7_75t_L g9127 ( 
.A(n_8153),
.Y(n_9127)
);

INVx2_ASAP7_75t_L g9128 ( 
.A(n_8153),
.Y(n_9128)
);

CKINVDCx6p67_ASAP7_75t_R g9129 ( 
.A(n_8387),
.Y(n_9129)
);

CKINVDCx5p33_ASAP7_75t_R g9130 ( 
.A(n_8017),
.Y(n_9130)
);

AND2x6_ASAP7_75t_L g9131 ( 
.A(n_8383),
.B(n_7093),
.Y(n_9131)
);

BUFx6f_ASAP7_75t_L g9132 ( 
.A(n_8044),
.Y(n_9132)
);

INVx3_ASAP7_75t_L g9133 ( 
.A(n_8571),
.Y(n_9133)
);

AND2x2_ASAP7_75t_L g9134 ( 
.A(n_8630),
.B(n_8573),
.Y(n_9134)
);

INVx1_ASAP7_75t_L g9135 ( 
.A(n_8551),
.Y(n_9135)
);

INVx2_ASAP7_75t_L g9136 ( 
.A(n_8594),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_8564),
.Y(n_9137)
);

CKINVDCx5p33_ASAP7_75t_R g9138 ( 
.A(n_8868),
.Y(n_9138)
);

INVx1_ASAP7_75t_L g9139 ( 
.A(n_8565),
.Y(n_9139)
);

AND2x4_ASAP7_75t_L g9140 ( 
.A(n_9066),
.B(n_6292),
.Y(n_9140)
);

INVxp67_ASAP7_75t_SL g9141 ( 
.A(n_8666),
.Y(n_9141)
);

NAND2xp5_ASAP7_75t_L g9142 ( 
.A(n_8783),
.B(n_7267),
.Y(n_9142)
);

CKINVDCx5p33_ASAP7_75t_R g9143 ( 
.A(n_8963),
.Y(n_9143)
);

CKINVDCx5p33_ASAP7_75t_R g9144 ( 
.A(n_9086),
.Y(n_9144)
);

NAND2xp5_ASAP7_75t_SL g9145 ( 
.A(n_8641),
.B(n_6655),
.Y(n_9145)
);

INVx1_ASAP7_75t_L g9146 ( 
.A(n_8569),
.Y(n_9146)
);

BUFx6f_ASAP7_75t_L g9147 ( 
.A(n_9098),
.Y(n_9147)
);

INVx3_ASAP7_75t_L g9148 ( 
.A(n_8574),
.Y(n_9148)
);

BUFx6f_ASAP7_75t_L g9149 ( 
.A(n_9124),
.Y(n_9149)
);

CKINVDCx5p33_ASAP7_75t_R g9150 ( 
.A(n_9130),
.Y(n_9150)
);

BUFx6f_ASAP7_75t_L g9151 ( 
.A(n_8555),
.Y(n_9151)
);

AND2x2_ASAP7_75t_L g9152 ( 
.A(n_8602),
.B(n_6737),
.Y(n_9152)
);

CKINVDCx5p33_ASAP7_75t_R g9153 ( 
.A(n_8549),
.Y(n_9153)
);

AND2x6_ASAP7_75t_L g9154 ( 
.A(n_8936),
.B(n_7270),
.Y(n_9154)
);

NAND2xp5_ASAP7_75t_L g9155 ( 
.A(n_8656),
.B(n_7315),
.Y(n_9155)
);

INVx1_ASAP7_75t_L g9156 ( 
.A(n_8570),
.Y(n_9156)
);

AND2x6_ASAP7_75t_L g9157 ( 
.A(n_8960),
.B(n_7337),
.Y(n_9157)
);

CKINVDCx5p33_ASAP7_75t_R g9158 ( 
.A(n_9119),
.Y(n_9158)
);

INVx2_ASAP7_75t_L g9159 ( 
.A(n_8600),
.Y(n_9159)
);

INVx1_ASAP7_75t_L g9160 ( 
.A(n_8577),
.Y(n_9160)
);

BUFx3_ASAP7_75t_L g9161 ( 
.A(n_8585),
.Y(n_9161)
);

NAND2xp5_ASAP7_75t_SL g9162 ( 
.A(n_8706),
.B(n_6688),
.Y(n_9162)
);

NOR2xp33_ASAP7_75t_L g9163 ( 
.A(n_9089),
.B(n_7135),
.Y(n_9163)
);

INVx2_ASAP7_75t_L g9164 ( 
.A(n_8601),
.Y(n_9164)
);

CKINVDCx5p33_ASAP7_75t_R g9165 ( 
.A(n_8621),
.Y(n_9165)
);

CKINVDCx20_ASAP7_75t_R g9166 ( 
.A(n_8615),
.Y(n_9166)
);

INVx1_ASAP7_75t_L g9167 ( 
.A(n_8581),
.Y(n_9167)
);

NOR2xp33_ASAP7_75t_L g9168 ( 
.A(n_9115),
.B(n_7197),
.Y(n_9168)
);

BUFx3_ASAP7_75t_L g9169 ( 
.A(n_8587),
.Y(n_9169)
);

INVx2_ASAP7_75t_L g9170 ( 
.A(n_8608),
.Y(n_9170)
);

INVx4_ASAP7_75t_L g9171 ( 
.A(n_9090),
.Y(n_9171)
);

HB1xp67_ASAP7_75t_L g9172 ( 
.A(n_8603),
.Y(n_9172)
);

CKINVDCx20_ASAP7_75t_R g9173 ( 
.A(n_8755),
.Y(n_9173)
);

BUFx6f_ASAP7_75t_L g9174 ( 
.A(n_8561),
.Y(n_9174)
);

BUFx3_ASAP7_75t_L g9175 ( 
.A(n_8781),
.Y(n_9175)
);

BUFx6f_ASAP7_75t_L g9176 ( 
.A(n_8566),
.Y(n_9176)
);

AND2x2_ASAP7_75t_L g9177 ( 
.A(n_9077),
.B(n_6737),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_8583),
.Y(n_9178)
);

INVx1_ASAP7_75t_L g9179 ( 
.A(n_8586),
.Y(n_9179)
);

BUFx6f_ASAP7_75t_L g9180 ( 
.A(n_9082),
.Y(n_9180)
);

CKINVDCx20_ASAP7_75t_R g9181 ( 
.A(n_8830),
.Y(n_9181)
);

CKINVDCx5p33_ASAP7_75t_R g9182 ( 
.A(n_8659),
.Y(n_9182)
);

INVx2_ASAP7_75t_L g9183 ( 
.A(n_8611),
.Y(n_9183)
);

AND2x2_ASAP7_75t_L g9184 ( 
.A(n_9113),
.B(n_6771),
.Y(n_9184)
);

INVx1_ASAP7_75t_L g9185 ( 
.A(n_8595),
.Y(n_9185)
);

INVx1_ASAP7_75t_L g9186 ( 
.A(n_8604),
.Y(n_9186)
);

BUFx6f_ASAP7_75t_L g9187 ( 
.A(n_9088),
.Y(n_9187)
);

BUFx2_ASAP7_75t_L g9188 ( 
.A(n_9120),
.Y(n_9188)
);

NOR2xp33_ASAP7_75t_SL g9189 ( 
.A(n_8853),
.B(n_6887),
.Y(n_9189)
);

INVx1_ASAP7_75t_L g9190 ( 
.A(n_8609),
.Y(n_9190)
);

CKINVDCx5p33_ASAP7_75t_R g9191 ( 
.A(n_8681),
.Y(n_9191)
);

NAND2xp5_ASAP7_75t_L g9192 ( 
.A(n_8940),
.B(n_7346),
.Y(n_9192)
);

INVx2_ASAP7_75t_L g9193 ( 
.A(n_8613),
.Y(n_9193)
);

INVx1_ASAP7_75t_L g9194 ( 
.A(n_8610),
.Y(n_9194)
);

HB1xp67_ASAP7_75t_L g9195 ( 
.A(n_8584),
.Y(n_9195)
);

INVx1_ASAP7_75t_L g9196 ( 
.A(n_8612),
.Y(n_9196)
);

AND2x4_ASAP7_75t_L g9197 ( 
.A(n_8639),
.B(n_6294),
.Y(n_9197)
);

INVx1_ASAP7_75t_L g9198 ( 
.A(n_8622),
.Y(n_9198)
);

CKINVDCx11_ASAP7_75t_R g9199 ( 
.A(n_8873),
.Y(n_9199)
);

INVx2_ASAP7_75t_L g9200 ( 
.A(n_8614),
.Y(n_9200)
);

NAND2xp5_ASAP7_75t_L g9201 ( 
.A(n_8947),
.B(n_7349),
.Y(n_9201)
);

INVx2_ASAP7_75t_L g9202 ( 
.A(n_8620),
.Y(n_9202)
);

INVx1_ASAP7_75t_L g9203 ( 
.A(n_8635),
.Y(n_9203)
);

INVx1_ASAP7_75t_L g9204 ( 
.A(n_8643),
.Y(n_9204)
);

HB1xp67_ASAP7_75t_L g9205 ( 
.A(n_9079),
.Y(n_9205)
);

INVx2_ASAP7_75t_L g9206 ( 
.A(n_8576),
.Y(n_9206)
);

INVx1_ASAP7_75t_L g9207 ( 
.A(n_8646),
.Y(n_9207)
);

INVx1_ASAP7_75t_L g9208 ( 
.A(n_8658),
.Y(n_9208)
);

BUFx6f_ASAP7_75t_L g9209 ( 
.A(n_9095),
.Y(n_9209)
);

BUFx2_ASAP7_75t_L g9210 ( 
.A(n_8871),
.Y(n_9210)
);

CKINVDCx5p33_ASAP7_75t_R g9211 ( 
.A(n_8724),
.Y(n_9211)
);

INVx1_ASAP7_75t_L g9212 ( 
.A(n_8661),
.Y(n_9212)
);

INVx1_ASAP7_75t_L g9213 ( 
.A(n_8662),
.Y(n_9213)
);

HB1xp67_ASAP7_75t_L g9214 ( 
.A(n_9091),
.Y(n_9214)
);

INVx2_ASAP7_75t_L g9215 ( 
.A(n_8592),
.Y(n_9215)
);

CKINVDCx5p33_ASAP7_75t_R g9216 ( 
.A(n_8738),
.Y(n_9216)
);

BUFx2_ASAP7_75t_L g9217 ( 
.A(n_8559),
.Y(n_9217)
);

CKINVDCx5p33_ASAP7_75t_R g9218 ( 
.A(n_8832),
.Y(n_9218)
);

BUFx6f_ASAP7_75t_L g9219 ( 
.A(n_9099),
.Y(n_9219)
);

INVx2_ASAP7_75t_L g9220 ( 
.A(n_8588),
.Y(n_9220)
);

INVx2_ASAP7_75t_L g9221 ( 
.A(n_8898),
.Y(n_9221)
);

NAND2xp5_ASAP7_75t_SL g9222 ( 
.A(n_8558),
.B(n_6688),
.Y(n_9222)
);

BUFx6f_ASAP7_75t_L g9223 ( 
.A(n_9105),
.Y(n_9223)
);

CKINVDCx5p33_ASAP7_75t_R g9224 ( 
.A(n_8910),
.Y(n_9224)
);

INVx1_ASAP7_75t_L g9225 ( 
.A(n_8669),
.Y(n_9225)
);

CKINVDCx5p33_ASAP7_75t_R g9226 ( 
.A(n_8928),
.Y(n_9226)
);

INVx3_ASAP7_75t_L g9227 ( 
.A(n_9069),
.Y(n_9227)
);

INVx2_ASAP7_75t_L g9228 ( 
.A(n_8899),
.Y(n_9228)
);

INVx1_ASAP7_75t_L g9229 ( 
.A(n_8686),
.Y(n_9229)
);

AND2x4_ASAP7_75t_L g9230 ( 
.A(n_8660),
.B(n_6296),
.Y(n_9230)
);

INVx1_ASAP7_75t_L g9231 ( 
.A(n_8688),
.Y(n_9231)
);

INVx1_ASAP7_75t_L g9232 ( 
.A(n_8696),
.Y(n_9232)
);

CKINVDCx20_ASAP7_75t_R g9233 ( 
.A(n_8842),
.Y(n_9233)
);

INVx1_ASAP7_75t_L g9234 ( 
.A(n_8701),
.Y(n_9234)
);

CKINVDCx5p33_ASAP7_75t_R g9235 ( 
.A(n_8937),
.Y(n_9235)
);

INVx2_ASAP7_75t_L g9236 ( 
.A(n_8900),
.Y(n_9236)
);

NAND2xp5_ASAP7_75t_L g9237 ( 
.A(n_8949),
.B(n_7372),
.Y(n_9237)
);

CKINVDCx5p33_ASAP7_75t_R g9238 ( 
.A(n_8979),
.Y(n_9238)
);

CKINVDCx5p33_ASAP7_75t_R g9239 ( 
.A(n_8998),
.Y(n_9239)
);

CKINVDCx5p33_ASAP7_75t_R g9240 ( 
.A(n_9071),
.Y(n_9240)
);

INVx1_ASAP7_75t_L g9241 ( 
.A(n_8704),
.Y(n_9241)
);

INVx1_ASAP7_75t_L g9242 ( 
.A(n_9067),
.Y(n_9242)
);

INVxp67_ASAP7_75t_SL g9243 ( 
.A(n_8619),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_9072),
.Y(n_9244)
);

CKINVDCx5p33_ASAP7_75t_R g9245 ( 
.A(n_8767),
.Y(n_9245)
);

INVx1_ASAP7_75t_L g9246 ( 
.A(n_9073),
.Y(n_9246)
);

BUFx6f_ASAP7_75t_L g9247 ( 
.A(n_9110),
.Y(n_9247)
);

INVx3_ASAP7_75t_L g9248 ( 
.A(n_9108),
.Y(n_9248)
);

NAND2xp5_ASAP7_75t_L g9249 ( 
.A(n_8950),
.B(n_7532),
.Y(n_9249)
);

INVx3_ASAP7_75t_L g9250 ( 
.A(n_9114),
.Y(n_9250)
);

CKINVDCx5p33_ASAP7_75t_R g9251 ( 
.A(n_9064),
.Y(n_9251)
);

NOR2xp33_ASAP7_75t_R g9252 ( 
.A(n_8914),
.B(n_6924),
.Y(n_9252)
);

AND2x2_ASAP7_75t_L g9253 ( 
.A(n_9097),
.B(n_6771),
.Y(n_9253)
);

INVx1_ASAP7_75t_L g9254 ( 
.A(n_9074),
.Y(n_9254)
);

XNOR2x2_ASAP7_75t_L g9255 ( 
.A(n_9122),
.B(n_7273),
.Y(n_9255)
);

CKINVDCx5p33_ASAP7_75t_R g9256 ( 
.A(n_8627),
.Y(n_9256)
);

BUFx2_ASAP7_75t_L g9257 ( 
.A(n_8598),
.Y(n_9257)
);

INVx1_ASAP7_75t_L g9258 ( 
.A(n_9075),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_9076),
.Y(n_9259)
);

BUFx6f_ASAP7_75t_L g9260 ( 
.A(n_9118),
.Y(n_9260)
);

CKINVDCx5p33_ASAP7_75t_R g9261 ( 
.A(n_8671),
.Y(n_9261)
);

AND2x2_ASAP7_75t_L g9262 ( 
.A(n_9112),
.B(n_6839),
.Y(n_9262)
);

OA21x2_ASAP7_75t_L g9263 ( 
.A1(n_8563),
.A2(n_6305),
.B(n_6304),
.Y(n_9263)
);

CKINVDCx5p33_ASAP7_75t_R g9264 ( 
.A(n_8709),
.Y(n_9264)
);

CKINVDCx5p33_ASAP7_75t_R g9265 ( 
.A(n_8712),
.Y(n_9265)
);

NAND2xp5_ASAP7_75t_L g9266 ( 
.A(n_8951),
.B(n_7022),
.Y(n_9266)
);

INVx1_ASAP7_75t_L g9267 ( 
.A(n_9087),
.Y(n_9267)
);

INVx2_ASAP7_75t_L g9268 ( 
.A(n_8904),
.Y(n_9268)
);

INVx2_ASAP7_75t_L g9269 ( 
.A(n_8905),
.Y(n_9269)
);

INVx1_ASAP7_75t_L g9270 ( 
.A(n_9092),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_8929),
.Y(n_9271)
);

INVx1_ASAP7_75t_L g9272 ( 
.A(n_8931),
.Y(n_9272)
);

CKINVDCx5p33_ASAP7_75t_R g9273 ( 
.A(n_8856),
.Y(n_9273)
);

NOR2xp33_ASAP7_75t_R g9274 ( 
.A(n_8942),
.B(n_6926),
.Y(n_9274)
);

AND2x2_ASAP7_75t_L g9275 ( 
.A(n_9103),
.B(n_6839),
.Y(n_9275)
);

CKINVDCx5p33_ASAP7_75t_R g9276 ( 
.A(n_8961),
.Y(n_9276)
);

CKINVDCx5p33_ASAP7_75t_R g9277 ( 
.A(n_8967),
.Y(n_9277)
);

INVx2_ASAP7_75t_L g9278 ( 
.A(n_8912),
.Y(n_9278)
);

NAND2xp5_ASAP7_75t_L g9279 ( 
.A(n_8971),
.B(n_7022),
.Y(n_9279)
);

CKINVDCx5p33_ASAP7_75t_R g9280 ( 
.A(n_8974),
.Y(n_9280)
);

INVx2_ASAP7_75t_L g9281 ( 
.A(n_8875),
.Y(n_9281)
);

INVx1_ASAP7_75t_L g9282 ( 
.A(n_8933),
.Y(n_9282)
);

INVx1_ASAP7_75t_L g9283 ( 
.A(n_8735),
.Y(n_9283)
);

INVx1_ASAP7_75t_L g9284 ( 
.A(n_8740),
.Y(n_9284)
);

CKINVDCx20_ASAP7_75t_R g9285 ( 
.A(n_9116),
.Y(n_9285)
);

CKINVDCx5p33_ASAP7_75t_R g9286 ( 
.A(n_9019),
.Y(n_9286)
);

INVx1_ASAP7_75t_L g9287 ( 
.A(n_8741),
.Y(n_9287)
);

OAI21x1_ASAP7_75t_L g9288 ( 
.A1(n_8667),
.A2(n_6247),
.B(n_6245),
.Y(n_9288)
);

INVxp67_ASAP7_75t_L g9289 ( 
.A(n_8684),
.Y(n_9289)
);

CKINVDCx20_ASAP7_75t_R g9290 ( 
.A(n_9050),
.Y(n_9290)
);

INVx2_ASAP7_75t_L g9291 ( 
.A(n_8888),
.Y(n_9291)
);

INVx1_ASAP7_75t_L g9292 ( 
.A(n_8742),
.Y(n_9292)
);

INVx2_ASAP7_75t_L g9293 ( 
.A(n_8665),
.Y(n_9293)
);

INVx3_ASAP7_75t_L g9294 ( 
.A(n_9121),
.Y(n_9294)
);

INVx3_ASAP7_75t_L g9295 ( 
.A(n_9126),
.Y(n_9295)
);

INVx4_ASAP7_75t_L g9296 ( 
.A(n_8917),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_8748),
.Y(n_9297)
);

INVx1_ASAP7_75t_L g9298 ( 
.A(n_8751),
.Y(n_9298)
);

INVx3_ASAP7_75t_L g9299 ( 
.A(n_9132),
.Y(n_9299)
);

CKINVDCx5p33_ASAP7_75t_R g9300 ( 
.A(n_9084),
.Y(n_9300)
);

CKINVDCx20_ASAP7_75t_R g9301 ( 
.A(n_8982),
.Y(n_9301)
);

INVx1_ASAP7_75t_L g9302 ( 
.A(n_8762),
.Y(n_9302)
);

INVx1_ASAP7_75t_L g9303 ( 
.A(n_8769),
.Y(n_9303)
);

INVx2_ASAP7_75t_L g9304 ( 
.A(n_8670),
.Y(n_9304)
);

INVxp67_ASAP7_75t_L g9305 ( 
.A(n_9106),
.Y(n_9305)
);

INVx1_ASAP7_75t_L g9306 ( 
.A(n_8777),
.Y(n_9306)
);

CKINVDCx5p33_ASAP7_75t_R g9307 ( 
.A(n_9101),
.Y(n_9307)
);

NAND2xp33_ASAP7_75t_R g9308 ( 
.A(n_8676),
.B(n_6135),
.Y(n_9308)
);

BUFx6f_ASAP7_75t_L g9309 ( 
.A(n_8927),
.Y(n_9309)
);

CKINVDCx5p33_ASAP7_75t_R g9310 ( 
.A(n_8925),
.Y(n_9310)
);

NOR2xp33_ASAP7_75t_R g9311 ( 
.A(n_8572),
.B(n_9104),
.Y(n_9311)
);

INVx2_ASAP7_75t_L g9312 ( 
.A(n_8672),
.Y(n_9312)
);

NAND2xp5_ASAP7_75t_L g9313 ( 
.A(n_8981),
.B(n_7495),
.Y(n_9313)
);

HB1xp67_ASAP7_75t_L g9314 ( 
.A(n_8903),
.Y(n_9314)
);

INVx1_ASAP7_75t_L g9315 ( 
.A(n_8780),
.Y(n_9315)
);

INVx2_ASAP7_75t_L g9316 ( 
.A(n_8687),
.Y(n_9316)
);

CKINVDCx5p33_ASAP7_75t_R g9317 ( 
.A(n_9052),
.Y(n_9317)
);

INVx2_ASAP7_75t_L g9318 ( 
.A(n_8689),
.Y(n_9318)
);

INVx1_ASAP7_75t_L g9319 ( 
.A(n_8784),
.Y(n_9319)
);

NOR2xp33_ASAP7_75t_R g9320 ( 
.A(n_9012),
.B(n_6936),
.Y(n_9320)
);

INVx1_ASAP7_75t_L g9321 ( 
.A(n_8787),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_8796),
.Y(n_9322)
);

CKINVDCx5p33_ASAP7_75t_R g9323 ( 
.A(n_9008),
.Y(n_9323)
);

INVx3_ASAP7_75t_L g9324 ( 
.A(n_8562),
.Y(n_9324)
);

NAND2xp5_ASAP7_75t_L g9325 ( 
.A(n_8816),
.B(n_7495),
.Y(n_9325)
);

INVx1_ASAP7_75t_L g9326 ( 
.A(n_8825),
.Y(n_9326)
);

INVx1_ASAP7_75t_L g9327 ( 
.A(n_8828),
.Y(n_9327)
);

INVx1_ASAP7_75t_L g9328 ( 
.A(n_8841),
.Y(n_9328)
);

AND2x2_ASAP7_75t_L g9329 ( 
.A(n_8776),
.B(n_7083),
.Y(n_9329)
);

AND2x2_ASAP7_75t_L g9330 ( 
.A(n_8815),
.B(n_7083),
.Y(n_9330)
);

AND2x2_ASAP7_75t_L g9331 ( 
.A(n_8730),
.B(n_7125),
.Y(n_9331)
);

INVx1_ASAP7_75t_L g9332 ( 
.A(n_8843),
.Y(n_9332)
);

INVx1_ASAP7_75t_L g9333 ( 
.A(n_8860),
.Y(n_9333)
);

INVx1_ASAP7_75t_L g9334 ( 
.A(n_8862),
.Y(n_9334)
);

NAND2xp5_ASAP7_75t_L g9335 ( 
.A(n_8919),
.B(n_7495),
.Y(n_9335)
);

BUFx8_ASAP7_75t_L g9336 ( 
.A(n_9015),
.Y(n_9336)
);

BUFx6f_ASAP7_75t_L g9337 ( 
.A(n_8590),
.Y(n_9337)
);

CKINVDCx5p33_ASAP7_75t_R g9338 ( 
.A(n_9024),
.Y(n_9338)
);

INVx1_ASAP7_75t_L g9339 ( 
.A(n_8897),
.Y(n_9339)
);

AND2x4_ASAP7_75t_L g9340 ( 
.A(n_8567),
.B(n_6310),
.Y(n_9340)
);

NOR2xp33_ASAP7_75t_R g9341 ( 
.A(n_8579),
.B(n_6940),
.Y(n_9341)
);

INVx1_ASAP7_75t_L g9342 ( 
.A(n_8901),
.Y(n_9342)
);

OA21x2_ASAP7_75t_L g9343 ( 
.A1(n_9068),
.A2(n_6318),
.B(n_6316),
.Y(n_9343)
);

INVx2_ASAP7_75t_L g9344 ( 
.A(n_8692),
.Y(n_9344)
);

INVx4_ASAP7_75t_L g9345 ( 
.A(n_9026),
.Y(n_9345)
);

INVx1_ASAP7_75t_L g9346 ( 
.A(n_8906),
.Y(n_9346)
);

NAND2xp5_ASAP7_75t_L g9347 ( 
.A(n_8924),
.B(n_7495),
.Y(n_9347)
);

INVx1_ASAP7_75t_L g9348 ( 
.A(n_8907),
.Y(n_9348)
);

NAND2xp5_ASAP7_75t_SL g9349 ( 
.A(n_8941),
.B(n_6688),
.Y(n_9349)
);

INVx3_ASAP7_75t_L g9350 ( 
.A(n_8679),
.Y(n_9350)
);

INVx2_ASAP7_75t_L g9351 ( 
.A(n_8699),
.Y(n_9351)
);

CKINVDCx20_ASAP7_75t_R g9352 ( 
.A(n_8605),
.Y(n_9352)
);

CKINVDCx5p33_ASAP7_75t_R g9353 ( 
.A(n_9029),
.Y(n_9353)
);

BUFx6f_ASAP7_75t_L g9354 ( 
.A(n_8682),
.Y(n_9354)
);

CKINVDCx16_ASAP7_75t_R g9355 ( 
.A(n_8807),
.Y(n_9355)
);

CKINVDCx5p33_ASAP7_75t_R g9356 ( 
.A(n_9041),
.Y(n_9356)
);

NAND2xp5_ASAP7_75t_SL g9357 ( 
.A(n_8958),
.B(n_6870),
.Y(n_9357)
);

AND2x2_ASAP7_75t_L g9358 ( 
.A(n_8739),
.B(n_7125),
.Y(n_9358)
);

BUFx3_ASAP7_75t_L g9359 ( 
.A(n_8718),
.Y(n_9359)
);

CKINVDCx5p33_ASAP7_75t_R g9360 ( 
.A(n_9043),
.Y(n_9360)
);

INVx1_ASAP7_75t_L g9361 ( 
.A(n_8673),
.Y(n_9361)
);

CKINVDCx20_ASAP7_75t_R g9362 ( 
.A(n_9129),
.Y(n_9362)
);

AND2x2_ASAP7_75t_L g9363 ( 
.A(n_8764),
.B(n_7251),
.Y(n_9363)
);

AND2x2_ASAP7_75t_L g9364 ( 
.A(n_8782),
.B(n_7251),
.Y(n_9364)
);

AND2x2_ASAP7_75t_L g9365 ( 
.A(n_8803),
.B(n_7440),
.Y(n_9365)
);

CKINVDCx5p33_ASAP7_75t_R g9366 ( 
.A(n_9046),
.Y(n_9366)
);

CKINVDCx5p33_ASAP7_75t_R g9367 ( 
.A(n_8723),
.Y(n_9367)
);

NAND2xp5_ASAP7_75t_L g9368 ( 
.A(n_8930),
.B(n_7495),
.Y(n_9368)
);

CKINVDCx20_ASAP7_75t_R g9369 ( 
.A(n_8773),
.Y(n_9369)
);

CKINVDCx5p33_ASAP7_75t_R g9370 ( 
.A(n_8920),
.Y(n_9370)
);

INVx1_ASAP7_75t_L g9371 ( 
.A(n_8678),
.Y(n_9371)
);

INVx1_ASAP7_75t_L g9372 ( 
.A(n_8702),
.Y(n_9372)
);

INVx1_ASAP7_75t_L g9373 ( 
.A(n_8703),
.Y(n_9373)
);

INVx1_ASAP7_75t_L g9374 ( 
.A(n_8705),
.Y(n_9374)
);

CKINVDCx5p33_ASAP7_75t_R g9375 ( 
.A(n_8959),
.Y(n_9375)
);

INVx1_ASAP7_75t_L g9376 ( 
.A(n_8711),
.Y(n_9376)
);

INVx3_ASAP7_75t_L g9377 ( 
.A(n_8683),
.Y(n_9377)
);

CKINVDCx5p33_ASAP7_75t_R g9378 ( 
.A(n_9034),
.Y(n_9378)
);

BUFx6f_ASAP7_75t_L g9379 ( 
.A(n_8693),
.Y(n_9379)
);

INVx1_ASAP7_75t_L g9380 ( 
.A(n_8728),
.Y(n_9380)
);

INVx2_ASAP7_75t_L g9381 ( 
.A(n_8734),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_8743),
.Y(n_9382)
);

INVx1_ASAP7_75t_L g9383 ( 
.A(n_8746),
.Y(n_9383)
);

HB1xp67_ASAP7_75t_L g9384 ( 
.A(n_8691),
.Y(n_9384)
);

AND2x4_ASAP7_75t_L g9385 ( 
.A(n_8685),
.B(n_6326),
.Y(n_9385)
);

NOR2xp33_ASAP7_75t_R g9386 ( 
.A(n_9017),
.B(n_6946),
.Y(n_9386)
);

INVx1_ASAP7_75t_L g9387 ( 
.A(n_8747),
.Y(n_9387)
);

CKINVDCx5p33_ASAP7_75t_R g9388 ( 
.A(n_9045),
.Y(n_9388)
);

INVx1_ASAP7_75t_L g9389 ( 
.A(n_8749),
.Y(n_9389)
);

CKINVDCx5p33_ASAP7_75t_R g9390 ( 
.A(n_8580),
.Y(n_9390)
);

INVx1_ASAP7_75t_L g9391 ( 
.A(n_8753),
.Y(n_9391)
);

CKINVDCx5p33_ASAP7_75t_R g9392 ( 
.A(n_8758),
.Y(n_9392)
);

NAND2xp33_ASAP7_75t_R g9393 ( 
.A(n_8855),
.B(n_6140),
.Y(n_9393)
);

OA21x2_ASAP7_75t_L g9394 ( 
.A1(n_9081),
.A2(n_6329),
.B(n_6328),
.Y(n_9394)
);

INVx1_ASAP7_75t_L g9395 ( 
.A(n_8754),
.Y(n_9395)
);

INVx1_ASAP7_75t_L g9396 ( 
.A(n_8761),
.Y(n_9396)
);

INVx1_ASAP7_75t_L g9397 ( 
.A(n_8775),
.Y(n_9397)
);

AND2x2_ASAP7_75t_L g9398 ( 
.A(n_8966),
.B(n_7464),
.Y(n_9398)
);

NOR2xp33_ASAP7_75t_R g9399 ( 
.A(n_9037),
.B(n_8756),
.Y(n_9399)
);

CKINVDCx5p33_ASAP7_75t_R g9400 ( 
.A(n_8879),
.Y(n_9400)
);

INVx2_ASAP7_75t_L g9401 ( 
.A(n_8786),
.Y(n_9401)
);

AND2x2_ASAP7_75t_L g9402 ( 
.A(n_8881),
.B(n_7494),
.Y(n_9402)
);

BUFx3_ASAP7_75t_L g9403 ( 
.A(n_8617),
.Y(n_9403)
);

INVx2_ASAP7_75t_L g9404 ( 
.A(n_8792),
.Y(n_9404)
);

INVx3_ASAP7_75t_L g9405 ( 
.A(n_8695),
.Y(n_9405)
);

INVx3_ASAP7_75t_L g9406 ( 
.A(n_8893),
.Y(n_9406)
);

INVx3_ASAP7_75t_L g9407 ( 
.A(n_8894),
.Y(n_9407)
);

NAND2xp33_ASAP7_75t_R g9408 ( 
.A(n_8885),
.B(n_6141),
.Y(n_9408)
);

NAND2xp5_ASAP7_75t_L g9409 ( 
.A(n_8939),
.B(n_6870),
.Y(n_9409)
);

INVxp67_ASAP7_75t_L g9410 ( 
.A(n_8760),
.Y(n_9410)
);

AND2x2_ASAP7_75t_L g9411 ( 
.A(n_8698),
.B(n_6971),
.Y(n_9411)
);

CKINVDCx5p33_ASAP7_75t_R g9412 ( 
.A(n_8895),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_8813),
.Y(n_9413)
);

CKINVDCx5p33_ASAP7_75t_R g9414 ( 
.A(n_8988),
.Y(n_9414)
);

CKINVDCx5p33_ASAP7_75t_R g9415 ( 
.A(n_9011),
.Y(n_9415)
);

INVx1_ASAP7_75t_L g9416 ( 
.A(n_8814),
.Y(n_9416)
);

CKINVDCx16_ASAP7_75t_R g9417 ( 
.A(n_9070),
.Y(n_9417)
);

CKINVDCx5p33_ASAP7_75t_R g9418 ( 
.A(n_9039),
.Y(n_9418)
);

CKINVDCx5p33_ASAP7_75t_R g9419 ( 
.A(n_8995),
.Y(n_9419)
);

CKINVDCx20_ASAP7_75t_R g9420 ( 
.A(n_8801),
.Y(n_9420)
);

OAI22xp5_ASAP7_75t_L g9421 ( 
.A1(n_8794),
.A2(n_8859),
.B1(n_8866),
.B2(n_8663),
.Y(n_9421)
);

INVx2_ASAP7_75t_L g9422 ( 
.A(n_8829),
.Y(n_9422)
);

INVx2_ASAP7_75t_L g9423 ( 
.A(n_8833),
.Y(n_9423)
);

XOR2xp5_ASAP7_75t_L g9424 ( 
.A(n_8991),
.B(n_6985),
.Y(n_9424)
);

NAND2xp33_ASAP7_75t_SL g9425 ( 
.A(n_8789),
.B(n_7013),
.Y(n_9425)
);

NAND2xp5_ASAP7_75t_L g9426 ( 
.A(n_8943),
.B(n_6870),
.Y(n_9426)
);

INVx2_ASAP7_75t_L g9427 ( 
.A(n_8837),
.Y(n_9427)
);

INVx1_ASAP7_75t_L g9428 ( 
.A(n_8848),
.Y(n_9428)
);

CKINVDCx20_ASAP7_75t_R g9429 ( 
.A(n_9018),
.Y(n_9429)
);

INVx2_ASAP7_75t_L g9430 ( 
.A(n_8851),
.Y(n_9430)
);

INVx1_ASAP7_75t_L g9431 ( 
.A(n_8863),
.Y(n_9431)
);

CKINVDCx5p33_ASAP7_75t_R g9432 ( 
.A(n_9033),
.Y(n_9432)
);

INVx1_ASAP7_75t_L g9433 ( 
.A(n_8864),
.Y(n_9433)
);

CKINVDCx5p33_ASAP7_75t_R g9434 ( 
.A(n_9042),
.Y(n_9434)
);

NOR2xp33_ASAP7_75t_L g9435 ( 
.A(n_8993),
.B(n_6144),
.Y(n_9435)
);

CKINVDCx5p33_ASAP7_75t_R g9436 ( 
.A(n_9051),
.Y(n_9436)
);

CKINVDCx5p33_ASAP7_75t_R g9437 ( 
.A(n_8593),
.Y(n_9437)
);

NOR2xp33_ASAP7_75t_R g9438 ( 
.A(n_8845),
.B(n_7051),
.Y(n_9438)
);

INVx3_ASAP7_75t_L g9439 ( 
.A(n_8896),
.Y(n_9439)
);

CKINVDCx20_ASAP7_75t_R g9440 ( 
.A(n_9030),
.Y(n_9440)
);

CKINVDCx5p33_ASAP7_75t_R g9441 ( 
.A(n_9093),
.Y(n_9441)
);

CKINVDCx5p33_ASAP7_75t_R g9442 ( 
.A(n_9125),
.Y(n_9442)
);

NAND2xp5_ASAP7_75t_SL g9443 ( 
.A(n_8962),
.B(n_7086),
.Y(n_9443)
);

INVx1_ASAP7_75t_L g9444 ( 
.A(n_8878),
.Y(n_9444)
);

CKINVDCx5p33_ASAP7_75t_R g9445 ( 
.A(n_8997),
.Y(n_9445)
);

INVxp67_ASAP7_75t_L g9446 ( 
.A(n_8798),
.Y(n_9446)
);

NAND2xp5_ASAP7_75t_L g9447 ( 
.A(n_8944),
.B(n_7086),
.Y(n_9447)
);

CKINVDCx20_ASAP7_75t_R g9448 ( 
.A(n_8716),
.Y(n_9448)
);

INVx1_ASAP7_75t_L g9449 ( 
.A(n_8880),
.Y(n_9449)
);

INVx1_ASAP7_75t_L g9450 ( 
.A(n_8886),
.Y(n_9450)
);

INVxp67_ASAP7_75t_L g9451 ( 
.A(n_8811),
.Y(n_9451)
);

AND2x2_ASAP7_75t_L g9452 ( 
.A(n_8729),
.B(n_7068),
.Y(n_9452)
);

CKINVDCx5p33_ASAP7_75t_R g9453 ( 
.A(n_9062),
.Y(n_9453)
);

CKINVDCx5p33_ASAP7_75t_R g9454 ( 
.A(n_9048),
.Y(n_9454)
);

INVx1_ASAP7_75t_L g9455 ( 
.A(n_8887),
.Y(n_9455)
);

INVx4_ASAP7_75t_L g9456 ( 
.A(n_8902),
.Y(n_9456)
);

INVx1_ASAP7_75t_L g9457 ( 
.A(n_8908),
.Y(n_9457)
);

INVx2_ASAP7_75t_L g9458 ( 
.A(n_8560),
.Y(n_9458)
);

BUFx6f_ASAP7_75t_L g9459 ( 
.A(n_8909),
.Y(n_9459)
);

CKINVDCx20_ASAP7_75t_R g9460 ( 
.A(n_8719),
.Y(n_9460)
);

INVx1_ASAP7_75t_L g9461 ( 
.A(n_8911),
.Y(n_9461)
);

INVx1_ASAP7_75t_L g9462 ( 
.A(n_8883),
.Y(n_9462)
);

INVx2_ASAP7_75t_L g9463 ( 
.A(n_8892),
.Y(n_9463)
);

INVx3_ASAP7_75t_L g9464 ( 
.A(n_8915),
.Y(n_9464)
);

CKINVDCx5p33_ASAP7_75t_R g9465 ( 
.A(n_8623),
.Y(n_9465)
);

AND2x2_ASAP7_75t_L g9466 ( 
.A(n_8731),
.B(n_8976),
.Y(n_9466)
);

CKINVDCx5p33_ASAP7_75t_R g9467 ( 
.A(n_8634),
.Y(n_9467)
);

BUFx6f_ASAP7_75t_L g9468 ( 
.A(n_8589),
.Y(n_9468)
);

CKINVDCx5p33_ASAP7_75t_R g9469 ( 
.A(n_9065),
.Y(n_9469)
);

INVx1_ASAP7_75t_L g9470 ( 
.A(n_8921),
.Y(n_9470)
);

HB1xp67_ASAP7_75t_L g9471 ( 
.A(n_8694),
.Y(n_9471)
);

AND2x2_ASAP7_75t_L g9472 ( 
.A(n_8827),
.B(n_7075),
.Y(n_9472)
);

CKINVDCx5p33_ASAP7_75t_R g9473 ( 
.A(n_8994),
.Y(n_9473)
);

BUFx6f_ASAP7_75t_L g9474 ( 
.A(n_8606),
.Y(n_9474)
);

INVx1_ASAP7_75t_L g9475 ( 
.A(n_8935),
.Y(n_9475)
);

CKINVDCx20_ASAP7_75t_R g9476 ( 
.A(n_8922),
.Y(n_9476)
);

BUFx10_ASAP7_75t_L g9477 ( 
.A(n_9000),
.Y(n_9477)
);

AND2x4_ASAP7_75t_L g9478 ( 
.A(n_9080),
.B(n_9085),
.Y(n_9478)
);

CKINVDCx20_ASAP7_75t_R g9479 ( 
.A(n_8973),
.Y(n_9479)
);

BUFx6f_ASAP7_75t_L g9480 ( 
.A(n_8616),
.Y(n_9480)
);

INVx1_ASAP7_75t_L g9481 ( 
.A(n_8624),
.Y(n_9481)
);

BUFx6f_ASAP7_75t_L g9482 ( 
.A(n_8626),
.Y(n_9482)
);

INVx1_ASAP7_75t_SL g9483 ( 
.A(n_8839),
.Y(n_9483)
);

INVx1_ASAP7_75t_L g9484 ( 
.A(n_8632),
.Y(n_9484)
);

INVx1_ASAP7_75t_L g9485 ( 
.A(n_8636),
.Y(n_9485)
);

BUFx6f_ASAP7_75t_L g9486 ( 
.A(n_8628),
.Y(n_9486)
);

INVx1_ASAP7_75t_L g9487 ( 
.A(n_8637),
.Y(n_9487)
);

CKINVDCx5p33_ASAP7_75t_R g9488 ( 
.A(n_8996),
.Y(n_9488)
);

INVx3_ASAP7_75t_L g9489 ( 
.A(n_8575),
.Y(n_9489)
);

BUFx2_ASAP7_75t_L g9490 ( 
.A(n_8644),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_8638),
.Y(n_9491)
);

INVxp67_ASAP7_75t_L g9492 ( 
.A(n_8821),
.Y(n_9492)
);

INVx1_ASAP7_75t_L g9493 ( 
.A(n_8647),
.Y(n_9493)
);

HB1xp67_ASAP7_75t_L g9494 ( 
.A(n_9005),
.Y(n_9494)
);

CKINVDCx5p33_ASAP7_75t_R g9495 ( 
.A(n_8999),
.Y(n_9495)
);

INVx1_ASAP7_75t_L g9496 ( 
.A(n_8653),
.Y(n_9496)
);

NOR2xp33_ASAP7_75t_L g9497 ( 
.A(n_9014),
.B(n_6145),
.Y(n_9497)
);

INVx2_ASAP7_75t_L g9498 ( 
.A(n_8657),
.Y(n_9498)
);

NOR2xp33_ASAP7_75t_R g9499 ( 
.A(n_9059),
.B(n_7097),
.Y(n_9499)
);

BUFx2_ASAP7_75t_L g9500 ( 
.A(n_8697),
.Y(n_9500)
);

INVx2_ASAP7_75t_L g9501 ( 
.A(n_8649),
.Y(n_9501)
);

INVx2_ASAP7_75t_L g9502 ( 
.A(n_8655),
.Y(n_9502)
);

NAND2xp5_ASAP7_75t_L g9503 ( 
.A(n_8952),
.B(n_7086),
.Y(n_9503)
);

CKINVDCx5p33_ASAP7_75t_R g9504 ( 
.A(n_9025),
.Y(n_9504)
);

NOR2xp67_ASAP7_75t_L g9505 ( 
.A(n_8884),
.B(n_4549),
.Y(n_9505)
);

INVx3_ASAP7_75t_L g9506 ( 
.A(n_8650),
.Y(n_9506)
);

INVx2_ASAP7_75t_L g9507 ( 
.A(n_8550),
.Y(n_9507)
);

INVx1_ASAP7_75t_L g9508 ( 
.A(n_8819),
.Y(n_9508)
);

INVx3_ASAP7_75t_L g9509 ( 
.A(n_8651),
.Y(n_9509)
);

INVx2_ASAP7_75t_L g9510 ( 
.A(n_8553),
.Y(n_9510)
);

AND2x4_ASAP7_75t_L g9511 ( 
.A(n_8568),
.B(n_6332),
.Y(n_9511)
);

BUFx2_ASAP7_75t_L g9512 ( 
.A(n_8697),
.Y(n_9512)
);

INVx1_ASAP7_75t_L g9513 ( 
.A(n_8953),
.Y(n_9513)
);

AND2x2_ASAP7_75t_L g9514 ( 
.A(n_8918),
.B(n_7111),
.Y(n_9514)
);

HB1xp67_ASAP7_75t_L g9515 ( 
.A(n_8707),
.Y(n_9515)
);

INVx2_ASAP7_75t_L g9516 ( 
.A(n_8557),
.Y(n_9516)
);

CKINVDCx5p33_ASAP7_75t_R g9517 ( 
.A(n_9027),
.Y(n_9517)
);

INVx1_ASAP7_75t_L g9518 ( 
.A(n_8965),
.Y(n_9518)
);

AND2x4_ASAP7_75t_L g9519 ( 
.A(n_8844),
.B(n_6341),
.Y(n_9519)
);

AND2x2_ASAP7_75t_L g9520 ( 
.A(n_8932),
.B(n_7126),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8714),
.Y(n_9521)
);

AND2x6_ASAP7_75t_L g9522 ( 
.A(n_8972),
.B(n_7122),
.Y(n_9522)
);

INVx1_ASAP7_75t_L g9523 ( 
.A(n_8766),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_8768),
.Y(n_9524)
);

INVx1_ASAP7_75t_L g9525 ( 
.A(n_8788),
.Y(n_9525)
);

INVx1_ASAP7_75t_L g9526 ( 
.A(n_8795),
.Y(n_9526)
);

NAND2xp5_ASAP7_75t_L g9527 ( 
.A(n_8578),
.B(n_7122),
.Y(n_9527)
);

CKINVDCx5p33_ASAP7_75t_R g9528 ( 
.A(n_9028),
.Y(n_9528)
);

INVx1_ASAP7_75t_L g9529 ( 
.A(n_8809),
.Y(n_9529)
);

CKINVDCx5p33_ASAP7_75t_R g9530 ( 
.A(n_9044),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_8840),
.Y(n_9531)
);

INVx1_ASAP7_75t_L g9532 ( 
.A(n_8849),
.Y(n_9532)
);

BUFx3_ASAP7_75t_L g9533 ( 
.A(n_8964),
.Y(n_9533)
);

BUFx6f_ASAP7_75t_L g9534 ( 
.A(n_8664),
.Y(n_9534)
);

CKINVDCx5p33_ASAP7_75t_R g9535 ( 
.A(n_9047),
.Y(n_9535)
);

INVx2_ASAP7_75t_L g9536 ( 
.A(n_9078),
.Y(n_9536)
);

AND2x2_ASAP7_75t_L g9537 ( 
.A(n_8732),
.B(n_9058),
.Y(n_9537)
);

INVx1_ASAP7_75t_L g9538 ( 
.A(n_8854),
.Y(n_9538)
);

CKINVDCx5p33_ASAP7_75t_R g9539 ( 
.A(n_9054),
.Y(n_9539)
);

INVx2_ASAP7_75t_L g9540 ( 
.A(n_9096),
.Y(n_9540)
);

INVx1_ASAP7_75t_L g9541 ( 
.A(n_8847),
.Y(n_9541)
);

INVxp67_ASAP7_75t_L g9542 ( 
.A(n_9056),
.Y(n_9542)
);

INVx1_ASAP7_75t_L g9543 ( 
.A(n_8852),
.Y(n_9543)
);

CKINVDCx5p33_ASAP7_75t_R g9544 ( 
.A(n_9002),
.Y(n_9544)
);

INVx2_ASAP7_75t_L g9545 ( 
.A(n_9107),
.Y(n_9545)
);

BUFx6f_ASAP7_75t_L g9546 ( 
.A(n_8710),
.Y(n_9546)
);

CKINVDCx5p33_ASAP7_75t_R g9547 ( 
.A(n_9006),
.Y(n_9547)
);

INVx2_ASAP7_75t_L g9548 ( 
.A(n_9109),
.Y(n_9548)
);

INVx4_ASAP7_75t_L g9549 ( 
.A(n_8717),
.Y(n_9549)
);

INVx1_ASAP7_75t_L g9550 ( 
.A(n_8861),
.Y(n_9550)
);

NOR2xp33_ASAP7_75t_R g9551 ( 
.A(n_9007),
.B(n_7171),
.Y(n_9551)
);

INVx2_ASAP7_75t_L g9552 ( 
.A(n_9127),
.Y(n_9552)
);

NAND2xp5_ASAP7_75t_L g9553 ( 
.A(n_8934),
.B(n_7122),
.Y(n_9553)
);

NOR2xp67_ASAP7_75t_L g9554 ( 
.A(n_9009),
.B(n_4551),
.Y(n_9554)
);

CKINVDCx20_ASAP7_75t_R g9555 ( 
.A(n_9004),
.Y(n_9555)
);

INVx3_ASAP7_75t_L g9556 ( 
.A(n_8721),
.Y(n_9556)
);

INVx3_ASAP7_75t_L g9557 ( 
.A(n_8744),
.Y(n_9557)
);

NAND2xp5_ASAP7_75t_SL g9558 ( 
.A(n_8607),
.B(n_7322),
.Y(n_9558)
);

HB1xp67_ASAP7_75t_L g9559 ( 
.A(n_9001),
.Y(n_9559)
);

INVx2_ASAP7_75t_L g9560 ( 
.A(n_9128),
.Y(n_9560)
);

INVx1_ASAP7_75t_L g9561 ( 
.A(n_8889),
.Y(n_9561)
);

NAND2xp5_ASAP7_75t_SL g9562 ( 
.A(n_8654),
.B(n_7322),
.Y(n_9562)
);

INVx5_ASAP7_75t_L g9563 ( 
.A(n_8810),
.Y(n_9563)
);

OAI22xp5_ASAP7_75t_L g9564 ( 
.A1(n_8986),
.A2(n_8957),
.B1(n_8938),
.B2(n_8715),
.Y(n_9564)
);

INVx2_ASAP7_75t_L g9565 ( 
.A(n_8737),
.Y(n_9565)
);

CKINVDCx20_ASAP7_75t_R g9566 ( 
.A(n_8763),
.Y(n_9566)
);

INVx1_ASAP7_75t_L g9567 ( 
.A(n_8923),
.Y(n_9567)
);

CKINVDCx20_ASAP7_75t_R g9568 ( 
.A(n_9057),
.Y(n_9568)
);

INVx2_ASAP7_75t_L g9569 ( 
.A(n_8745),
.Y(n_9569)
);

CKINVDCx5p33_ASAP7_75t_R g9570 ( 
.A(n_9010),
.Y(n_9570)
);

INVx1_ASAP7_75t_L g9571 ( 
.A(n_8955),
.Y(n_9571)
);

CKINVDCx20_ASAP7_75t_R g9572 ( 
.A(n_8891),
.Y(n_9572)
);

INVx2_ASAP7_75t_L g9573 ( 
.A(n_8752),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_8822),
.Y(n_9574)
);

CKINVDCx20_ASAP7_75t_R g9575 ( 
.A(n_8945),
.Y(n_9575)
);

INVx2_ASAP7_75t_L g9576 ( 
.A(n_8759),
.Y(n_9576)
);

BUFx3_ASAP7_75t_L g9577 ( 
.A(n_8765),
.Y(n_9577)
);

INVx1_ASAP7_75t_L g9578 ( 
.A(n_9111),
.Y(n_9578)
);

CKINVDCx5p33_ASAP7_75t_R g9579 ( 
.A(n_9013),
.Y(n_9579)
);

INVx2_ASAP7_75t_L g9580 ( 
.A(n_8770),
.Y(n_9580)
);

AND2x2_ASAP7_75t_L g9581 ( 
.A(n_8690),
.B(n_7189),
.Y(n_9581)
);

INVx3_ASAP7_75t_L g9582 ( 
.A(n_8772),
.Y(n_9582)
);

NOR2xp33_ASAP7_75t_SL g9583 ( 
.A(n_8987),
.B(n_7194),
.Y(n_9583)
);

INVx1_ASAP7_75t_L g9584 ( 
.A(n_8778),
.Y(n_9584)
);

CKINVDCx5p33_ASAP7_75t_R g9585 ( 
.A(n_9016),
.Y(n_9585)
);

AND2x6_ASAP7_75t_L g9586 ( 
.A(n_8970),
.B(n_7322),
.Y(n_9586)
);

INVx1_ASAP7_75t_L g9587 ( 
.A(n_8779),
.Y(n_9587)
);

NAND2xp5_ASAP7_75t_L g9588 ( 
.A(n_8582),
.B(n_7415),
.Y(n_9588)
);

INVx2_ASAP7_75t_L g9589 ( 
.A(n_8793),
.Y(n_9589)
);

INVx1_ASAP7_75t_L g9590 ( 
.A(n_8800),
.Y(n_9590)
);

NAND2xp5_ASAP7_75t_L g9591 ( 
.A(n_8591),
.B(n_8968),
.Y(n_9591)
);

HB1xp67_ASAP7_75t_L g9592 ( 
.A(n_8736),
.Y(n_9592)
);

INVx2_ASAP7_75t_L g9593 ( 
.A(n_8802),
.Y(n_9593)
);

AND2x2_ASAP7_75t_L g9594 ( 
.A(n_8989),
.B(n_7203),
.Y(n_9594)
);

INVx1_ASAP7_75t_L g9595 ( 
.A(n_8806),
.Y(n_9595)
);

BUFx6f_ASAP7_75t_L g9596 ( 
.A(n_8808),
.Y(n_9596)
);

AND2x2_ASAP7_75t_SL g9597 ( 
.A(n_8983),
.B(n_6289),
.Y(n_9597)
);

NOR2xp33_ASAP7_75t_R g9598 ( 
.A(n_9020),
.B(n_7224),
.Y(n_9598)
);

NAND2xp5_ASAP7_75t_L g9599 ( 
.A(n_8969),
.B(n_7415),
.Y(n_9599)
);

CKINVDCx5p33_ASAP7_75t_R g9600 ( 
.A(n_9021),
.Y(n_9600)
);

CKINVDCx5p33_ASAP7_75t_R g9601 ( 
.A(n_9023),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_8812),
.Y(n_9602)
);

BUFx6f_ASAP7_75t_L g9603 ( 
.A(n_8824),
.Y(n_9603)
);

CKINVDCx5p33_ASAP7_75t_R g9604 ( 
.A(n_9035),
.Y(n_9604)
);

CKINVDCx20_ASAP7_75t_R g9605 ( 
.A(n_9038),
.Y(n_9605)
);

INVxp67_ASAP7_75t_L g9606 ( 
.A(n_8750),
.Y(n_9606)
);

INVx1_ASAP7_75t_L g9607 ( 
.A(n_8834),
.Y(n_9607)
);

INVx1_ASAP7_75t_L g9608 ( 
.A(n_8850),
.Y(n_9608)
);

CKINVDCx5p33_ASAP7_75t_R g9609 ( 
.A(n_9040),
.Y(n_9609)
);

INVx2_ASAP7_75t_L g9610 ( 
.A(n_8857),
.Y(n_9610)
);

INVx2_ASAP7_75t_L g9611 ( 
.A(n_8858),
.Y(n_9611)
);

INVx1_ASAP7_75t_L g9612 ( 
.A(n_8876),
.Y(n_9612)
);

INVx1_ASAP7_75t_L g9613 ( 
.A(n_8890),
.Y(n_9613)
);

AND2x2_ASAP7_75t_SL g9614 ( 
.A(n_9022),
.B(n_6306),
.Y(n_9614)
);

CKINVDCx5p33_ASAP7_75t_R g9615 ( 
.A(n_9053),
.Y(n_9615)
);

CKINVDCx5p33_ASAP7_75t_R g9616 ( 
.A(n_9055),
.Y(n_9616)
);

INVx1_ASAP7_75t_L g9617 ( 
.A(n_8700),
.Y(n_9617)
);

CKINVDCx5p33_ASAP7_75t_R g9618 ( 
.A(n_8865),
.Y(n_9618)
);

CKINVDCx5p33_ASAP7_75t_R g9619 ( 
.A(n_8865),
.Y(n_9619)
);

CKINVDCx20_ASAP7_75t_R g9620 ( 
.A(n_8913),
.Y(n_9620)
);

CKINVDCx20_ASAP7_75t_R g9621 ( 
.A(n_8984),
.Y(n_9621)
);

BUFx6f_ASAP7_75t_L g9622 ( 
.A(n_9049),
.Y(n_9622)
);

CKINVDCx5p33_ASAP7_75t_R g9623 ( 
.A(n_8805),
.Y(n_9623)
);

NOR2xp33_ASAP7_75t_R g9624 ( 
.A(n_8992),
.B(n_7236),
.Y(n_9624)
);

CKINVDCx20_ASAP7_75t_R g9625 ( 
.A(n_8990),
.Y(n_9625)
);

INVx2_ASAP7_75t_L g9626 ( 
.A(n_8713),
.Y(n_9626)
);

CKINVDCx5p33_ASAP7_75t_R g9627 ( 
.A(n_8674),
.Y(n_9627)
);

CKINVDCx5p33_ASAP7_75t_R g9628 ( 
.A(n_9032),
.Y(n_9628)
);

CKINVDCx20_ASAP7_75t_R g9629 ( 
.A(n_8835),
.Y(n_9629)
);

CKINVDCx5p33_ASAP7_75t_R g9630 ( 
.A(n_8916),
.Y(n_9630)
);

HB1xp67_ASAP7_75t_L g9631 ( 
.A(n_8771),
.Y(n_9631)
);

BUFx10_ASAP7_75t_L g9632 ( 
.A(n_9003),
.Y(n_9632)
);

BUFx6f_ASAP7_75t_L g9633 ( 
.A(n_8596),
.Y(n_9633)
);

INVx1_ASAP7_75t_L g9634 ( 
.A(n_8722),
.Y(n_9634)
);

INVx1_ASAP7_75t_SL g9635 ( 
.A(n_9060),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_8556),
.Y(n_9636)
);

INVx3_ASAP7_75t_L g9637 ( 
.A(n_8797),
.Y(n_9637)
);

CKINVDCx20_ASAP7_75t_R g9638 ( 
.A(n_9031),
.Y(n_9638)
);

INVx1_ASAP7_75t_L g9639 ( 
.A(n_8726),
.Y(n_9639)
);

CKINVDCx5p33_ASAP7_75t_R g9640 ( 
.A(n_9131),
.Y(n_9640)
);

INVx1_ASAP7_75t_L g9641 ( 
.A(n_8757),
.Y(n_9641)
);

CKINVDCx5p33_ASAP7_75t_R g9642 ( 
.A(n_8810),
.Y(n_9642)
);

AND2x2_ASAP7_75t_L g9643 ( 
.A(n_9123),
.B(n_7239),
.Y(n_9643)
);

HB1xp67_ASAP7_75t_L g9644 ( 
.A(n_8826),
.Y(n_9644)
);

CKINVDCx5p33_ASAP7_75t_R g9645 ( 
.A(n_9131),
.Y(n_9645)
);

AND2x2_ASAP7_75t_L g9646 ( 
.A(n_8831),
.B(n_7284),
.Y(n_9646)
);

INVx1_ASAP7_75t_L g9647 ( 
.A(n_8785),
.Y(n_9647)
);

CKINVDCx20_ASAP7_75t_R g9648 ( 
.A(n_8804),
.Y(n_9648)
);

CKINVDCx5p33_ASAP7_75t_R g9649 ( 
.A(n_8869),
.Y(n_9649)
);

BUFx6f_ASAP7_75t_L g9650 ( 
.A(n_8629),
.Y(n_9650)
);

INVx1_ASAP7_75t_L g9651 ( 
.A(n_8836),
.Y(n_9651)
);

INVx1_ASAP7_75t_L g9652 ( 
.A(n_8631),
.Y(n_9652)
);

INVx3_ASAP7_75t_L g9653 ( 
.A(n_8633),
.Y(n_9653)
);

INVx2_ASAP7_75t_L g9654 ( 
.A(n_8733),
.Y(n_9654)
);

INVx1_ASAP7_75t_L g9655 ( 
.A(n_8645),
.Y(n_9655)
);

NAND2xp5_ASAP7_75t_L g9656 ( 
.A(n_8791),
.B(n_7415),
.Y(n_9656)
);

CKINVDCx5p33_ASAP7_75t_R g9657 ( 
.A(n_8869),
.Y(n_9657)
);

NAND2xp5_ASAP7_75t_L g9658 ( 
.A(n_8877),
.B(n_8625),
.Y(n_9658)
);

CKINVDCx5p33_ASAP7_75t_R g9659 ( 
.A(n_8552),
.Y(n_9659)
);

INVx1_ASAP7_75t_L g9660 ( 
.A(n_8720),
.Y(n_9660)
);

INVx1_ASAP7_75t_L g9661 ( 
.A(n_8725),
.Y(n_9661)
);

CKINVDCx5p33_ASAP7_75t_R g9662 ( 
.A(n_8774),
.Y(n_9662)
);

CKINVDCx5p33_ASAP7_75t_R g9663 ( 
.A(n_8946),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_8790),
.Y(n_9664)
);

OA21x2_ASAP7_75t_L g9665 ( 
.A1(n_9094),
.A2(n_9102),
.B(n_8977),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_8867),
.Y(n_9666)
);

OAI22xp5_ASAP7_75t_L g9667 ( 
.A1(n_9117),
.A2(n_7451),
.B1(n_6148),
.B2(n_6150),
.Y(n_9667)
);

INVx1_ASAP7_75t_L g9668 ( 
.A(n_8872),
.Y(n_9668)
);

CKINVDCx5p33_ASAP7_75t_R g9669 ( 
.A(n_8948),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_SL g9670 ( 
.A(n_8640),
.B(n_7451),
.Y(n_9670)
);

INVx1_ASAP7_75t_L g9671 ( 
.A(n_9083),
.Y(n_9671)
);

CKINVDCx5p33_ASAP7_75t_R g9672 ( 
.A(n_8956),
.Y(n_9672)
);

AND2x4_ASAP7_75t_L g9673 ( 
.A(n_8648),
.B(n_6344),
.Y(n_9673)
);

CKINVDCx20_ASAP7_75t_R g9674 ( 
.A(n_9063),
.Y(n_9674)
);

BUFx6f_ASAP7_75t_L g9675 ( 
.A(n_8975),
.Y(n_9675)
);

INVx1_ASAP7_75t_L g9676 ( 
.A(n_9100),
.Y(n_9676)
);

CKINVDCx5p33_ASAP7_75t_R g9677 ( 
.A(n_8554),
.Y(n_9677)
);

INVx2_ASAP7_75t_L g9678 ( 
.A(n_8708),
.Y(n_9678)
);

INVx1_ASAP7_75t_L g9679 ( 
.A(n_8985),
.Y(n_9679)
);

AND2x2_ASAP7_75t_L g9680 ( 
.A(n_8727),
.B(n_7295),
.Y(n_9680)
);

INVx1_ASAP7_75t_L g9681 ( 
.A(n_8597),
.Y(n_9681)
);

INVx1_ASAP7_75t_L g9682 ( 
.A(n_8668),
.Y(n_9682)
);

BUFx6f_ASAP7_75t_L g9683 ( 
.A(n_8799),
.Y(n_9683)
);

OAI21x1_ASAP7_75t_L g9684 ( 
.A1(n_8817),
.A2(n_6361),
.B(n_6314),
.Y(n_9684)
);

AND2x2_ASAP7_75t_L g9685 ( 
.A(n_8820),
.B(n_7298),
.Y(n_9685)
);

CKINVDCx20_ASAP7_75t_R g9686 ( 
.A(n_9036),
.Y(n_9686)
);

OAI21x1_ASAP7_75t_L g9687 ( 
.A1(n_8870),
.A2(n_6399),
.B(n_6363),
.Y(n_9687)
);

CKINVDCx5p33_ASAP7_75t_R g9688 ( 
.A(n_8980),
.Y(n_9688)
);

CKINVDCx20_ASAP7_75t_R g9689 ( 
.A(n_8846),
.Y(n_9689)
);

INVx2_ASAP7_75t_L g9690 ( 
.A(n_8675),
.Y(n_9690)
);

INVx1_ASAP7_75t_L g9691 ( 
.A(n_8680),
.Y(n_9691)
);

NAND2x1_ASAP7_75t_L g9692 ( 
.A(n_8818),
.B(n_7451),
.Y(n_9692)
);

NAND2xp5_ASAP7_75t_SL g9693 ( 
.A(n_8642),
.B(n_6147),
.Y(n_9693)
);

CKINVDCx20_ASAP7_75t_R g9694 ( 
.A(n_8954),
.Y(n_9694)
);

NAND2xp5_ASAP7_75t_L g9695 ( 
.A(n_8652),
.B(n_6152),
.Y(n_9695)
);

CKINVDCx5p33_ASAP7_75t_R g9696 ( 
.A(n_8823),
.Y(n_9696)
);

BUFx6f_ASAP7_75t_L g9697 ( 
.A(n_9337),
.Y(n_9697)
);

INVx2_ASAP7_75t_L g9698 ( 
.A(n_9136),
.Y(n_9698)
);

NAND2xp5_ASAP7_75t_L g9699 ( 
.A(n_9639),
.B(n_9591),
.Y(n_9699)
);

INVx1_ASAP7_75t_SL g9700 ( 
.A(n_9483),
.Y(n_9700)
);

INVx1_ASAP7_75t_L g9701 ( 
.A(n_9135),
.Y(n_9701)
);

AND2x2_ASAP7_75t_L g9702 ( 
.A(n_9134),
.B(n_9398),
.Y(n_9702)
);

HB1xp67_ASAP7_75t_L g9703 ( 
.A(n_9172),
.Y(n_9703)
);

INVxp67_ASAP7_75t_L g9704 ( 
.A(n_9152),
.Y(n_9704)
);

OAI22xp5_ASAP7_75t_SL g9705 ( 
.A1(n_9555),
.A2(n_7313),
.B1(n_7325),
.B2(n_7312),
.Y(n_9705)
);

AND2x2_ASAP7_75t_L g9706 ( 
.A(n_9365),
.B(n_8978),
.Y(n_9706)
);

INVxp67_ASAP7_75t_L g9707 ( 
.A(n_9188),
.Y(n_9707)
);

INVxp67_ASAP7_75t_L g9708 ( 
.A(n_9330),
.Y(n_9708)
);

OAI22xp5_ASAP7_75t_SL g9709 ( 
.A1(n_9566),
.A2(n_7393),
.B1(n_7399),
.B2(n_7385),
.Y(n_9709)
);

BUFx2_ASAP7_75t_L g9710 ( 
.A(n_9217),
.Y(n_9710)
);

INVxp67_ASAP7_75t_L g9711 ( 
.A(n_9402),
.Y(n_9711)
);

INVx2_ASAP7_75t_L g9712 ( 
.A(n_9159),
.Y(n_9712)
);

INVx2_ASAP7_75t_L g9713 ( 
.A(n_9164),
.Y(n_9713)
);

INVx2_ASAP7_75t_L g9714 ( 
.A(n_9170),
.Y(n_9714)
);

OAI22xp5_ASAP7_75t_SL g9715 ( 
.A1(n_9424),
.A2(n_7481),
.B1(n_7518),
.B2(n_7419),
.Y(n_9715)
);

INVx2_ASAP7_75t_L g9716 ( 
.A(n_9183),
.Y(n_9716)
);

INVx2_ASAP7_75t_L g9717 ( 
.A(n_9193),
.Y(n_9717)
);

NAND2xp33_ASAP7_75t_SL g9718 ( 
.A(n_9399),
.B(n_8926),
.Y(n_9718)
);

INVx1_ASAP7_75t_L g9719 ( 
.A(n_9137),
.Y(n_9719)
);

BUFx2_ASAP7_75t_L g9720 ( 
.A(n_9257),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_9139),
.Y(n_9721)
);

BUFx6f_ASAP7_75t_L g9722 ( 
.A(n_9337),
.Y(n_9722)
);

HB1xp67_ASAP7_75t_L g9723 ( 
.A(n_9210),
.Y(n_9723)
);

OAI22xp5_ASAP7_75t_SL g9724 ( 
.A1(n_9686),
.A2(n_6158),
.B1(n_6159),
.B2(n_6156),
.Y(n_9724)
);

OAI22xp5_ASAP7_75t_SL g9725 ( 
.A1(n_9689),
.A2(n_6164),
.B1(n_6168),
.B2(n_6161),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_9146),
.Y(n_9726)
);

INVx2_ASAP7_75t_L g9727 ( 
.A(n_9200),
.Y(n_9727)
);

INVx2_ASAP7_75t_L g9728 ( 
.A(n_9202),
.Y(n_9728)
);

INVx1_ASAP7_75t_L g9729 ( 
.A(n_9156),
.Y(n_9729)
);

NAND2xp33_ASAP7_75t_SL g9730 ( 
.A(n_9618),
.B(n_8618),
.Y(n_9730)
);

INVx1_ASAP7_75t_L g9731 ( 
.A(n_9160),
.Y(n_9731)
);

OAI21x1_ASAP7_75t_L g9732 ( 
.A1(n_9288),
.A2(n_8838),
.B(n_8874),
.Y(n_9732)
);

INVx2_ASAP7_75t_L g9733 ( 
.A(n_9206),
.Y(n_9733)
);

INVx1_ASAP7_75t_L g9734 ( 
.A(n_9167),
.Y(n_9734)
);

NAND2xp5_ASAP7_75t_SL g9735 ( 
.A(n_9628),
.B(n_8677),
.Y(n_9735)
);

BUFx6f_ASAP7_75t_L g9736 ( 
.A(n_9359),
.Y(n_9736)
);

NAND2xp5_ASAP7_75t_SL g9737 ( 
.A(n_9421),
.B(n_8599),
.Y(n_9737)
);

OAI22xp33_ASAP7_75t_L g9738 ( 
.A1(n_9155),
.A2(n_8882),
.B1(n_6170),
.B2(n_6171),
.Y(n_9738)
);

INVx1_ASAP7_75t_L g9739 ( 
.A(n_9178),
.Y(n_9739)
);

BUFx6f_ASAP7_75t_L g9740 ( 
.A(n_9354),
.Y(n_9740)
);

AND2x2_ASAP7_75t_L g9741 ( 
.A(n_9466),
.B(n_9061),
.Y(n_9741)
);

BUFx6f_ASAP7_75t_L g9742 ( 
.A(n_9354),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_9215),
.Y(n_9743)
);

INVx2_ASAP7_75t_L g9744 ( 
.A(n_9179),
.Y(n_9744)
);

NAND2xp5_ASAP7_75t_SL g9745 ( 
.A(n_9630),
.B(n_6169),
.Y(n_9745)
);

INVx1_ASAP7_75t_L g9746 ( 
.A(n_9185),
.Y(n_9746)
);

OAI22xp5_ASAP7_75t_SL g9747 ( 
.A1(n_9694),
.A2(n_6179),
.B1(n_6181),
.B2(n_6175),
.Y(n_9747)
);

INVx2_ASAP7_75t_L g9748 ( 
.A(n_9186),
.Y(n_9748)
);

AND2x2_ASAP7_75t_L g9749 ( 
.A(n_9275),
.B(n_6183),
.Y(n_9749)
);

INVx2_ASAP7_75t_L g9750 ( 
.A(n_9190),
.Y(n_9750)
);

INVx2_ASAP7_75t_L g9751 ( 
.A(n_9194),
.Y(n_9751)
);

BUFx6f_ASAP7_75t_L g9752 ( 
.A(n_9379),
.Y(n_9752)
);

INVx2_ASAP7_75t_L g9753 ( 
.A(n_9196),
.Y(n_9753)
);

INVx1_ASAP7_75t_L g9754 ( 
.A(n_9198),
.Y(n_9754)
);

NAND2xp5_ASAP7_75t_L g9755 ( 
.A(n_9578),
.B(n_6871),
.Y(n_9755)
);

INVx1_ASAP7_75t_L g9756 ( 
.A(n_9203),
.Y(n_9756)
);

INVxp67_ASAP7_75t_L g9757 ( 
.A(n_9177),
.Y(n_9757)
);

INVx2_ASAP7_75t_L g9758 ( 
.A(n_9204),
.Y(n_9758)
);

BUFx6f_ASAP7_75t_L g9759 ( 
.A(n_9379),
.Y(n_9759)
);

INVx1_ASAP7_75t_L g9760 ( 
.A(n_9207),
.Y(n_9760)
);

BUFx6f_ASAP7_75t_L g9761 ( 
.A(n_9546),
.Y(n_9761)
);

INVx1_ASAP7_75t_L g9762 ( 
.A(n_9208),
.Y(n_9762)
);

INVx2_ASAP7_75t_L g9763 ( 
.A(n_9212),
.Y(n_9763)
);

INVx1_ASAP7_75t_L g9764 ( 
.A(n_9213),
.Y(n_9764)
);

INVx1_ASAP7_75t_SL g9765 ( 
.A(n_9490),
.Y(n_9765)
);

INVx1_ASAP7_75t_L g9766 ( 
.A(n_9225),
.Y(n_9766)
);

INVx1_ASAP7_75t_L g9767 ( 
.A(n_9229),
.Y(n_9767)
);

INVx1_ASAP7_75t_L g9768 ( 
.A(n_9231),
.Y(n_9768)
);

NAND2xp5_ASAP7_75t_L g9769 ( 
.A(n_9243),
.B(n_7167),
.Y(n_9769)
);

INVx1_ASAP7_75t_L g9770 ( 
.A(n_9232),
.Y(n_9770)
);

NAND2xp5_ASAP7_75t_SL g9771 ( 
.A(n_9305),
.B(n_6187),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_9234),
.Y(n_9772)
);

INVx2_ASAP7_75t_L g9773 ( 
.A(n_9241),
.Y(n_9773)
);

NAND2xp5_ASAP7_75t_L g9774 ( 
.A(n_9660),
.B(n_6191),
.Y(n_9774)
);

OAI22xp5_ASAP7_75t_SL g9775 ( 
.A1(n_9688),
.A2(n_6197),
.B1(n_6198),
.B2(n_6194),
.Y(n_9775)
);

INVx1_ASAP7_75t_L g9776 ( 
.A(n_9242),
.Y(n_9776)
);

INVx1_ASAP7_75t_L g9777 ( 
.A(n_9244),
.Y(n_9777)
);

AND2x4_ASAP7_75t_L g9778 ( 
.A(n_9533),
.B(n_6346),
.Y(n_9778)
);

INVx2_ASAP7_75t_L g9779 ( 
.A(n_9246),
.Y(n_9779)
);

INVx1_ASAP7_75t_L g9780 ( 
.A(n_9254),
.Y(n_9780)
);

INVx3_ASAP7_75t_L g9781 ( 
.A(n_9546),
.Y(n_9781)
);

INVx2_ASAP7_75t_L g9782 ( 
.A(n_9258),
.Y(n_9782)
);

AND2x6_ASAP7_75t_L g9783 ( 
.A(n_9661),
.B(n_6349),
.Y(n_9783)
);

INVx2_ASAP7_75t_L g9784 ( 
.A(n_9259),
.Y(n_9784)
);

INVx2_ASAP7_75t_L g9785 ( 
.A(n_9267),
.Y(n_9785)
);

INVx1_ASAP7_75t_L g9786 ( 
.A(n_9270),
.Y(n_9786)
);

INVx1_ASAP7_75t_L g9787 ( 
.A(n_9283),
.Y(n_9787)
);

NAND2xp5_ASAP7_75t_SL g9788 ( 
.A(n_9597),
.B(n_6200),
.Y(n_9788)
);

INVx3_ASAP7_75t_L g9789 ( 
.A(n_9596),
.Y(n_9789)
);

INVxp67_ASAP7_75t_L g9790 ( 
.A(n_9184),
.Y(n_9790)
);

INVx2_ASAP7_75t_L g9791 ( 
.A(n_9284),
.Y(n_9791)
);

INVx2_ASAP7_75t_L g9792 ( 
.A(n_9287),
.Y(n_9792)
);

NAND2xp5_ASAP7_75t_SL g9793 ( 
.A(n_9614),
.B(n_6202),
.Y(n_9793)
);

INVx1_ASAP7_75t_L g9794 ( 
.A(n_9292),
.Y(n_9794)
);

INVx1_ASAP7_75t_L g9795 ( 
.A(n_9297),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_9298),
.Y(n_9796)
);

INVx2_ASAP7_75t_L g9797 ( 
.A(n_9302),
.Y(n_9797)
);

INVx2_ASAP7_75t_L g9798 ( 
.A(n_9303),
.Y(n_9798)
);

OAI22xp5_ASAP7_75t_SL g9799 ( 
.A1(n_9623),
.A2(n_6208),
.B1(n_6210),
.B2(n_6206),
.Y(n_9799)
);

INVx1_ASAP7_75t_L g9800 ( 
.A(n_9306),
.Y(n_9800)
);

AND2x2_ASAP7_75t_L g9801 ( 
.A(n_9331),
.B(n_6213),
.Y(n_9801)
);

INVxp67_ASAP7_75t_L g9802 ( 
.A(n_9329),
.Y(n_9802)
);

OAI22xp5_ASAP7_75t_L g9803 ( 
.A1(n_9542),
.A2(n_6217),
.B1(n_6219),
.B2(n_6215),
.Y(n_9803)
);

INVx1_ASAP7_75t_L g9804 ( 
.A(n_9315),
.Y(n_9804)
);

NAND2xp33_ASAP7_75t_SL g9805 ( 
.A(n_9619),
.B(n_6222),
.Y(n_9805)
);

INVx1_ASAP7_75t_L g9806 ( 
.A(n_9319),
.Y(n_9806)
);

INVx2_ASAP7_75t_L g9807 ( 
.A(n_9321),
.Y(n_9807)
);

NOR2xp33_ASAP7_75t_L g9808 ( 
.A(n_9606),
.B(n_6224),
.Y(n_9808)
);

INVx2_ASAP7_75t_L g9809 ( 
.A(n_9322),
.Y(n_9809)
);

HB1xp67_ASAP7_75t_L g9810 ( 
.A(n_9314),
.Y(n_9810)
);

INVx3_ASAP7_75t_L g9811 ( 
.A(n_9596),
.Y(n_9811)
);

INVx1_ASAP7_75t_L g9812 ( 
.A(n_9326),
.Y(n_9812)
);

INVx1_ASAP7_75t_L g9813 ( 
.A(n_9327),
.Y(n_9813)
);

INVxp67_ASAP7_75t_L g9814 ( 
.A(n_9163),
.Y(n_9814)
);

INVx2_ASAP7_75t_L g9815 ( 
.A(n_9328),
.Y(n_9815)
);

INVx1_ASAP7_75t_L g9816 ( 
.A(n_9332),
.Y(n_9816)
);

NAND2xp5_ASAP7_75t_L g9817 ( 
.A(n_9664),
.B(n_6226),
.Y(n_9817)
);

INVx2_ASAP7_75t_L g9818 ( 
.A(n_9333),
.Y(n_9818)
);

INVx1_ASAP7_75t_L g9819 ( 
.A(n_9334),
.Y(n_9819)
);

NAND2xp5_ASAP7_75t_SL g9820 ( 
.A(n_9473),
.B(n_6229),
.Y(n_9820)
);

INVx1_ASAP7_75t_SL g9821 ( 
.A(n_9205),
.Y(n_9821)
);

INVx2_ASAP7_75t_L g9822 ( 
.A(n_9458),
.Y(n_9822)
);

NAND2xp5_ASAP7_75t_SL g9823 ( 
.A(n_9488),
.B(n_6232),
.Y(n_9823)
);

INVxp67_ASAP7_75t_L g9824 ( 
.A(n_9168),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_9339),
.Y(n_9825)
);

NAND2xp5_ASAP7_75t_L g9826 ( 
.A(n_9658),
.B(n_6238),
.Y(n_9826)
);

INVx1_ASAP7_75t_L g9827 ( 
.A(n_9342),
.Y(n_9827)
);

OAI22xp5_ASAP7_75t_L g9828 ( 
.A1(n_9636),
.A2(n_6243),
.B1(n_6244),
.B2(n_6240),
.Y(n_9828)
);

BUFx6f_ASAP7_75t_L g9829 ( 
.A(n_9603),
.Y(n_9829)
);

INVx2_ASAP7_75t_L g9830 ( 
.A(n_9346),
.Y(n_9830)
);

INVx1_ASAP7_75t_L g9831 ( 
.A(n_9348),
.Y(n_9831)
);

OAI21x1_ASAP7_75t_L g9832 ( 
.A1(n_9684),
.A2(n_6432),
.B(n_6417),
.Y(n_9832)
);

NAND2xp5_ASAP7_75t_L g9833 ( 
.A(n_9435),
.B(n_9497),
.Y(n_9833)
);

AND2x4_ASAP7_75t_L g9834 ( 
.A(n_9345),
.B(n_6355),
.Y(n_9834)
);

INVx2_ASAP7_75t_L g9835 ( 
.A(n_9293),
.Y(n_9835)
);

OAI22xp5_ASAP7_75t_L g9836 ( 
.A1(n_9142),
.A2(n_6252),
.B1(n_6256),
.B2(n_6248),
.Y(n_9836)
);

INVx1_ASAP7_75t_L g9837 ( 
.A(n_9513),
.Y(n_9837)
);

BUFx6f_ASAP7_75t_L g9838 ( 
.A(n_9603),
.Y(n_9838)
);

HB1xp67_ASAP7_75t_L g9839 ( 
.A(n_9384),
.Y(n_9839)
);

HB1xp67_ASAP7_75t_L g9840 ( 
.A(n_9214),
.Y(n_9840)
);

AND2x2_ASAP7_75t_L g9841 ( 
.A(n_9358),
.B(n_6262),
.Y(n_9841)
);

BUFx6f_ASAP7_75t_SL g9842 ( 
.A(n_9296),
.Y(n_9842)
);

INVx1_ASAP7_75t_SL g9843 ( 
.A(n_9195),
.Y(n_9843)
);

INVx1_ASAP7_75t_L g9844 ( 
.A(n_9518),
.Y(n_9844)
);

INVx2_ASAP7_75t_L g9845 ( 
.A(n_9304),
.Y(n_9845)
);

AND2x4_ASAP7_75t_L g9846 ( 
.A(n_9161),
.B(n_9169),
.Y(n_9846)
);

BUFx6f_ASAP7_75t_L g9847 ( 
.A(n_9151),
.Y(n_9847)
);

INVx2_ASAP7_75t_L g9848 ( 
.A(n_9312),
.Y(n_9848)
);

NAND2xp5_ASAP7_75t_SL g9849 ( 
.A(n_9495),
.B(n_6268),
.Y(n_9849)
);

INVx1_ASAP7_75t_L g9850 ( 
.A(n_9281),
.Y(n_9850)
);

NAND2xp5_ASAP7_75t_L g9851 ( 
.A(n_9695),
.B(n_6272),
.Y(n_9851)
);

CKINVDCx16_ASAP7_75t_R g9852 ( 
.A(n_9311),
.Y(n_9852)
);

INVx2_ASAP7_75t_L g9853 ( 
.A(n_9316),
.Y(n_9853)
);

INVx1_ASAP7_75t_L g9854 ( 
.A(n_9291),
.Y(n_9854)
);

INVx1_ASAP7_75t_L g9855 ( 
.A(n_9372),
.Y(n_9855)
);

INVx1_ASAP7_75t_L g9856 ( 
.A(n_9373),
.Y(n_9856)
);

XOR2xp5_ASAP7_75t_L g9857 ( 
.A(n_9166),
.B(n_4552),
.Y(n_9857)
);

INVx2_ASAP7_75t_L g9858 ( 
.A(n_9318),
.Y(n_9858)
);

INVx2_ASAP7_75t_L g9859 ( 
.A(n_9344),
.Y(n_9859)
);

INVx1_ASAP7_75t_L g9860 ( 
.A(n_9374),
.Y(n_9860)
);

INVx1_ASAP7_75t_L g9861 ( 
.A(n_9376),
.Y(n_9861)
);

AOI22xp5_ASAP7_75t_L g9862 ( 
.A1(n_9289),
.A2(n_6274),
.B1(n_6275),
.B2(n_6273),
.Y(n_9862)
);

OAI22xp33_ASAP7_75t_L g9863 ( 
.A1(n_9659),
.A2(n_6282),
.B1(n_6284),
.B2(n_6280),
.Y(n_9863)
);

INVx1_ASAP7_75t_L g9864 ( 
.A(n_9380),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_9382),
.Y(n_9865)
);

AND2x2_ASAP7_75t_L g9866 ( 
.A(n_9363),
.B(n_6290),
.Y(n_9866)
);

INVx1_ASAP7_75t_SL g9867 ( 
.A(n_9572),
.Y(n_9867)
);

INVxp33_ASAP7_75t_L g9868 ( 
.A(n_9252),
.Y(n_9868)
);

INVx1_ASAP7_75t_L g9869 ( 
.A(n_9383),
.Y(n_9869)
);

NOR2xp33_ASAP7_75t_L g9870 ( 
.A(n_9492),
.B(n_6291),
.Y(n_9870)
);

INVx2_ASAP7_75t_L g9871 ( 
.A(n_9351),
.Y(n_9871)
);

INVx2_ASAP7_75t_L g9872 ( 
.A(n_9381),
.Y(n_9872)
);

INVx1_ASAP7_75t_L g9873 ( 
.A(n_9387),
.Y(n_9873)
);

INVxp67_ASAP7_75t_L g9874 ( 
.A(n_9364),
.Y(n_9874)
);

INVx1_ASAP7_75t_L g9875 ( 
.A(n_9389),
.Y(n_9875)
);

INVx1_ASAP7_75t_L g9876 ( 
.A(n_9391),
.Y(n_9876)
);

INVx1_ASAP7_75t_L g9877 ( 
.A(n_9395),
.Y(n_9877)
);

INVx2_ASAP7_75t_L g9878 ( 
.A(n_9401),
.Y(n_9878)
);

NAND3xp33_ASAP7_75t_SL g9879 ( 
.A(n_9499),
.B(n_6295),
.C(n_6293),
.Y(n_9879)
);

INVx1_ASAP7_75t_L g9880 ( 
.A(n_9396),
.Y(n_9880)
);

NAND2xp33_ASAP7_75t_SL g9881 ( 
.A(n_9390),
.B(n_6297),
.Y(n_9881)
);

INVx1_ASAP7_75t_L g9882 ( 
.A(n_9397),
.Y(n_9882)
);

AND2x4_ASAP7_75t_L g9883 ( 
.A(n_9403),
.B(n_6359),
.Y(n_9883)
);

INVx1_ASAP7_75t_L g9884 ( 
.A(n_9413),
.Y(n_9884)
);

INVx2_ASAP7_75t_L g9885 ( 
.A(n_9404),
.Y(n_9885)
);

INVx2_ASAP7_75t_L g9886 ( 
.A(n_9422),
.Y(n_9886)
);

INVx1_ASAP7_75t_SL g9887 ( 
.A(n_9575),
.Y(n_9887)
);

BUFx6f_ASAP7_75t_L g9888 ( 
.A(n_9151),
.Y(n_9888)
);

INVx1_ASAP7_75t_L g9889 ( 
.A(n_9416),
.Y(n_9889)
);

CKINVDCx20_ASAP7_75t_R g9890 ( 
.A(n_9290),
.Y(n_9890)
);

INVx2_ASAP7_75t_L g9891 ( 
.A(n_9423),
.Y(n_9891)
);

INVxp67_ASAP7_75t_L g9892 ( 
.A(n_9253),
.Y(n_9892)
);

AOI22x1_ASAP7_75t_L g9893 ( 
.A1(n_9641),
.A2(n_6302),
.B1(n_6307),
.B2(n_6300),
.Y(n_9893)
);

INVx1_ASAP7_75t_L g9894 ( 
.A(n_9428),
.Y(n_9894)
);

INVx1_ASAP7_75t_SL g9895 ( 
.A(n_9471),
.Y(n_9895)
);

INVx1_ASAP7_75t_L g9896 ( 
.A(n_9431),
.Y(n_9896)
);

INVx2_ASAP7_75t_L g9897 ( 
.A(n_9427),
.Y(n_9897)
);

INVx1_ASAP7_75t_L g9898 ( 
.A(n_9433),
.Y(n_9898)
);

OAI22xp5_ASAP7_75t_SL g9899 ( 
.A1(n_9677),
.A2(n_6320),
.B1(n_6323),
.B2(n_6308),
.Y(n_9899)
);

INVx2_ASAP7_75t_L g9900 ( 
.A(n_9430),
.Y(n_9900)
);

NAND2xp5_ASAP7_75t_L g9901 ( 
.A(n_9553),
.B(n_6325),
.Y(n_9901)
);

INVx1_ASAP7_75t_L g9902 ( 
.A(n_9444),
.Y(n_9902)
);

INVx2_ASAP7_75t_L g9903 ( 
.A(n_9221),
.Y(n_9903)
);

INVx1_ASAP7_75t_L g9904 ( 
.A(n_9449),
.Y(n_9904)
);

INVx1_ASAP7_75t_L g9905 ( 
.A(n_9450),
.Y(n_9905)
);

INVx2_ASAP7_75t_L g9906 ( 
.A(n_9228),
.Y(n_9906)
);

INVx3_ASAP7_75t_L g9907 ( 
.A(n_9459),
.Y(n_9907)
);

NAND2xp5_ASAP7_75t_L g9908 ( 
.A(n_9192),
.B(n_6335),
.Y(n_9908)
);

AND2x6_ASAP7_75t_L g9909 ( 
.A(n_9622),
.B(n_6365),
.Y(n_9909)
);

INVx1_ASAP7_75t_L g9910 ( 
.A(n_9455),
.Y(n_9910)
);

AOI22xp5_ASAP7_75t_L g9911 ( 
.A1(n_9559),
.A2(n_6338),
.B1(n_6339),
.B2(n_6337),
.Y(n_9911)
);

INVx3_ASAP7_75t_L g9912 ( 
.A(n_9459),
.Y(n_9912)
);

NAND2xp5_ASAP7_75t_L g9913 ( 
.A(n_9201),
.B(n_6340),
.Y(n_9913)
);

INVx1_ASAP7_75t_L g9914 ( 
.A(n_9271),
.Y(n_9914)
);

INVx2_ASAP7_75t_L g9915 ( 
.A(n_9236),
.Y(n_9915)
);

NAND2xp5_ASAP7_75t_L g9916 ( 
.A(n_9237),
.B(n_6342),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_9272),
.Y(n_9917)
);

INVx2_ASAP7_75t_L g9918 ( 
.A(n_9268),
.Y(n_9918)
);

AOI22xp5_ASAP7_75t_L g9919 ( 
.A1(n_9696),
.A2(n_9635),
.B1(n_9574),
.B2(n_9564),
.Y(n_9919)
);

INVx2_ASAP7_75t_L g9920 ( 
.A(n_9269),
.Y(n_9920)
);

AND2x4_ASAP7_75t_L g9921 ( 
.A(n_9577),
.B(n_6367),
.Y(n_9921)
);

OAI22xp5_ASAP7_75t_SL g9922 ( 
.A1(n_9629),
.A2(n_9638),
.B1(n_9479),
.B2(n_9476),
.Y(n_9922)
);

INVx1_ASAP7_75t_L g9923 ( 
.A(n_9282),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_9481),
.Y(n_9924)
);

NAND2xp33_ASAP7_75t_SL g9925 ( 
.A(n_9392),
.B(n_6345),
.Y(n_9925)
);

INVx3_ASAP7_75t_L g9926 ( 
.A(n_9468),
.Y(n_9926)
);

BUFx6f_ASAP7_75t_L g9927 ( 
.A(n_9174),
.Y(n_9927)
);

NAND2xp33_ASAP7_75t_SL g9928 ( 
.A(n_9400),
.B(n_9412),
.Y(n_9928)
);

BUFx6f_ASAP7_75t_L g9929 ( 
.A(n_9174),
.Y(n_9929)
);

INVx1_ASAP7_75t_L g9930 ( 
.A(n_9484),
.Y(n_9930)
);

INVx3_ASAP7_75t_L g9931 ( 
.A(n_9468),
.Y(n_9931)
);

INVx1_ASAP7_75t_L g9932 ( 
.A(n_9485),
.Y(n_9932)
);

INVxp67_ASAP7_75t_L g9933 ( 
.A(n_9262),
.Y(n_9933)
);

AND2x2_ASAP7_75t_L g9934 ( 
.A(n_9515),
.B(n_6348),
.Y(n_9934)
);

INVx2_ASAP7_75t_SL g9935 ( 
.A(n_9537),
.Y(n_9935)
);

NAND2xp5_ASAP7_75t_SL g9936 ( 
.A(n_9504),
.B(n_6351),
.Y(n_9936)
);

INVx2_ASAP7_75t_L g9937 ( 
.A(n_9278),
.Y(n_9937)
);

INVx1_ASAP7_75t_L g9938 ( 
.A(n_9487),
.Y(n_9938)
);

INVx1_ASAP7_75t_L g9939 ( 
.A(n_9491),
.Y(n_9939)
);

INVx2_ASAP7_75t_L g9940 ( 
.A(n_9498),
.Y(n_9940)
);

BUFx6f_ASAP7_75t_L g9941 ( 
.A(n_9176),
.Y(n_9941)
);

INVx2_ASAP7_75t_L g9942 ( 
.A(n_9493),
.Y(n_9942)
);

INVx1_ASAP7_75t_L g9943 ( 
.A(n_9496),
.Y(n_9943)
);

INVx1_ASAP7_75t_L g9944 ( 
.A(n_9507),
.Y(n_9944)
);

INVx2_ASAP7_75t_L g9945 ( 
.A(n_9220),
.Y(n_9945)
);

INVx1_ASAP7_75t_L g9946 ( 
.A(n_9510),
.Y(n_9946)
);

INVx2_ASAP7_75t_L g9947 ( 
.A(n_9565),
.Y(n_9947)
);

NAND2xp5_ASAP7_75t_SL g9948 ( 
.A(n_9517),
.B(n_6352),
.Y(n_9948)
);

INVx3_ASAP7_75t_L g9949 ( 
.A(n_9474),
.Y(n_9949)
);

BUFx6f_ASAP7_75t_L g9950 ( 
.A(n_9176),
.Y(n_9950)
);

AND2x2_ASAP7_75t_L g9951 ( 
.A(n_9508),
.B(n_6358),
.Y(n_9951)
);

AND2x2_ASAP7_75t_L g9952 ( 
.A(n_9514),
.B(n_6364),
.Y(n_9952)
);

INVx1_ASAP7_75t_L g9953 ( 
.A(n_9516),
.Y(n_9953)
);

INVx1_ASAP7_75t_L g9954 ( 
.A(n_9536),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_L g9955 ( 
.A(n_9249),
.B(n_6369),
.Y(n_9955)
);

INVx1_ASAP7_75t_L g9956 ( 
.A(n_9540),
.Y(n_9956)
);

INVx1_ASAP7_75t_L g9957 ( 
.A(n_9545),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_9548),
.Y(n_9958)
);

INVx2_ASAP7_75t_L g9959 ( 
.A(n_9552),
.Y(n_9959)
);

INVx1_ASAP7_75t_L g9960 ( 
.A(n_9560),
.Y(n_9960)
);

INVx1_ASAP7_75t_L g9961 ( 
.A(n_9457),
.Y(n_9961)
);

OAI22xp5_ASAP7_75t_L g9962 ( 
.A1(n_9554),
.A2(n_6371),
.B1(n_6372),
.B2(n_6370),
.Y(n_9962)
);

INVx2_ASAP7_75t_L g9963 ( 
.A(n_9501),
.Y(n_9963)
);

BUFx6f_ASAP7_75t_L g9964 ( 
.A(n_9180),
.Y(n_9964)
);

INVx1_ASAP7_75t_L g9965 ( 
.A(n_9461),
.Y(n_9965)
);

INVx2_ASAP7_75t_L g9966 ( 
.A(n_9502),
.Y(n_9966)
);

NAND2xp5_ASAP7_75t_L g9967 ( 
.A(n_9141),
.B(n_6375),
.Y(n_9967)
);

INVx1_ASAP7_75t_L g9968 ( 
.A(n_9462),
.Y(n_9968)
);

INVx1_ASAP7_75t_L g9969 ( 
.A(n_9361),
.Y(n_9969)
);

INVx1_ASAP7_75t_L g9970 ( 
.A(n_9371),
.Y(n_9970)
);

INVx2_ASAP7_75t_L g9971 ( 
.A(n_9489),
.Y(n_9971)
);

AOI22xp5_ASAP7_75t_L g9972 ( 
.A1(n_9335),
.A2(n_6376),
.B1(n_6378),
.B2(n_6377),
.Y(n_9972)
);

INVx1_ASAP7_75t_L g9973 ( 
.A(n_9521),
.Y(n_9973)
);

INVx2_ASAP7_75t_L g9974 ( 
.A(n_9523),
.Y(n_9974)
);

INVx2_ASAP7_75t_L g9975 ( 
.A(n_9524),
.Y(n_9975)
);

AOI22xp5_ASAP7_75t_L g9976 ( 
.A1(n_9347),
.A2(n_6379),
.B1(n_6386),
.B2(n_6380),
.Y(n_9976)
);

INVx2_ASAP7_75t_L g9977 ( 
.A(n_9525),
.Y(n_9977)
);

INVx1_ASAP7_75t_L g9978 ( 
.A(n_9526),
.Y(n_9978)
);

AND2x2_ASAP7_75t_L g9979 ( 
.A(n_9520),
.B(n_6387),
.Y(n_9979)
);

NAND2xp33_ASAP7_75t_SL g9980 ( 
.A(n_9414),
.B(n_6389),
.Y(n_9980)
);

NOR2x1_ASAP7_75t_L g9981 ( 
.A(n_9456),
.B(n_6374),
.Y(n_9981)
);

INVx1_ASAP7_75t_L g9982 ( 
.A(n_9529),
.Y(n_9982)
);

INVx1_ASAP7_75t_L g9983 ( 
.A(n_9531),
.Y(n_9983)
);

INVx1_ASAP7_75t_L g9984 ( 
.A(n_9532),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_9538),
.Y(n_9985)
);

BUFx6f_ASAP7_75t_L g9986 ( 
.A(n_9180),
.Y(n_9986)
);

INVx1_ASAP7_75t_L g9987 ( 
.A(n_9266),
.Y(n_9987)
);

INVx1_ASAP7_75t_L g9988 ( 
.A(n_9279),
.Y(n_9988)
);

NAND2x1p5_ASAP7_75t_L g9989 ( 
.A(n_9549),
.B(n_6384),
.Y(n_9989)
);

BUFx6f_ASAP7_75t_L g9990 ( 
.A(n_9187),
.Y(n_9990)
);

BUFx2_ASAP7_75t_L g9991 ( 
.A(n_9625),
.Y(n_9991)
);

INVx1_ASAP7_75t_L g9992 ( 
.A(n_9313),
.Y(n_9992)
);

HB1xp67_ASAP7_75t_L g9993 ( 
.A(n_9410),
.Y(n_9993)
);

NOR2xp33_ASAP7_75t_L g9994 ( 
.A(n_9446),
.B(n_6392),
.Y(n_9994)
);

INVx1_ASAP7_75t_L g9995 ( 
.A(n_9368),
.Y(n_9995)
);

INVx1_ASAP7_75t_L g9996 ( 
.A(n_9197),
.Y(n_9996)
);

INVx1_ASAP7_75t_L g9997 ( 
.A(n_9230),
.Y(n_9997)
);

NAND2xp5_ASAP7_75t_SL g9998 ( 
.A(n_9528),
.B(n_6393),
.Y(n_9998)
);

BUFx6f_ASAP7_75t_L g9999 ( 
.A(n_9187),
.Y(n_9999)
);

INVx2_ASAP7_75t_L g10000 ( 
.A(n_9690),
.Y(n_10000)
);

INVx1_ASAP7_75t_L g10001 ( 
.A(n_9325),
.Y(n_10001)
);

BUFx2_ASAP7_75t_L g10002 ( 
.A(n_9274),
.Y(n_10002)
);

INVx1_ASAP7_75t_L g10003 ( 
.A(n_9470),
.Y(n_10003)
);

INVx1_ASAP7_75t_L g10004 ( 
.A(n_9475),
.Y(n_10004)
);

INVxp67_ASAP7_75t_L g10005 ( 
.A(n_9594),
.Y(n_10005)
);

INVx3_ASAP7_75t_L g10006 ( 
.A(n_9474),
.Y(n_10006)
);

AND2x6_ASAP7_75t_L g10007 ( 
.A(n_9622),
.B(n_6390),
.Y(n_10007)
);

INVx2_ASAP7_75t_L g10008 ( 
.A(n_9678),
.Y(n_10008)
);

XOR2xp5_ASAP7_75t_L g10009 ( 
.A(n_9173),
.B(n_4553),
.Y(n_10009)
);

NAND2xp5_ASAP7_75t_SL g10010 ( 
.A(n_9530),
.B(n_6396),
.Y(n_10010)
);

INVx1_ASAP7_75t_L g10011 ( 
.A(n_9409),
.Y(n_10011)
);

INVx1_ASAP7_75t_L g10012 ( 
.A(n_9426),
.Y(n_10012)
);

INVx1_ASAP7_75t_L g10013 ( 
.A(n_9447),
.Y(n_10013)
);

INVx1_ASAP7_75t_SL g10014 ( 
.A(n_9411),
.Y(n_10014)
);

INVx2_ASAP7_75t_L g10015 ( 
.A(n_9681),
.Y(n_10015)
);

NAND2xp5_ASAP7_75t_L g10016 ( 
.A(n_9656),
.B(n_6401),
.Y(n_10016)
);

INVx1_ASAP7_75t_L g10017 ( 
.A(n_9503),
.Y(n_10017)
);

INVx1_ASAP7_75t_SL g10018 ( 
.A(n_9452),
.Y(n_10018)
);

INVx2_ASAP7_75t_L g10019 ( 
.A(n_9682),
.Y(n_10019)
);

INVx2_ASAP7_75t_L g10020 ( 
.A(n_9691),
.Y(n_10020)
);

AOI22xp5_ASAP7_75t_L g10021 ( 
.A1(n_9535),
.A2(n_6404),
.B1(n_6405),
.B2(n_6403),
.Y(n_10021)
);

INVx1_ASAP7_75t_L g10022 ( 
.A(n_9541),
.Y(n_10022)
);

AND2x2_ASAP7_75t_L g10023 ( 
.A(n_9472),
.B(n_6409),
.Y(n_10023)
);

INVx3_ASAP7_75t_L g10024 ( 
.A(n_9480),
.Y(n_10024)
);

INVx1_ASAP7_75t_L g10025 ( 
.A(n_9543),
.Y(n_10025)
);

OAI22xp5_ASAP7_75t_L g10026 ( 
.A1(n_9539),
.A2(n_6419),
.B1(n_6421),
.B2(n_6410),
.Y(n_10026)
);

INVx3_ASAP7_75t_L g10027 ( 
.A(n_9480),
.Y(n_10027)
);

OAI21x1_ASAP7_75t_L g10028 ( 
.A1(n_9626),
.A2(n_6451),
.B(n_6447),
.Y(n_10028)
);

INVx2_ASAP7_75t_L g10029 ( 
.A(n_9647),
.Y(n_10029)
);

INVx1_ASAP7_75t_L g10030 ( 
.A(n_9550),
.Y(n_10030)
);

BUFx6f_ASAP7_75t_L g10031 ( 
.A(n_9209),
.Y(n_10031)
);

INVx1_ASAP7_75t_L g10032 ( 
.A(n_9561),
.Y(n_10032)
);

OAI22xp5_ASAP7_75t_SL g10033 ( 
.A1(n_9388),
.A2(n_6425),
.B1(n_6426),
.B2(n_6422),
.Y(n_10033)
);

NOR2xp33_ASAP7_75t_L g10034 ( 
.A(n_9451),
.B(n_6427),
.Y(n_10034)
);

INVx1_ASAP7_75t_SL g10035 ( 
.A(n_9419),
.Y(n_10035)
);

OAI22xp5_ASAP7_75t_L g10036 ( 
.A1(n_9679),
.A2(n_6433),
.B1(n_6435),
.B2(n_6429),
.Y(n_10036)
);

INVx3_ASAP7_75t_L g10037 ( 
.A(n_9482),
.Y(n_10037)
);

CKINVDCx8_ASAP7_75t_R g10038 ( 
.A(n_9150),
.Y(n_10038)
);

NAND2xp33_ASAP7_75t_SL g10039 ( 
.A(n_9415),
.B(n_6440),
.Y(n_10039)
);

NAND2xp5_ASAP7_75t_L g10040 ( 
.A(n_9154),
.B(n_6443),
.Y(n_10040)
);

INVx2_ASAP7_75t_L g10041 ( 
.A(n_9651),
.Y(n_10041)
);

AND2x4_ASAP7_75t_L g10042 ( 
.A(n_9324),
.B(n_6394),
.Y(n_10042)
);

OA21x2_ASAP7_75t_L g10043 ( 
.A1(n_9671),
.A2(n_6398),
.B(n_6395),
.Y(n_10043)
);

INVx2_ASAP7_75t_L g10044 ( 
.A(n_9666),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9567),
.Y(n_10045)
);

BUFx6f_ASAP7_75t_L g10046 ( 
.A(n_9209),
.Y(n_10046)
);

INVx1_ASAP7_75t_L g10047 ( 
.A(n_9571),
.Y(n_10047)
);

NOR3xp33_ASAP7_75t_SL g10048 ( 
.A(n_9393),
.B(n_6450),
.C(n_6446),
.Y(n_10048)
);

INVx1_ASAP7_75t_L g10049 ( 
.A(n_9340),
.Y(n_10049)
);

INVx5_ASAP7_75t_L g10050 ( 
.A(n_9632),
.Y(n_10050)
);

BUFx6f_ASAP7_75t_SL g10051 ( 
.A(n_9175),
.Y(n_10051)
);

INVx1_ASAP7_75t_L g10052 ( 
.A(n_9511),
.Y(n_10052)
);

INVx1_ASAP7_75t_L g10053 ( 
.A(n_9227),
.Y(n_10053)
);

INVx2_ASAP7_75t_L g10054 ( 
.A(n_9668),
.Y(n_10054)
);

INVx2_ASAP7_75t_L g10055 ( 
.A(n_9676),
.Y(n_10055)
);

HB1xp67_ASAP7_75t_L g10056 ( 
.A(n_9494),
.Y(n_10056)
);

INVx1_ASAP7_75t_L g10057 ( 
.A(n_9248),
.Y(n_10057)
);

NAND2xp5_ASAP7_75t_SL g10058 ( 
.A(n_9454),
.B(n_6455),
.Y(n_10058)
);

INVx1_ASAP7_75t_L g10059 ( 
.A(n_9250),
.Y(n_10059)
);

NAND2xp5_ASAP7_75t_L g10060 ( 
.A(n_9154),
.B(n_6458),
.Y(n_10060)
);

NAND2xp5_ASAP7_75t_L g10061 ( 
.A(n_9154),
.B(n_6461),
.Y(n_10061)
);

INVx3_ASAP7_75t_L g10062 ( 
.A(n_9482),
.Y(n_10062)
);

INVx2_ASAP7_75t_L g10063 ( 
.A(n_9654),
.Y(n_10063)
);

OAI22xp5_ASAP7_75t_SL g10064 ( 
.A1(n_9417),
.A2(n_6480),
.B1(n_6482),
.B2(n_6463),
.Y(n_10064)
);

INVx2_ASAP7_75t_L g10065 ( 
.A(n_9463),
.Y(n_10065)
);

AND3x1_ASAP7_75t_L g10066 ( 
.A(n_9583),
.B(n_6408),
.C(n_6406),
.Y(n_10066)
);

AND2x4_ASAP7_75t_L g10067 ( 
.A(n_9506),
.B(n_6412),
.Y(n_10067)
);

AOI22xp5_ASAP7_75t_L g10068 ( 
.A1(n_9693),
.A2(n_6486),
.B1(n_6488),
.B2(n_6485),
.Y(n_10068)
);

INVx1_ASAP7_75t_L g10069 ( 
.A(n_9584),
.Y(n_10069)
);

INVx8_ASAP7_75t_L g10070 ( 
.A(n_9323),
.Y(n_10070)
);

INVx2_ASAP7_75t_L g10071 ( 
.A(n_9569),
.Y(n_10071)
);

INVx2_ASAP7_75t_L g10072 ( 
.A(n_9573),
.Y(n_10072)
);

AND2x2_ASAP7_75t_L g10073 ( 
.A(n_9581),
.B(n_6491),
.Y(n_10073)
);

NAND2xp5_ASAP7_75t_L g10074 ( 
.A(n_9157),
.B(n_6492),
.Y(n_10074)
);

INVx2_ASAP7_75t_L g10075 ( 
.A(n_9576),
.Y(n_10075)
);

INVx2_ASAP7_75t_L g10076 ( 
.A(n_9580),
.Y(n_10076)
);

AND2x4_ASAP7_75t_L g10077 ( 
.A(n_9509),
.B(n_6416),
.Y(n_10077)
);

INVx1_ASAP7_75t_L g10078 ( 
.A(n_9587),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_9590),
.Y(n_10079)
);

HB1xp67_ASAP7_75t_L g10080 ( 
.A(n_9140),
.Y(n_10080)
);

INVx1_ASAP7_75t_L g10081 ( 
.A(n_9595),
.Y(n_10081)
);

INVx1_ASAP7_75t_L g10082 ( 
.A(n_9607),
.Y(n_10082)
);

AND2x2_ASAP7_75t_SL g10083 ( 
.A(n_9189),
.B(n_6474),
.Y(n_10083)
);

INVx3_ASAP7_75t_L g10084 ( 
.A(n_9486),
.Y(n_10084)
);

BUFx8_ASAP7_75t_L g10085 ( 
.A(n_9500),
.Y(n_10085)
);

INVx1_ASAP7_75t_L g10086 ( 
.A(n_9608),
.Y(n_10086)
);

INVx2_ASAP7_75t_L g10087 ( 
.A(n_9589),
.Y(n_10087)
);

OAI22xp5_ASAP7_75t_SL g10088 ( 
.A1(n_9662),
.A2(n_6499),
.B1(n_6503),
.B2(n_6497),
.Y(n_10088)
);

NAND2xp5_ASAP7_75t_L g10089 ( 
.A(n_9157),
.B(n_6505),
.Y(n_10089)
);

INVx1_ASAP7_75t_L g10090 ( 
.A(n_9612),
.Y(n_10090)
);

AND2x2_ASAP7_75t_L g10091 ( 
.A(n_9477),
.B(n_9680),
.Y(n_10091)
);

INVx1_ASAP7_75t_SL g10092 ( 
.A(n_9432),
.Y(n_10092)
);

OAI22xp5_ASAP7_75t_L g10093 ( 
.A1(n_9544),
.A2(n_6508),
.B1(n_6510),
.B2(n_6506),
.Y(n_10093)
);

INVx1_ASAP7_75t_L g10094 ( 
.A(n_9613),
.Y(n_10094)
);

INVx2_ASAP7_75t_L g10095 ( 
.A(n_9593),
.Y(n_10095)
);

OAI22xp33_ASAP7_75t_L g10096 ( 
.A1(n_9547),
.A2(n_6515),
.B1(n_6516),
.B2(n_6512),
.Y(n_10096)
);

NAND2xp33_ASAP7_75t_SL g10097 ( 
.A(n_9418),
.B(n_6523),
.Y(n_10097)
);

NAND2xp33_ASAP7_75t_L g10098 ( 
.A(n_9157),
.B(n_6524),
.Y(n_10098)
);

INVx1_ASAP7_75t_L g10099 ( 
.A(n_9602),
.Y(n_10099)
);

INVx1_ASAP7_75t_L g10100 ( 
.A(n_9610),
.Y(n_10100)
);

OAI22xp5_ASAP7_75t_L g10101 ( 
.A1(n_9570),
.A2(n_6526),
.B1(n_6527),
.B2(n_6525),
.Y(n_10101)
);

INVx1_ASAP7_75t_L g10102 ( 
.A(n_9611),
.Y(n_10102)
);

AND2x2_ASAP7_75t_L g10103 ( 
.A(n_9646),
.B(n_6528),
.Y(n_10103)
);

OAI22xp5_ASAP7_75t_L g10104 ( 
.A1(n_9579),
.A2(n_6531),
.B1(n_6532),
.B2(n_6529),
.Y(n_10104)
);

INVx2_ASAP7_75t_L g10105 ( 
.A(n_9133),
.Y(n_10105)
);

INVx2_ASAP7_75t_L g10106 ( 
.A(n_9148),
.Y(n_10106)
);

INVx1_ASAP7_75t_L g10107 ( 
.A(n_9519),
.Y(n_10107)
);

CKINVDCx8_ASAP7_75t_R g10108 ( 
.A(n_9153),
.Y(n_10108)
);

NAND2xp5_ASAP7_75t_SL g10109 ( 
.A(n_9563),
.B(n_6539),
.Y(n_10109)
);

AOI22xp5_ASAP7_75t_L g10110 ( 
.A1(n_9585),
.A2(n_6543),
.B1(n_6544),
.B2(n_6540),
.Y(n_10110)
);

INVx2_ASAP7_75t_L g10111 ( 
.A(n_9486),
.Y(n_10111)
);

INVxp67_ASAP7_75t_L g10112 ( 
.A(n_9631),
.Y(n_10112)
);

INVx1_ASAP7_75t_L g10113 ( 
.A(n_9617),
.Y(n_10113)
);

NOR2xp33_ASAP7_75t_L g10114 ( 
.A(n_9600),
.B(n_6547),
.Y(n_10114)
);

AOI22xp5_ASAP7_75t_L g10115 ( 
.A1(n_9601),
.A2(n_6554),
.B1(n_6557),
.B2(n_6548),
.Y(n_10115)
);

NAND2xp5_ASAP7_75t_SL g10116 ( 
.A(n_9563),
.B(n_6563),
.Y(n_10116)
);

INVx2_ASAP7_75t_L g10117 ( 
.A(n_9534),
.Y(n_10117)
);

AND2x2_ASAP7_75t_L g10118 ( 
.A(n_9604),
.B(n_6569),
.Y(n_10118)
);

INVx1_ASAP7_75t_SL g10119 ( 
.A(n_9434),
.Y(n_10119)
);

HB1xp67_ASAP7_75t_L g10120 ( 
.A(n_9644),
.Y(n_10120)
);

INVx1_ASAP7_75t_L g10121 ( 
.A(n_9634),
.Y(n_10121)
);

OAI22xp5_ASAP7_75t_SL g10122 ( 
.A1(n_9663),
.A2(n_6576),
.B1(n_6577),
.B2(n_6574),
.Y(n_10122)
);

BUFx6f_ASAP7_75t_L g10123 ( 
.A(n_9219),
.Y(n_10123)
);

INVx1_ASAP7_75t_L g10124 ( 
.A(n_9673),
.Y(n_10124)
);

INVx1_ASAP7_75t_L g10125 ( 
.A(n_9652),
.Y(n_10125)
);

NAND2xp33_ASAP7_75t_SL g10126 ( 
.A(n_9386),
.B(n_6579),
.Y(n_10126)
);

INVx1_ASAP7_75t_L g10127 ( 
.A(n_9655),
.Y(n_10127)
);

OAI22xp5_ASAP7_75t_SL g10128 ( 
.A1(n_9669),
.A2(n_6590),
.B1(n_6591),
.B2(n_6581),
.Y(n_10128)
);

INVx2_ASAP7_75t_L g10129 ( 
.A(n_9534),
.Y(n_10129)
);

HB1xp67_ASAP7_75t_L g10130 ( 
.A(n_9592),
.Y(n_10130)
);

INVx1_ASAP7_75t_L g10131 ( 
.A(n_9350),
.Y(n_10131)
);

AOI22xp5_ASAP7_75t_L g10132 ( 
.A1(n_9609),
.A2(n_6600),
.B1(n_6601),
.B2(n_6592),
.Y(n_10132)
);

AND2x4_ASAP7_75t_L g10133 ( 
.A(n_9406),
.B(n_6418),
.Y(n_10133)
);

NAND2xp5_ASAP7_75t_L g10134 ( 
.A(n_9588),
.B(n_6602),
.Y(n_10134)
);

INVx2_ASAP7_75t_L g10135 ( 
.A(n_9407),
.Y(n_10135)
);

BUFx6f_ASAP7_75t_L g10136 ( 
.A(n_9219),
.Y(n_10136)
);

BUFx6f_ASAP7_75t_L g10137 ( 
.A(n_9223),
.Y(n_10137)
);

INVx1_ASAP7_75t_L g10138 ( 
.A(n_9377),
.Y(n_10138)
);

INVx3_ASAP7_75t_L g10139 ( 
.A(n_9309),
.Y(n_10139)
);

CKINVDCx8_ASAP7_75t_R g10140 ( 
.A(n_9158),
.Y(n_10140)
);

INVx2_ASAP7_75t_L g10141 ( 
.A(n_9439),
.Y(n_10141)
);

INVx1_ASAP7_75t_L g10142 ( 
.A(n_9405),
.Y(n_10142)
);

INVx2_ASAP7_75t_L g10143 ( 
.A(n_9464),
.Y(n_10143)
);

INVx1_ASAP7_75t_L g10144 ( 
.A(n_9556),
.Y(n_10144)
);

AND2x2_ASAP7_75t_L g10145 ( 
.A(n_9615),
.B(n_6606),
.Y(n_10145)
);

INVx3_ASAP7_75t_L g10146 ( 
.A(n_9309),
.Y(n_10146)
);

INVx2_ASAP7_75t_L g10147 ( 
.A(n_9263),
.Y(n_10147)
);

INVx1_ASAP7_75t_L g10148 ( 
.A(n_9557),
.Y(n_10148)
);

BUFx6f_ASAP7_75t_L g10149 ( 
.A(n_9223),
.Y(n_10149)
);

INVx1_ASAP7_75t_L g10150 ( 
.A(n_9582),
.Y(n_10150)
);

CKINVDCx5p33_ASAP7_75t_R g10151 ( 
.A(n_9165),
.Y(n_10151)
);

OAI22xp5_ASAP7_75t_SL g10152 ( 
.A1(n_9672),
.A2(n_6610),
.B1(n_6616),
.B2(n_6607),
.Y(n_10152)
);

INVx1_ASAP7_75t_L g10153 ( 
.A(n_9637),
.Y(n_10153)
);

INVx2_ASAP7_75t_L g10154 ( 
.A(n_9247),
.Y(n_10154)
);

OAI22xp5_ASAP7_75t_L g10155 ( 
.A1(n_9616),
.A2(n_6619),
.B1(n_6625),
.B2(n_6618),
.Y(n_10155)
);

INVx2_ASAP7_75t_L g10156 ( 
.A(n_9247),
.Y(n_10156)
);

NAND2xp5_ASAP7_75t_L g10157 ( 
.A(n_9527),
.B(n_6626),
.Y(n_10157)
);

BUFx2_ASAP7_75t_L g10158 ( 
.A(n_9621),
.Y(n_10158)
);

INVx1_ASAP7_75t_L g10159 ( 
.A(n_9294),
.Y(n_10159)
);

INVxp67_ASAP7_75t_L g10160 ( 
.A(n_9408),
.Y(n_10160)
);

INVx1_ASAP7_75t_L g10161 ( 
.A(n_9295),
.Y(n_10161)
);

INVx2_ASAP7_75t_L g10162 ( 
.A(n_9260),
.Y(n_10162)
);

AND2x6_ASAP7_75t_L g10163 ( 
.A(n_9675),
.B(n_9478),
.Y(n_10163)
);

INVx1_ASAP7_75t_L g10164 ( 
.A(n_9299),
.Y(n_10164)
);

INVx2_ASAP7_75t_L g10165 ( 
.A(n_9260),
.Y(n_10165)
);

INVx2_ASAP7_75t_L g10166 ( 
.A(n_9343),
.Y(n_10166)
);

NAND2xp33_ASAP7_75t_SL g10167 ( 
.A(n_9551),
.B(n_6630),
.Y(n_10167)
);

OA21x2_ASAP7_75t_L g10168 ( 
.A1(n_9687),
.A2(n_6441),
.B(n_6420),
.Y(n_10168)
);

BUFx6f_ASAP7_75t_L g10169 ( 
.A(n_9147),
.Y(n_10169)
);

INVx1_ASAP7_75t_L g10170 ( 
.A(n_9653),
.Y(n_10170)
);

INVx2_ASAP7_75t_L g10171 ( 
.A(n_9394),
.Y(n_10171)
);

HB1xp67_ASAP7_75t_L g10172 ( 
.A(n_9385),
.Y(n_10172)
);

NAND2xp33_ASAP7_75t_SL g10173 ( 
.A(n_9598),
.B(n_6635),
.Y(n_10173)
);

CKINVDCx8_ASAP7_75t_R g10174 ( 
.A(n_9182),
.Y(n_10174)
);

INVx1_ASAP7_75t_L g10175 ( 
.A(n_9670),
.Y(n_10175)
);

AND2x2_ASAP7_75t_L g10176 ( 
.A(n_9643),
.B(n_6636),
.Y(n_10176)
);

AND2x4_ASAP7_75t_L g10177 ( 
.A(n_9147),
.B(n_6456),
.Y(n_10177)
);

INVxp67_ASAP7_75t_L g10178 ( 
.A(n_9308),
.Y(n_10178)
);

BUFx6f_ASAP7_75t_L g10179 ( 
.A(n_9149),
.Y(n_10179)
);

AND2x2_ASAP7_75t_L g10180 ( 
.A(n_9685),
.B(n_6644),
.Y(n_10180)
);

OAI22xp5_ASAP7_75t_SL g10181 ( 
.A1(n_9648),
.A2(n_9355),
.B1(n_9568),
.B2(n_9674),
.Y(n_10181)
);

AND2x4_ASAP7_75t_L g10182 ( 
.A(n_9149),
.B(n_6459),
.Y(n_10182)
);

INVx1_ASAP7_75t_L g10183 ( 
.A(n_9599),
.Y(n_10183)
);

INVx1_ASAP7_75t_L g10184 ( 
.A(n_9349),
.Y(n_10184)
);

NAND2xp5_ASAP7_75t_SL g10185 ( 
.A(n_9465),
.B(n_6646),
.Y(n_10185)
);

INVx1_ASAP7_75t_L g10186 ( 
.A(n_9357),
.Y(n_10186)
);

INVx2_ASAP7_75t_L g10187 ( 
.A(n_9683),
.Y(n_10187)
);

INVx1_ASAP7_75t_L g10188 ( 
.A(n_9443),
.Y(n_10188)
);

INVx2_ASAP7_75t_L g10189 ( 
.A(n_9683),
.Y(n_10189)
);

AOI22xp5_ASAP7_75t_L g10190 ( 
.A1(n_9425),
.A2(n_6658),
.B1(n_6660),
.B2(n_6650),
.Y(n_10190)
);

INVx2_ASAP7_75t_L g10191 ( 
.A(n_9675),
.Y(n_10191)
);

NAND3xp33_ASAP7_75t_SL g10192 ( 
.A(n_9624),
.B(n_6668),
.C(n_6664),
.Y(n_10192)
);

INVxp67_ASAP7_75t_L g10193 ( 
.A(n_9512),
.Y(n_10193)
);

INVx1_ASAP7_75t_L g10194 ( 
.A(n_9558),
.Y(n_10194)
);

INVx2_ASAP7_75t_L g10195 ( 
.A(n_9665),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_9562),
.Y(n_10196)
);

OA21x2_ASAP7_75t_L g10197 ( 
.A1(n_9145),
.A2(n_6465),
.B(n_6462),
.Y(n_10197)
);

INVx2_ASAP7_75t_L g10198 ( 
.A(n_9692),
.Y(n_10198)
);

INVx2_ASAP7_75t_L g10199 ( 
.A(n_9633),
.Y(n_10199)
);

INVx2_ASAP7_75t_L g10200 ( 
.A(n_9633),
.Y(n_10200)
);

INVx1_ASAP7_75t_L g10201 ( 
.A(n_9650),
.Y(n_10201)
);

INVxp67_ASAP7_75t_L g10202 ( 
.A(n_9222),
.Y(n_10202)
);

AND2x2_ASAP7_75t_L g10203 ( 
.A(n_9338),
.B(n_6669),
.Y(n_10203)
);

BUFx6f_ASAP7_75t_L g10204 ( 
.A(n_9650),
.Y(n_10204)
);

INVx2_ASAP7_75t_L g10205 ( 
.A(n_9255),
.Y(n_10205)
);

INVx1_ASAP7_75t_SL g10206 ( 
.A(n_9436),
.Y(n_10206)
);

INVx1_ASAP7_75t_L g10207 ( 
.A(n_9667),
.Y(n_10207)
);

INVx1_ASAP7_75t_L g10208 ( 
.A(n_9162),
.Y(n_10208)
);

AND2x6_ASAP7_75t_L g10209 ( 
.A(n_9353),
.B(n_6467),
.Y(n_10209)
);

INVx2_ASAP7_75t_L g10210 ( 
.A(n_9522),
.Y(n_10210)
);

BUFx6f_ASAP7_75t_L g10211 ( 
.A(n_9199),
.Y(n_10211)
);

OAI22xp5_ASAP7_75t_SL g10212 ( 
.A1(n_9429),
.A2(n_9440),
.B1(n_9233),
.B2(n_9285),
.Y(n_10212)
);

NAND2x1_ASAP7_75t_L g10213 ( 
.A(n_9522),
.B(n_9171),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_9522),
.Y(n_10214)
);

INVx1_ASAP7_75t_L g10215 ( 
.A(n_9586),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_9586),
.Y(n_10216)
);

OAI22xp5_ASAP7_75t_L g10217 ( 
.A1(n_9467),
.A2(n_6672),
.B1(n_6673),
.B2(n_6671),
.Y(n_10217)
);

AND2x6_ASAP7_75t_L g10218 ( 
.A(n_9356),
.B(n_6472),
.Y(n_10218)
);

INVx2_ASAP7_75t_L g10219 ( 
.A(n_9586),
.Y(n_10219)
);

NAND2xp5_ASAP7_75t_L g10220 ( 
.A(n_9505),
.B(n_6674),
.Y(n_10220)
);

INVx1_ASAP7_75t_L g10221 ( 
.A(n_9605),
.Y(n_10221)
);

BUFx2_ASAP7_75t_L g10222 ( 
.A(n_9181),
.Y(n_10222)
);

INVx1_ASAP7_75t_L g10223 ( 
.A(n_9360),
.Y(n_10223)
);

BUFx2_ASAP7_75t_L g10224 ( 
.A(n_9438),
.Y(n_10224)
);

INVx2_ASAP7_75t_L g10225 ( 
.A(n_9366),
.Y(n_10225)
);

INVx1_ASAP7_75t_L g10226 ( 
.A(n_9367),
.Y(n_10226)
);

INVx1_ASAP7_75t_L g10227 ( 
.A(n_9370),
.Y(n_10227)
);

INVx2_ASAP7_75t_L g10228 ( 
.A(n_9620),
.Y(n_10228)
);

INVx1_ASAP7_75t_L g10229 ( 
.A(n_9375),
.Y(n_10229)
);

BUFx2_ASAP7_75t_L g10230 ( 
.A(n_9320),
.Y(n_10230)
);

BUFx2_ASAP7_75t_L g10231 ( 
.A(n_9369),
.Y(n_10231)
);

INVx1_ASAP7_75t_L g10232 ( 
.A(n_9378),
.Y(n_10232)
);

HB1xp67_ASAP7_75t_L g10233 ( 
.A(n_9469),
.Y(n_10233)
);

AND3x1_ASAP7_75t_L g10234 ( 
.A(n_9341),
.B(n_6476),
.C(n_6475),
.Y(n_10234)
);

INVx1_ASAP7_75t_L g10235 ( 
.A(n_9640),
.Y(n_10235)
);

BUFx2_ASAP7_75t_L g10236 ( 
.A(n_9336),
.Y(n_10236)
);

INVx1_ASAP7_75t_L g10237 ( 
.A(n_9642),
.Y(n_10237)
);

INVx1_ASAP7_75t_L g10238 ( 
.A(n_9645),
.Y(n_10238)
);

INVx2_ASAP7_75t_L g10239 ( 
.A(n_9649),
.Y(n_10239)
);

INVx1_ASAP7_75t_L g10240 ( 
.A(n_9657),
.Y(n_10240)
);

NAND2xp5_ASAP7_75t_L g10241 ( 
.A(n_9191),
.B(n_6684),
.Y(n_10241)
);

NAND2xp5_ASAP7_75t_L g10242 ( 
.A(n_9211),
.B(n_6685),
.Y(n_10242)
);

INVx1_ASAP7_75t_L g10243 ( 
.A(n_9216),
.Y(n_10243)
);

HB1xp67_ASAP7_75t_L g10244 ( 
.A(n_9218),
.Y(n_10244)
);

AOI22xp5_ASAP7_75t_L g10245 ( 
.A1(n_9224),
.A2(n_6687),
.B1(n_6690),
.B2(n_6686),
.Y(n_10245)
);

INVx1_ASAP7_75t_L g10246 ( 
.A(n_9226),
.Y(n_10246)
);

NAND2xp33_ASAP7_75t_SL g10247 ( 
.A(n_9235),
.B(n_6691),
.Y(n_10247)
);

BUFx2_ASAP7_75t_L g10248 ( 
.A(n_9301),
.Y(n_10248)
);

INVx1_ASAP7_75t_L g10249 ( 
.A(n_9238),
.Y(n_10249)
);

INVx1_ASAP7_75t_L g10250 ( 
.A(n_9239),
.Y(n_10250)
);

BUFx6f_ASAP7_75t_L g10251 ( 
.A(n_9240),
.Y(n_10251)
);

INVx2_ASAP7_75t_L g10252 ( 
.A(n_9445),
.Y(n_10252)
);

AOI22xp5_ASAP7_75t_L g10253 ( 
.A1(n_9833),
.A2(n_9251),
.B1(n_9310),
.B2(n_9317),
.Y(n_10253)
);

INVx4_ASAP7_75t_L g10254 ( 
.A(n_10070),
.Y(n_10254)
);

INVx1_ASAP7_75t_L g10255 ( 
.A(n_9837),
.Y(n_10255)
);

INVx2_ASAP7_75t_L g10256 ( 
.A(n_9947),
.Y(n_10256)
);

BUFx2_ASAP7_75t_L g10257 ( 
.A(n_9710),
.Y(n_10257)
);

INVx1_ASAP7_75t_L g10258 ( 
.A(n_9844),
.Y(n_10258)
);

INVx4_ASAP7_75t_L g10259 ( 
.A(n_10070),
.Y(n_10259)
);

BUFx3_ASAP7_75t_L g10260 ( 
.A(n_9736),
.Y(n_10260)
);

NAND2xp5_ASAP7_75t_SL g10261 ( 
.A(n_9699),
.B(n_9453),
.Y(n_10261)
);

INVx1_ASAP7_75t_SL g10262 ( 
.A(n_9700),
.Y(n_10262)
);

CKINVDCx20_ASAP7_75t_R g10263 ( 
.A(n_9890),
.Y(n_10263)
);

BUFx4f_ASAP7_75t_L g10264 ( 
.A(n_10211),
.Y(n_10264)
);

NAND2xp5_ASAP7_75t_L g10265 ( 
.A(n_9826),
.B(n_6695),
.Y(n_10265)
);

NOR2xp33_ASAP7_75t_L g10266 ( 
.A(n_9814),
.B(n_9138),
.Y(n_10266)
);

BUFx3_ASAP7_75t_L g10267 ( 
.A(n_9736),
.Y(n_10267)
);

AND2x4_ASAP7_75t_L g10268 ( 
.A(n_9846),
.B(n_10050),
.Y(n_10268)
);

AND2x2_ASAP7_75t_L g10269 ( 
.A(n_9702),
.B(n_9256),
.Y(n_10269)
);

NAND2xp5_ASAP7_75t_L g10270 ( 
.A(n_9824),
.B(n_6703),
.Y(n_10270)
);

NAND2xp5_ASAP7_75t_L g10271 ( 
.A(n_9995),
.B(n_6704),
.Y(n_10271)
);

INVx1_ASAP7_75t_L g10272 ( 
.A(n_9701),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_9719),
.Y(n_10273)
);

BUFx3_ASAP7_75t_L g10274 ( 
.A(n_9847),
.Y(n_10274)
);

INVx1_ASAP7_75t_L g10275 ( 
.A(n_9721),
.Y(n_10275)
);

INVx2_ASAP7_75t_L g10276 ( 
.A(n_10000),
.Y(n_10276)
);

INVx2_ASAP7_75t_L g10277 ( 
.A(n_10008),
.Y(n_10277)
);

INVxp33_ASAP7_75t_SL g10278 ( 
.A(n_10212),
.Y(n_10278)
);

INVxp67_ASAP7_75t_SL g10279 ( 
.A(n_9723),
.Y(n_10279)
);

NAND2xp5_ASAP7_75t_L g10280 ( 
.A(n_9851),
.B(n_6706),
.Y(n_10280)
);

INVx1_ASAP7_75t_L g10281 ( 
.A(n_9726),
.Y(n_10281)
);

INVx3_ASAP7_75t_L g10282 ( 
.A(n_9740),
.Y(n_10282)
);

NAND2xp5_ASAP7_75t_L g10283 ( 
.A(n_9755),
.B(n_6708),
.Y(n_10283)
);

INVx1_ASAP7_75t_L g10284 ( 
.A(n_9729),
.Y(n_10284)
);

AND2x4_ASAP7_75t_L g10285 ( 
.A(n_10050),
.B(n_10204),
.Y(n_10285)
);

INVx1_ASAP7_75t_L g10286 ( 
.A(n_9731),
.Y(n_10286)
);

AND2x6_ASAP7_75t_L g10287 ( 
.A(n_9741),
.B(n_6478),
.Y(n_10287)
);

CKINVDCx5p33_ASAP7_75t_R g10288 ( 
.A(n_10151),
.Y(n_10288)
);

INVx3_ASAP7_75t_L g10289 ( 
.A(n_9740),
.Y(n_10289)
);

INVx2_ASAP7_75t_L g10290 ( 
.A(n_10015),
.Y(n_10290)
);

INVx4_ASAP7_75t_L g10291 ( 
.A(n_9742),
.Y(n_10291)
);

BUFx6f_ASAP7_75t_L g10292 ( 
.A(n_9742),
.Y(n_10292)
);

BUFx6f_ASAP7_75t_L g10293 ( 
.A(n_9752),
.Y(n_10293)
);

NOR2xp33_ASAP7_75t_L g10294 ( 
.A(n_10178),
.B(n_9143),
.Y(n_10294)
);

INVx3_ASAP7_75t_L g10295 ( 
.A(n_9759),
.Y(n_10295)
);

INVx4_ASAP7_75t_L g10296 ( 
.A(n_9752),
.Y(n_10296)
);

INVx2_ASAP7_75t_L g10297 ( 
.A(n_10019),
.Y(n_10297)
);

OAI22xp33_ASAP7_75t_L g10298 ( 
.A1(n_9919),
.A2(n_9261),
.B1(n_9265),
.B2(n_9264),
.Y(n_10298)
);

BUFx6f_ASAP7_75t_L g10299 ( 
.A(n_9759),
.Y(n_10299)
);

NAND2xp5_ASAP7_75t_SL g10300 ( 
.A(n_10083),
.B(n_9273),
.Y(n_10300)
);

AOI22xp33_ASAP7_75t_L g10301 ( 
.A1(n_10205),
.A2(n_6603),
.B1(n_6604),
.B2(n_6530),
.Y(n_10301)
);

INVxp67_ASAP7_75t_L g10302 ( 
.A(n_9720),
.Y(n_10302)
);

INVx2_ASAP7_75t_SL g10303 ( 
.A(n_9761),
.Y(n_10303)
);

NAND2xp5_ASAP7_75t_L g10304 ( 
.A(n_9769),
.B(n_6710),
.Y(n_10304)
);

BUFx3_ASAP7_75t_L g10305 ( 
.A(n_9847),
.Y(n_10305)
);

NAND2xp5_ASAP7_75t_SL g10306 ( 
.A(n_9735),
.B(n_9843),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_9734),
.Y(n_10307)
);

BUFx3_ASAP7_75t_L g10308 ( 
.A(n_9888),
.Y(n_10308)
);

INVx2_ASAP7_75t_L g10309 ( 
.A(n_10020),
.Y(n_10309)
);

INVx1_ASAP7_75t_L g10310 ( 
.A(n_9739),
.Y(n_10310)
);

INVx2_ASAP7_75t_SL g10311 ( 
.A(n_9761),
.Y(n_10311)
);

INVx3_ASAP7_75t_L g10312 ( 
.A(n_9829),
.Y(n_10312)
);

INVx1_ASAP7_75t_L g10313 ( 
.A(n_9746),
.Y(n_10313)
);

BUFx6f_ASAP7_75t_L g10314 ( 
.A(n_9829),
.Y(n_10314)
);

INVx1_ASAP7_75t_L g10315 ( 
.A(n_9754),
.Y(n_10315)
);

NAND2xp5_ASAP7_75t_L g10316 ( 
.A(n_9756),
.B(n_6711),
.Y(n_10316)
);

OAI22xp5_ASAP7_75t_L g10317 ( 
.A1(n_9737),
.A2(n_10001),
.B1(n_9987),
.B2(n_9992),
.Y(n_10317)
);

BUFx3_ASAP7_75t_L g10318 ( 
.A(n_9888),
.Y(n_10318)
);

AND2x4_ASAP7_75t_L g10319 ( 
.A(n_10204),
.B(n_9352),
.Y(n_10319)
);

AND2x4_ASAP7_75t_L g10320 ( 
.A(n_9935),
.B(n_9362),
.Y(n_10320)
);

INVx2_ASAP7_75t_L g10321 ( 
.A(n_9744),
.Y(n_10321)
);

INVx2_ASAP7_75t_L g10322 ( 
.A(n_9748),
.Y(n_10322)
);

INVx1_ASAP7_75t_L g10323 ( 
.A(n_9760),
.Y(n_10323)
);

INVx1_ASAP7_75t_SL g10324 ( 
.A(n_9765),
.Y(n_10324)
);

NOR3xp33_ASAP7_75t_L g10325 ( 
.A(n_9715),
.B(n_9627),
.C(n_9245),
.Y(n_10325)
);

BUFx4f_ASAP7_75t_L g10326 ( 
.A(n_10211),
.Y(n_10326)
);

INVx3_ASAP7_75t_R g10327 ( 
.A(n_10236),
.Y(n_10327)
);

NAND2xp5_ASAP7_75t_L g10328 ( 
.A(n_9762),
.B(n_6713),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_9764),
.Y(n_10329)
);

NAND2xp5_ASAP7_75t_SL g10330 ( 
.A(n_9895),
.B(n_9276),
.Y(n_10330)
);

NAND2xp5_ASAP7_75t_SL g10331 ( 
.A(n_10160),
.B(n_9277),
.Y(n_10331)
);

INVx6_ASAP7_75t_L g10332 ( 
.A(n_9697),
.Y(n_10332)
);

INVx1_ASAP7_75t_L g10333 ( 
.A(n_9766),
.Y(n_10333)
);

NAND2xp5_ASAP7_75t_SL g10334 ( 
.A(n_9708),
.B(n_9280),
.Y(n_10334)
);

INVx1_ASAP7_75t_L g10335 ( 
.A(n_9767),
.Y(n_10335)
);

AND2x4_ASAP7_75t_L g10336 ( 
.A(n_10199),
.B(n_9144),
.Y(n_10336)
);

INVx2_ASAP7_75t_L g10337 ( 
.A(n_9750),
.Y(n_10337)
);

CKINVDCx8_ASAP7_75t_R g10338 ( 
.A(n_9852),
.Y(n_10338)
);

OR2x2_ASAP7_75t_SL g10339 ( 
.A(n_10233),
.B(n_9437),
.Y(n_10339)
);

BUFx6f_ASAP7_75t_L g10340 ( 
.A(n_9838),
.Y(n_10340)
);

INVx2_ASAP7_75t_L g10341 ( 
.A(n_9751),
.Y(n_10341)
);

BUFx6f_ASAP7_75t_L g10342 ( 
.A(n_9838),
.Y(n_10342)
);

NAND2xp5_ASAP7_75t_L g10343 ( 
.A(n_9768),
.B(n_6714),
.Y(n_10343)
);

INVx1_ASAP7_75t_L g10344 ( 
.A(n_9770),
.Y(n_10344)
);

AND2x4_ASAP7_75t_L g10345 ( 
.A(n_10200),
.B(n_9286),
.Y(n_10345)
);

NAND2xp5_ASAP7_75t_L g10346 ( 
.A(n_9772),
.B(n_6715),
.Y(n_10346)
);

INVx1_ASAP7_75t_L g10347 ( 
.A(n_9776),
.Y(n_10347)
);

INVx2_ASAP7_75t_L g10348 ( 
.A(n_9753),
.Y(n_10348)
);

INVx2_ASAP7_75t_L g10349 ( 
.A(n_9758),
.Y(n_10349)
);

INVx1_ASAP7_75t_L g10350 ( 
.A(n_9777),
.Y(n_10350)
);

NAND2xp5_ASAP7_75t_SL g10351 ( 
.A(n_9874),
.B(n_9300),
.Y(n_10351)
);

INVx2_ASAP7_75t_L g10352 ( 
.A(n_9763),
.Y(n_10352)
);

NAND2xp5_ASAP7_75t_L g10353 ( 
.A(n_9780),
.B(n_6721),
.Y(n_10353)
);

INVx4_ASAP7_75t_L g10354 ( 
.A(n_9927),
.Y(n_10354)
);

INVx1_ASAP7_75t_L g10355 ( 
.A(n_9786),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_9787),
.Y(n_10356)
);

INVx3_ASAP7_75t_L g10357 ( 
.A(n_10169),
.Y(n_10357)
);

NOR2xp33_ASAP7_75t_L g10358 ( 
.A(n_9711),
.B(n_9307),
.Y(n_10358)
);

INVx1_ASAP7_75t_L g10359 ( 
.A(n_9794),
.Y(n_10359)
);

AND2x2_ASAP7_75t_L g10360 ( 
.A(n_9706),
.B(n_9441),
.Y(n_10360)
);

NAND2xp5_ASAP7_75t_L g10361 ( 
.A(n_9795),
.B(n_9796),
.Y(n_10361)
);

INVx2_ASAP7_75t_SL g10362 ( 
.A(n_9927),
.Y(n_10362)
);

INVx1_ASAP7_75t_L g10363 ( 
.A(n_9800),
.Y(n_10363)
);

AND2x2_ASAP7_75t_L g10364 ( 
.A(n_10176),
.B(n_9442),
.Y(n_10364)
);

INVx1_ASAP7_75t_L g10365 ( 
.A(n_9804),
.Y(n_10365)
);

INVx2_ASAP7_75t_L g10366 ( 
.A(n_9773),
.Y(n_10366)
);

NOR2xp33_ASAP7_75t_L g10367 ( 
.A(n_10014),
.B(n_9420),
.Y(n_10367)
);

INVx1_ASAP7_75t_L g10368 ( 
.A(n_9806),
.Y(n_10368)
);

NAND2xp5_ASAP7_75t_L g10369 ( 
.A(n_9812),
.B(n_9813),
.Y(n_10369)
);

OR2x2_ASAP7_75t_L g10370 ( 
.A(n_9821),
.B(n_6722),
.Y(n_10370)
);

NOR2xp33_ASAP7_75t_L g10371 ( 
.A(n_10018),
.B(n_6723),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_9816),
.Y(n_10372)
);

BUFx3_ASAP7_75t_L g10373 ( 
.A(n_9929),
.Y(n_10373)
);

AND2x2_ASAP7_75t_L g10374 ( 
.A(n_10180),
.B(n_6726),
.Y(n_10374)
);

BUFx4f_ASAP7_75t_L g10375 ( 
.A(n_9929),
.Y(n_10375)
);

NAND2xp5_ASAP7_75t_L g10376 ( 
.A(n_9819),
.B(n_6727),
.Y(n_10376)
);

INVx1_ASAP7_75t_L g10377 ( 
.A(n_9825),
.Y(n_10377)
);

NAND2xp5_ASAP7_75t_L g10378 ( 
.A(n_9827),
.B(n_9831),
.Y(n_10378)
);

INVx1_ASAP7_75t_L g10379 ( 
.A(n_9779),
.Y(n_10379)
);

INVx2_ASAP7_75t_L g10380 ( 
.A(n_9782),
.Y(n_10380)
);

INVx4_ASAP7_75t_L g10381 ( 
.A(n_9941),
.Y(n_10381)
);

AND2x4_ASAP7_75t_L g10382 ( 
.A(n_10052),
.B(n_9448),
.Y(n_10382)
);

OAI22xp5_ASAP7_75t_SL g10383 ( 
.A1(n_9705),
.A2(n_9460),
.B1(n_6730),
.B2(n_6733),
.Y(n_10383)
);

NAND2xp5_ASAP7_75t_SL g10384 ( 
.A(n_9802),
.B(n_6729),
.Y(n_10384)
);

AND2x4_ASAP7_75t_L g10385 ( 
.A(n_10049),
.B(n_6481),
.Y(n_10385)
);

INVx3_ASAP7_75t_L g10386 ( 
.A(n_10169),
.Y(n_10386)
);

NAND2xp5_ASAP7_75t_L g10387 ( 
.A(n_9784),
.B(n_6738),
.Y(n_10387)
);

NOR2xp33_ASAP7_75t_L g10388 ( 
.A(n_9707),
.B(n_6739),
.Y(n_10388)
);

INVx5_ASAP7_75t_L g10389 ( 
.A(n_10251),
.Y(n_10389)
);

AOI22xp5_ASAP7_75t_L g10390 ( 
.A1(n_9730),
.A2(n_6741),
.B1(n_6742),
.B2(n_6740),
.Y(n_10390)
);

AND2x4_ASAP7_75t_SL g10391 ( 
.A(n_10251),
.B(n_6487),
.Y(n_10391)
);

OR2x2_ASAP7_75t_L g10392 ( 
.A(n_9867),
.B(n_6747),
.Y(n_10392)
);

XOR2xp5_ASAP7_75t_SL g10393 ( 
.A(n_10244),
.B(n_6493),
.Y(n_10393)
);

INVx2_ASAP7_75t_L g10394 ( 
.A(n_9785),
.Y(n_10394)
);

OAI22xp5_ASAP7_75t_L g10395 ( 
.A1(n_9988),
.A2(n_6753),
.B1(n_6756),
.B2(n_6751),
.Y(n_10395)
);

CKINVDCx16_ASAP7_75t_R g10396 ( 
.A(n_10051),
.Y(n_10396)
);

AND2x6_ASAP7_75t_L g10397 ( 
.A(n_10243),
.B(n_6501),
.Y(n_10397)
);

INVxp33_ASAP7_75t_L g10398 ( 
.A(n_9703),
.Y(n_10398)
);

CKINVDCx20_ASAP7_75t_R g10399 ( 
.A(n_10038),
.Y(n_10399)
);

BUFx2_ASAP7_75t_L g10400 ( 
.A(n_9991),
.Y(n_10400)
);

OR2x6_ASAP7_75t_L g10401 ( 
.A(n_10179),
.B(n_6504),
.Y(n_10401)
);

BUFx3_ASAP7_75t_L g10402 ( 
.A(n_9941),
.Y(n_10402)
);

INVx2_ASAP7_75t_L g10403 ( 
.A(n_9791),
.Y(n_10403)
);

INVx2_ASAP7_75t_L g10404 ( 
.A(n_9792),
.Y(n_10404)
);

INVx1_ASAP7_75t_L g10405 ( 
.A(n_9797),
.Y(n_10405)
);

AND2x6_ASAP7_75t_L g10406 ( 
.A(n_10246),
.B(n_6518),
.Y(n_10406)
);

INVx3_ASAP7_75t_R g10407 ( 
.A(n_10158),
.Y(n_10407)
);

BUFx6f_ASAP7_75t_L g10408 ( 
.A(n_9950),
.Y(n_10408)
);

INVx1_ASAP7_75t_L g10409 ( 
.A(n_9798),
.Y(n_10409)
);

INVx1_ASAP7_75t_L g10410 ( 
.A(n_9807),
.Y(n_10410)
);

AND2x2_ASAP7_75t_L g10411 ( 
.A(n_10073),
.B(n_6760),
.Y(n_10411)
);

AOI22xp5_ASAP7_75t_L g10412 ( 
.A1(n_10005),
.A2(n_6762),
.B1(n_6763),
.B2(n_6761),
.Y(n_10412)
);

BUFx6f_ASAP7_75t_L g10413 ( 
.A(n_9950),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_9809),
.Y(n_10414)
);

INVx2_ASAP7_75t_SL g10415 ( 
.A(n_9964),
.Y(n_10415)
);

INVx4_ASAP7_75t_L g10416 ( 
.A(n_9964),
.Y(n_10416)
);

BUFx8_ASAP7_75t_SL g10417 ( 
.A(n_10231),
.Y(n_10417)
);

INVx3_ASAP7_75t_L g10418 ( 
.A(n_10179),
.Y(n_10418)
);

NOR2xp33_ASAP7_75t_R g10419 ( 
.A(n_9928),
.B(n_6766),
.Y(n_10419)
);

OR2x2_ASAP7_75t_L g10420 ( 
.A(n_9887),
.B(n_6767),
.Y(n_10420)
);

INVx1_ASAP7_75t_L g10421 ( 
.A(n_9815),
.Y(n_10421)
);

INVx4_ASAP7_75t_L g10422 ( 
.A(n_9986),
.Y(n_10422)
);

NAND2xp5_ASAP7_75t_SL g10423 ( 
.A(n_9704),
.B(n_6768),
.Y(n_10423)
);

INVx1_ASAP7_75t_SL g10424 ( 
.A(n_9839),
.Y(n_10424)
);

NAND2xp5_ASAP7_75t_L g10425 ( 
.A(n_9818),
.B(n_6772),
.Y(n_10425)
);

NOR2xp33_ASAP7_75t_L g10426 ( 
.A(n_10114),
.B(n_6773),
.Y(n_10426)
);

INVx2_ASAP7_75t_L g10427 ( 
.A(n_9830),
.Y(n_10427)
);

NAND3xp33_ASAP7_75t_L g10428 ( 
.A(n_9994),
.B(n_6775),
.C(n_6774),
.Y(n_10428)
);

AOI22xp33_ASAP7_75t_L g10429 ( 
.A1(n_10207),
.A2(n_6675),
.B1(n_6678),
.B2(n_6608),
.Y(n_10429)
);

BUFx6f_ASAP7_75t_L g10430 ( 
.A(n_9986),
.Y(n_10430)
);

AO21x2_ASAP7_75t_L g10431 ( 
.A1(n_9832),
.A2(n_6520),
.B(n_6519),
.Y(n_10431)
);

INVx4_ASAP7_75t_SL g10432 ( 
.A(n_10209),
.Y(n_10432)
);

INVx5_ASAP7_75t_L g10433 ( 
.A(n_9990),
.Y(n_10433)
);

AND2x4_ASAP7_75t_L g10434 ( 
.A(n_9781),
.B(n_6533),
.Y(n_10434)
);

BUFx6f_ASAP7_75t_L g10435 ( 
.A(n_9990),
.Y(n_10435)
);

INVx2_ASAP7_75t_L g10436 ( 
.A(n_10029),
.Y(n_10436)
);

INVx5_ASAP7_75t_L g10437 ( 
.A(n_9999),
.Y(n_10437)
);

NAND2xp5_ASAP7_75t_SL g10438 ( 
.A(n_9757),
.B(n_6779),
.Y(n_10438)
);

OAI22xp5_ASAP7_75t_L g10439 ( 
.A1(n_10011),
.A2(n_6783),
.B1(n_6785),
.B2(n_6782),
.Y(n_10439)
);

INVx4_ASAP7_75t_L g10440 ( 
.A(n_9999),
.Y(n_10440)
);

INVx2_ASAP7_75t_L g10441 ( 
.A(n_10041),
.Y(n_10441)
);

INVx2_ASAP7_75t_L g10442 ( 
.A(n_10044),
.Y(n_10442)
);

INVx2_ASAP7_75t_L g10443 ( 
.A(n_10054),
.Y(n_10443)
);

NAND2xp5_ASAP7_75t_L g10444 ( 
.A(n_9808),
.B(n_6790),
.Y(n_10444)
);

OR2x2_ASAP7_75t_L g10445 ( 
.A(n_9810),
.B(n_9840),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_10118),
.B(n_6798),
.Y(n_10446)
);

INVx4_ASAP7_75t_L g10447 ( 
.A(n_10031),
.Y(n_10447)
);

INVx1_ASAP7_75t_L g10448 ( 
.A(n_9855),
.Y(n_10448)
);

BUFx2_ASAP7_75t_L g10449 ( 
.A(n_10031),
.Y(n_10449)
);

NAND2xp5_ASAP7_75t_L g10450 ( 
.A(n_9783),
.B(n_6799),
.Y(n_10450)
);

INVx1_ASAP7_75t_L g10451 ( 
.A(n_9856),
.Y(n_10451)
);

NAND3xp33_ASAP7_75t_L g10452 ( 
.A(n_10034),
.B(n_6806),
.C(n_6804),
.Y(n_10452)
);

INVx1_ASAP7_75t_L g10453 ( 
.A(n_9860),
.Y(n_10453)
);

INVx2_ASAP7_75t_L g10454 ( 
.A(n_10055),
.Y(n_10454)
);

INVx3_ASAP7_75t_L g10455 ( 
.A(n_10108),
.Y(n_10455)
);

NAND2xp5_ASAP7_75t_SL g10456 ( 
.A(n_9790),
.B(n_6810),
.Y(n_10456)
);

INVx2_ASAP7_75t_L g10457 ( 
.A(n_10063),
.Y(n_10457)
);

INVxp67_ASAP7_75t_L g10458 ( 
.A(n_9993),
.Y(n_10458)
);

INVx2_ASAP7_75t_L g10459 ( 
.A(n_9698),
.Y(n_10459)
);

INVx2_ASAP7_75t_L g10460 ( 
.A(n_9712),
.Y(n_10460)
);

INVx1_ASAP7_75t_L g10461 ( 
.A(n_9861),
.Y(n_10461)
);

OR2x2_ASAP7_75t_L g10462 ( 
.A(n_10228),
.B(n_6811),
.Y(n_10462)
);

INVx1_ASAP7_75t_L g10463 ( 
.A(n_9864),
.Y(n_10463)
);

AND2x2_ASAP7_75t_L g10464 ( 
.A(n_10145),
.B(n_6814),
.Y(n_10464)
);

NAND2xp5_ASAP7_75t_L g10465 ( 
.A(n_9783),
.B(n_6816),
.Y(n_10465)
);

INVx1_ASAP7_75t_SL g10466 ( 
.A(n_10035),
.Y(n_10466)
);

AND2x2_ASAP7_75t_L g10467 ( 
.A(n_9749),
.B(n_9801),
.Y(n_10467)
);

OR2x2_ASAP7_75t_L g10468 ( 
.A(n_10248),
.B(n_6820),
.Y(n_10468)
);

INVx1_ASAP7_75t_L g10469 ( 
.A(n_9865),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_L g10470 ( 
.A(n_9783),
.B(n_6822),
.Y(n_10470)
);

AND2x2_ASAP7_75t_L g10471 ( 
.A(n_9841),
.B(n_6823),
.Y(n_10471)
);

BUFx6f_ASAP7_75t_L g10472 ( 
.A(n_10046),
.Y(n_10472)
);

NAND2xp5_ASAP7_75t_SL g10473 ( 
.A(n_10091),
.B(n_6828),
.Y(n_10473)
);

INVx2_ASAP7_75t_L g10474 ( 
.A(n_9713),
.Y(n_10474)
);

OAI22xp33_ASAP7_75t_L g10475 ( 
.A1(n_9892),
.A2(n_6831),
.B1(n_6832),
.B2(n_6829),
.Y(n_10475)
);

AND2x4_ASAP7_75t_L g10476 ( 
.A(n_9789),
.B(n_6536),
.Y(n_10476)
);

INVxp67_ASAP7_75t_L g10477 ( 
.A(n_10056),
.Y(n_10477)
);

INVx3_ASAP7_75t_L g10478 ( 
.A(n_10140),
.Y(n_10478)
);

NAND2xp5_ASAP7_75t_SL g10479 ( 
.A(n_9933),
.B(n_6840),
.Y(n_10479)
);

INVx1_ASAP7_75t_L g10480 ( 
.A(n_9869),
.Y(n_10480)
);

BUFx2_ASAP7_75t_L g10481 ( 
.A(n_10046),
.Y(n_10481)
);

INVx1_ASAP7_75t_L g10482 ( 
.A(n_9873),
.Y(n_10482)
);

BUFx10_ASAP7_75t_L g10483 ( 
.A(n_9842),
.Y(n_10483)
);

INVx1_ASAP7_75t_L g10484 ( 
.A(n_9875),
.Y(n_10484)
);

INVx1_ASAP7_75t_L g10485 ( 
.A(n_9876),
.Y(n_10485)
);

NAND2xp5_ASAP7_75t_SL g10486 ( 
.A(n_10226),
.B(n_6841),
.Y(n_10486)
);

INVxp67_ASAP7_75t_SL g10487 ( 
.A(n_10123),
.Y(n_10487)
);

AND2x2_ASAP7_75t_L g10488 ( 
.A(n_9866),
.B(n_6843),
.Y(n_10488)
);

BUFx6f_ASAP7_75t_L g10489 ( 
.A(n_10123),
.Y(n_10489)
);

OR2x2_ASAP7_75t_L g10490 ( 
.A(n_10002),
.B(n_6844),
.Y(n_10490)
);

OAI22xp33_ASAP7_75t_L g10491 ( 
.A1(n_10124),
.A2(n_6846),
.B1(n_6848),
.B2(n_6845),
.Y(n_10491)
);

NOR2xp33_ASAP7_75t_L g10492 ( 
.A(n_10241),
.B(n_6849),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_9877),
.Y(n_10493)
);

NOR2xp33_ASAP7_75t_L g10494 ( 
.A(n_10242),
.B(n_6851),
.Y(n_10494)
);

NAND2xp5_ASAP7_75t_L g10495 ( 
.A(n_9774),
.B(n_6854),
.Y(n_10495)
);

INVx2_ASAP7_75t_L g10496 ( 
.A(n_9714),
.Y(n_10496)
);

CKINVDCx5p33_ASAP7_75t_R g10497 ( 
.A(n_10174),
.Y(n_10497)
);

BUFx6f_ASAP7_75t_L g10498 ( 
.A(n_10136),
.Y(n_10498)
);

NAND2xp5_ASAP7_75t_L g10499 ( 
.A(n_9817),
.B(n_9908),
.Y(n_10499)
);

INVx1_ASAP7_75t_L g10500 ( 
.A(n_9880),
.Y(n_10500)
);

CKINVDCx20_ASAP7_75t_R g10501 ( 
.A(n_10222),
.Y(n_10501)
);

INVx1_ASAP7_75t_L g10502 ( 
.A(n_9882),
.Y(n_10502)
);

NAND2xp5_ASAP7_75t_SL g10503 ( 
.A(n_10227),
.B(n_6855),
.Y(n_10503)
);

NAND2xp5_ASAP7_75t_L g10504 ( 
.A(n_9913),
.B(n_6866),
.Y(n_10504)
);

INVx2_ASAP7_75t_L g10505 ( 
.A(n_9716),
.Y(n_10505)
);

INVx2_ASAP7_75t_L g10506 ( 
.A(n_9717),
.Y(n_10506)
);

NOR2xp33_ASAP7_75t_L g10507 ( 
.A(n_9868),
.B(n_6867),
.Y(n_10507)
);

AND2x4_ASAP7_75t_L g10508 ( 
.A(n_9811),
.B(n_6555),
.Y(n_10508)
);

AND2x2_ASAP7_75t_L g10509 ( 
.A(n_10023),
.B(n_6869),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9884),
.Y(n_10510)
);

INVx1_ASAP7_75t_L g10511 ( 
.A(n_9889),
.Y(n_10511)
);

NAND2xp33_ASAP7_75t_L g10512 ( 
.A(n_10163),
.B(n_6872),
.Y(n_10512)
);

NOR2xp33_ASAP7_75t_L g10513 ( 
.A(n_10229),
.B(n_6873),
.Y(n_10513)
);

AOI22xp33_ASAP7_75t_L g10514 ( 
.A1(n_9738),
.A2(n_6716),
.B1(n_6749),
.B2(n_6680),
.Y(n_10514)
);

AND2x4_ASAP7_75t_L g10515 ( 
.A(n_9907),
.B(n_6556),
.Y(n_10515)
);

INVx5_ASAP7_75t_L g10516 ( 
.A(n_10136),
.Y(n_10516)
);

BUFx10_ASAP7_75t_L g10517 ( 
.A(n_9870),
.Y(n_10517)
);

NOR2xp33_ASAP7_75t_L g10518 ( 
.A(n_10232),
.B(n_6875),
.Y(n_10518)
);

NAND2xp5_ASAP7_75t_L g10519 ( 
.A(n_9916),
.B(n_6876),
.Y(n_10519)
);

INVx1_ASAP7_75t_SL g10520 ( 
.A(n_10092),
.Y(n_10520)
);

HB1xp67_ASAP7_75t_L g10521 ( 
.A(n_10130),
.Y(n_10521)
);

NAND2xp5_ASAP7_75t_SL g10522 ( 
.A(n_10249),
.B(n_6878),
.Y(n_10522)
);

INVx1_ASAP7_75t_L g10523 ( 
.A(n_9894),
.Y(n_10523)
);

AND2x2_ASAP7_75t_L g10524 ( 
.A(n_9952),
.B(n_6882),
.Y(n_10524)
);

INVx2_ASAP7_75t_L g10525 ( 
.A(n_9727),
.Y(n_10525)
);

INVx1_ASAP7_75t_L g10526 ( 
.A(n_9896),
.Y(n_10526)
);

BUFx6f_ASAP7_75t_L g10527 ( 
.A(n_10137),
.Y(n_10527)
);

INVx5_ASAP7_75t_L g10528 ( 
.A(n_10137),
.Y(n_10528)
);

NOR2xp33_ASAP7_75t_L g10529 ( 
.A(n_9745),
.B(n_6884),
.Y(n_10529)
);

INVx6_ASAP7_75t_L g10530 ( 
.A(n_9697),
.Y(n_10530)
);

INVx2_ASAP7_75t_SL g10531 ( 
.A(n_10149),
.Y(n_10531)
);

INVx2_ASAP7_75t_L g10532 ( 
.A(n_9728),
.Y(n_10532)
);

AND2x2_ASAP7_75t_L g10533 ( 
.A(n_9979),
.B(n_6885),
.Y(n_10533)
);

NAND2xp5_ASAP7_75t_L g10534 ( 
.A(n_9955),
.B(n_6886),
.Y(n_10534)
);

NAND2xp5_ASAP7_75t_L g10535 ( 
.A(n_9850),
.B(n_9854),
.Y(n_10535)
);

AO21x2_ASAP7_75t_L g10536 ( 
.A1(n_10166),
.A2(n_10171),
.B(n_10147),
.Y(n_10536)
);

NOR2x1p5_ASAP7_75t_L g10537 ( 
.A(n_10225),
.B(n_6894),
.Y(n_10537)
);

OAI22xp5_ASAP7_75t_SL g10538 ( 
.A1(n_9709),
.A2(n_9922),
.B1(n_10181),
.B2(n_10066),
.Y(n_10538)
);

NAND2xp5_ASAP7_75t_SL g10539 ( 
.A(n_10250),
.B(n_6896),
.Y(n_10539)
);

BUFx6f_ASAP7_75t_L g10540 ( 
.A(n_10149),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_9898),
.Y(n_10541)
);

INVx4_ASAP7_75t_L g10542 ( 
.A(n_9722),
.Y(n_10542)
);

INVx4_ASAP7_75t_L g10543 ( 
.A(n_9722),
.Y(n_10543)
);

BUFx3_ASAP7_75t_L g10544 ( 
.A(n_9912),
.Y(n_10544)
);

NAND2xp5_ASAP7_75t_L g10545 ( 
.A(n_10012),
.B(n_6898),
.Y(n_10545)
);

NOR2xp33_ASAP7_75t_L g10546 ( 
.A(n_9863),
.B(n_10193),
.Y(n_10546)
);

INVx2_ASAP7_75t_L g10547 ( 
.A(n_9733),
.Y(n_10547)
);

AND2x2_ASAP7_75t_L g10548 ( 
.A(n_9951),
.B(n_6903),
.Y(n_10548)
);

INVx4_ASAP7_75t_SL g10549 ( 
.A(n_10209),
.Y(n_10549)
);

NOR2xp33_ASAP7_75t_L g10550 ( 
.A(n_10112),
.B(n_9820),
.Y(n_10550)
);

BUFx6f_ASAP7_75t_L g10551 ( 
.A(n_9926),
.Y(n_10551)
);

AND3x4_ASAP7_75t_L g10552 ( 
.A(n_10048),
.B(n_6777),
.C(n_6759),
.Y(n_10552)
);

HB1xp67_ASAP7_75t_L g10553 ( 
.A(n_10120),
.Y(n_10553)
);

NAND2xp5_ASAP7_75t_SL g10554 ( 
.A(n_9718),
.B(n_6904),
.Y(n_10554)
);

INVx6_ASAP7_75t_L g10555 ( 
.A(n_10085),
.Y(n_10555)
);

OR2x6_ASAP7_75t_L g10556 ( 
.A(n_10172),
.B(n_6559),
.Y(n_10556)
);

INVx1_ASAP7_75t_L g10557 ( 
.A(n_9902),
.Y(n_10557)
);

AND2x2_ASAP7_75t_L g10558 ( 
.A(n_9934),
.B(n_6905),
.Y(n_10558)
);

AND2x6_ASAP7_75t_L g10559 ( 
.A(n_10235),
.B(n_6562),
.Y(n_10559)
);

BUFx6f_ASAP7_75t_L g10560 ( 
.A(n_9931),
.Y(n_10560)
);

BUFx3_ASAP7_75t_L g10561 ( 
.A(n_9949),
.Y(n_10561)
);

INVx1_ASAP7_75t_L g10562 ( 
.A(n_9904),
.Y(n_10562)
);

INVx2_ASAP7_75t_L g10563 ( 
.A(n_9743),
.Y(n_10563)
);

INVx1_ASAP7_75t_L g10564 ( 
.A(n_9905),
.Y(n_10564)
);

BUFx3_ASAP7_75t_L g10565 ( 
.A(n_10006),
.Y(n_10565)
);

AND2x2_ASAP7_75t_L g10566 ( 
.A(n_10103),
.B(n_6906),
.Y(n_10566)
);

INVx1_ASAP7_75t_L g10567 ( 
.A(n_9910),
.Y(n_10567)
);

OR2x6_ASAP7_75t_L g10568 ( 
.A(n_10223),
.B(n_6565),
.Y(n_10568)
);

AOI22xp33_ASAP7_75t_L g10569 ( 
.A1(n_9893),
.A2(n_6827),
.B1(n_6842),
.B2(n_6815),
.Y(n_10569)
);

BUFx6f_ASAP7_75t_L g10570 ( 
.A(n_10024),
.Y(n_10570)
);

AND2x6_ASAP7_75t_L g10571 ( 
.A(n_10237),
.B(n_6566),
.Y(n_10571)
);

AND2x2_ASAP7_75t_L g10572 ( 
.A(n_10203),
.B(n_9996),
.Y(n_10572)
);

NOR2xp33_ASAP7_75t_L g10573 ( 
.A(n_9823),
.B(n_6909),
.Y(n_10573)
);

INVx4_ASAP7_75t_L g10574 ( 
.A(n_10027),
.Y(n_10574)
);

AND2x2_ASAP7_75t_L g10575 ( 
.A(n_9997),
.B(n_6910),
.Y(n_10575)
);

INVx1_ASAP7_75t_L g10576 ( 
.A(n_9914),
.Y(n_10576)
);

NAND2xp5_ASAP7_75t_L g10577 ( 
.A(n_10013),
.B(n_6914),
.Y(n_10577)
);

INVx4_ASAP7_75t_L g10578 ( 
.A(n_10037),
.Y(n_10578)
);

CKINVDCx5p33_ASAP7_75t_R g10579 ( 
.A(n_10119),
.Y(n_10579)
);

INVx2_ASAP7_75t_L g10580 ( 
.A(n_9822),
.Y(n_10580)
);

INVxp67_ASAP7_75t_L g10581 ( 
.A(n_10221),
.Y(n_10581)
);

BUFx2_ASAP7_75t_L g10582 ( 
.A(n_10080),
.Y(n_10582)
);

NAND2xp5_ASAP7_75t_SL g10583 ( 
.A(n_9967),
.B(n_6916),
.Y(n_10583)
);

NAND2xp5_ASAP7_75t_L g10584 ( 
.A(n_10017),
.B(n_6917),
.Y(n_10584)
);

INVx1_ASAP7_75t_L g10585 ( 
.A(n_9917),
.Y(n_10585)
);

INVx2_ASAP7_75t_L g10586 ( 
.A(n_9835),
.Y(n_10586)
);

INVx1_ASAP7_75t_L g10587 ( 
.A(n_9923),
.Y(n_10587)
);

NAND2xp5_ASAP7_75t_L g10588 ( 
.A(n_10016),
.B(n_6918),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_9845),
.Y(n_10589)
);

AND2x2_ASAP7_75t_L g10590 ( 
.A(n_10177),
.B(n_6919),
.Y(n_10590)
);

BUFx3_ASAP7_75t_L g10591 ( 
.A(n_10062),
.Y(n_10591)
);

INVx1_ASAP7_75t_L g10592 ( 
.A(n_9924),
.Y(n_10592)
);

NAND2xp33_ASAP7_75t_L g10593 ( 
.A(n_10163),
.B(n_6922),
.Y(n_10593)
);

INVx1_ASAP7_75t_L g10594 ( 
.A(n_9930),
.Y(n_10594)
);

INVx2_ASAP7_75t_SL g10595 ( 
.A(n_10154),
.Y(n_10595)
);

BUFx6f_ASAP7_75t_L g10596 ( 
.A(n_10084),
.Y(n_10596)
);

INVx1_ASAP7_75t_SL g10597 ( 
.A(n_10206),
.Y(n_10597)
);

AND2x2_ASAP7_75t_L g10598 ( 
.A(n_10182),
.B(n_6927),
.Y(n_10598)
);

BUFx3_ASAP7_75t_L g10599 ( 
.A(n_10139),
.Y(n_10599)
);

INVx2_ASAP7_75t_L g10600 ( 
.A(n_9848),
.Y(n_10600)
);

INVx1_ASAP7_75t_L g10601 ( 
.A(n_9932),
.Y(n_10601)
);

INVx1_ASAP7_75t_L g10602 ( 
.A(n_9938),
.Y(n_10602)
);

INVx2_ASAP7_75t_L g10603 ( 
.A(n_9853),
.Y(n_10603)
);

INVx1_ASAP7_75t_L g10604 ( 
.A(n_9939),
.Y(n_10604)
);

INVx2_ASAP7_75t_SL g10605 ( 
.A(n_10156),
.Y(n_10605)
);

INVx2_ASAP7_75t_L g10606 ( 
.A(n_9858),
.Y(n_10606)
);

INVx2_ASAP7_75t_L g10607 ( 
.A(n_9859),
.Y(n_10607)
);

INVx3_ASAP7_75t_L g10608 ( 
.A(n_10146),
.Y(n_10608)
);

INVx1_ASAP7_75t_L g10609 ( 
.A(n_9943),
.Y(n_10609)
);

OR2x2_ASAP7_75t_SL g10610 ( 
.A(n_10192),
.B(n_6571),
.Y(n_10610)
);

NOR2xp33_ASAP7_75t_L g10611 ( 
.A(n_9849),
.B(n_6932),
.Y(n_10611)
);

BUFx6f_ASAP7_75t_L g10612 ( 
.A(n_10162),
.Y(n_10612)
);

BUFx6f_ASAP7_75t_L g10613 ( 
.A(n_10165),
.Y(n_10613)
);

INVx2_ASAP7_75t_L g10614 ( 
.A(n_9871),
.Y(n_10614)
);

INVx5_ASAP7_75t_L g10615 ( 
.A(n_10209),
.Y(n_10615)
);

AOI22xp33_ASAP7_75t_L g10616 ( 
.A1(n_10194),
.A2(n_6907),
.B1(n_6935),
.B2(n_6879),
.Y(n_10616)
);

INVx2_ASAP7_75t_L g10617 ( 
.A(n_9872),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_10022),
.Y(n_10618)
);

BUFx3_ASAP7_75t_L g10619 ( 
.A(n_10111),
.Y(n_10619)
);

INVx3_ASAP7_75t_L g10620 ( 
.A(n_10117),
.Y(n_10620)
);

INVx2_ASAP7_75t_L g10621 ( 
.A(n_9878),
.Y(n_10621)
);

OR2x2_ASAP7_75t_SL g10622 ( 
.A(n_9879),
.B(n_6575),
.Y(n_10622)
);

NAND2xp5_ASAP7_75t_L g10623 ( 
.A(n_9942),
.B(n_6934),
.Y(n_10623)
);

INVx1_ASAP7_75t_L g10624 ( 
.A(n_10025),
.Y(n_10624)
);

AND2x2_ASAP7_75t_L g10625 ( 
.A(n_9883),
.B(n_6938),
.Y(n_10625)
);

NOR2xp33_ASAP7_75t_L g10626 ( 
.A(n_9936),
.B(n_6942),
.Y(n_10626)
);

INVx2_ASAP7_75t_L g10627 ( 
.A(n_9885),
.Y(n_10627)
);

INVx2_ASAP7_75t_SL g10628 ( 
.A(n_10129),
.Y(n_10628)
);

NOR2xp33_ASAP7_75t_L g10629 ( 
.A(n_9948),
.B(n_6944),
.Y(n_10629)
);

BUFx6f_ASAP7_75t_L g10630 ( 
.A(n_10042),
.Y(n_10630)
);

NAND2xp5_ASAP7_75t_L g10631 ( 
.A(n_10196),
.B(n_6951),
.Y(n_10631)
);

NAND2xp5_ASAP7_75t_L g10632 ( 
.A(n_9886),
.B(n_6955),
.Y(n_10632)
);

INVx2_ASAP7_75t_L g10633 ( 
.A(n_9891),
.Y(n_10633)
);

INVx1_ASAP7_75t_L g10634 ( 
.A(n_10030),
.Y(n_10634)
);

NOR2xp33_ASAP7_75t_L g10635 ( 
.A(n_9998),
.B(n_6958),
.Y(n_10635)
);

BUFx6f_ASAP7_75t_L g10636 ( 
.A(n_9778),
.Y(n_10636)
);

NAND2xp5_ASAP7_75t_L g10637 ( 
.A(n_9897),
.B(n_6961),
.Y(n_10637)
);

INVx1_ASAP7_75t_L g10638 ( 
.A(n_10032),
.Y(n_10638)
);

INVx2_ASAP7_75t_L g10639 ( 
.A(n_9900),
.Y(n_10639)
);

AND2x2_ASAP7_75t_SL g10640 ( 
.A(n_10230),
.B(n_6964),
.Y(n_10640)
);

INVx3_ASAP7_75t_L g10641 ( 
.A(n_10135),
.Y(n_10641)
);

NAND2xp5_ASAP7_75t_L g10642 ( 
.A(n_9903),
.B(n_6962),
.Y(n_10642)
);

OR2x2_ASAP7_75t_L g10643 ( 
.A(n_10239),
.B(n_6967),
.Y(n_10643)
);

INVx2_ASAP7_75t_SL g10644 ( 
.A(n_9921),
.Y(n_10644)
);

INVx1_ASAP7_75t_L g10645 ( 
.A(n_10045),
.Y(n_10645)
);

AND2x2_ASAP7_75t_SL g10646 ( 
.A(n_10224),
.B(n_7036),
.Y(n_10646)
);

NOR2xp33_ASAP7_75t_L g10647 ( 
.A(n_10010),
.B(n_6969),
.Y(n_10647)
);

AND2x6_ASAP7_75t_L g10648 ( 
.A(n_10238),
.B(n_6578),
.Y(n_10648)
);

NOR2xp33_ASAP7_75t_L g10649 ( 
.A(n_9788),
.B(n_6970),
.Y(n_10649)
);

AND2x6_ASAP7_75t_L g10650 ( 
.A(n_10240),
.B(n_6582),
.Y(n_10650)
);

BUFx6f_ASAP7_75t_L g10651 ( 
.A(n_10067),
.Y(n_10651)
);

INVx2_ASAP7_75t_L g10652 ( 
.A(n_9906),
.Y(n_10652)
);

INVx1_ASAP7_75t_L g10653 ( 
.A(n_10047),
.Y(n_10653)
);

INVx2_ASAP7_75t_L g10654 ( 
.A(n_9915),
.Y(n_10654)
);

NAND2xp5_ASAP7_75t_L g10655 ( 
.A(n_9918),
.B(n_6978),
.Y(n_10655)
);

INVx2_ASAP7_75t_L g10656 ( 
.A(n_9920),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_9937),
.Y(n_10657)
);

AND2x2_ASAP7_75t_L g10658 ( 
.A(n_10110),
.B(n_6981),
.Y(n_10658)
);

INVx1_ASAP7_75t_L g10659 ( 
.A(n_9940),
.Y(n_10659)
);

INVx1_ASAP7_75t_L g10660 ( 
.A(n_9944),
.Y(n_10660)
);

NOR2xp33_ASAP7_75t_L g10661 ( 
.A(n_9793),
.B(n_6982),
.Y(n_10661)
);

OA22x2_ASAP7_75t_L g10662 ( 
.A1(n_9724),
.A2(n_6986),
.B1(n_6987),
.B2(n_6983),
.Y(n_10662)
);

OAI22xp33_ASAP7_75t_L g10663 ( 
.A1(n_9911),
.A2(n_6989),
.B1(n_6991),
.B2(n_6988),
.Y(n_10663)
);

INVx2_ASAP7_75t_L g10664 ( 
.A(n_9958),
.Y(n_10664)
);

BUFx6f_ASAP7_75t_L g10665 ( 
.A(n_10077),
.Y(n_10665)
);

NOR2xp33_ASAP7_75t_L g10666 ( 
.A(n_9775),
.B(n_6992),
.Y(n_10666)
);

NAND2xp5_ASAP7_75t_L g10667 ( 
.A(n_9901),
.B(n_6994),
.Y(n_10667)
);

NAND2xp5_ASAP7_75t_SL g10668 ( 
.A(n_9971),
.B(n_10040),
.Y(n_10668)
);

BUFx3_ASAP7_75t_L g10669 ( 
.A(n_10201),
.Y(n_10669)
);

INVx1_ASAP7_75t_L g10670 ( 
.A(n_9946),
.Y(n_10670)
);

AND2x2_ASAP7_75t_L g10671 ( 
.A(n_10115),
.B(n_6996),
.Y(n_10671)
);

INVx2_ASAP7_75t_L g10672 ( 
.A(n_9959),
.Y(n_10672)
);

AND2x4_ASAP7_75t_L g10673 ( 
.A(n_10107),
.B(n_6585),
.Y(n_10673)
);

INVx2_ASAP7_75t_L g10674 ( 
.A(n_9953),
.Y(n_10674)
);

INVx4_ASAP7_75t_L g10675 ( 
.A(n_10163),
.Y(n_10675)
);

NAND2xp5_ASAP7_75t_L g10676 ( 
.A(n_9961),
.B(n_6997),
.Y(n_10676)
);

NAND2xp5_ASAP7_75t_L g10677 ( 
.A(n_9965),
.B(n_7002),
.Y(n_10677)
);

NOR2xp33_ASAP7_75t_L g10678 ( 
.A(n_10033),
.B(n_7003),
.Y(n_10678)
);

AND2x2_ASAP7_75t_L g10679 ( 
.A(n_10132),
.B(n_7005),
.Y(n_10679)
);

BUFx3_ASAP7_75t_L g10680 ( 
.A(n_10252),
.Y(n_10680)
);

NAND2x1p5_ASAP7_75t_L g10681 ( 
.A(n_10053),
.B(n_10057),
.Y(n_10681)
);

BUFx6f_ASAP7_75t_L g10682 ( 
.A(n_10133),
.Y(n_10682)
);

INVx1_ASAP7_75t_L g10683 ( 
.A(n_9954),
.Y(n_10683)
);

INVx1_ASAP7_75t_L g10684 ( 
.A(n_9956),
.Y(n_10684)
);

AND2x6_ASAP7_75t_L g10685 ( 
.A(n_10219),
.B(n_6586),
.Y(n_10685)
);

BUFx6f_ASAP7_75t_L g10686 ( 
.A(n_10141),
.Y(n_10686)
);

INVx3_ASAP7_75t_L g10687 ( 
.A(n_10143),
.Y(n_10687)
);

INVx3_ASAP7_75t_L g10688 ( 
.A(n_10105),
.Y(n_10688)
);

INVx4_ASAP7_75t_L g10689 ( 
.A(n_10218),
.Y(n_10689)
);

BUFx6f_ASAP7_75t_L g10690 ( 
.A(n_9909),
.Y(n_10690)
);

NOR2xp33_ASAP7_75t_L g10691 ( 
.A(n_10058),
.B(n_7006),
.Y(n_10691)
);

OR2x6_ASAP7_75t_L g10692 ( 
.A(n_10213),
.B(n_9989),
.Y(n_10692)
);

AND2x2_ASAP7_75t_L g10693 ( 
.A(n_10021),
.B(n_7009),
.Y(n_10693)
);

INVx3_ASAP7_75t_L g10694 ( 
.A(n_10106),
.Y(n_10694)
);

BUFx3_ASAP7_75t_L g10695 ( 
.A(n_10159),
.Y(n_10695)
);

AOI22xp33_ASAP7_75t_L g10696 ( 
.A1(n_9974),
.A2(n_7115),
.B1(n_7146),
.B2(n_7069),
.Y(n_10696)
);

NOR2x1p5_ASAP7_75t_L g10697 ( 
.A(n_10060),
.B(n_7010),
.Y(n_10697)
);

INVx2_ASAP7_75t_SL g10698 ( 
.A(n_9834),
.Y(n_10698)
);

AND2x6_ASAP7_75t_L g10699 ( 
.A(n_10215),
.B(n_6588),
.Y(n_10699)
);

NOR2x1p5_ASAP7_75t_L g10700 ( 
.A(n_10061),
.B(n_7014),
.Y(n_10700)
);

INVx2_ASAP7_75t_L g10701 ( 
.A(n_9957),
.Y(n_10701)
);

INVx1_ASAP7_75t_L g10702 ( 
.A(n_9960),
.Y(n_10702)
);

AND2x4_ASAP7_75t_L g10703 ( 
.A(n_10131),
.B(n_6589),
.Y(n_10703)
);

BUFx2_ASAP7_75t_L g10704 ( 
.A(n_9909),
.Y(n_10704)
);

OR2x6_ASAP7_75t_L g10705 ( 
.A(n_10065),
.B(n_6611),
.Y(n_10705)
);

NAND2xp5_ASAP7_75t_SL g10706 ( 
.A(n_10074),
.B(n_7024),
.Y(n_10706)
);

BUFx3_ASAP7_75t_L g10707 ( 
.A(n_10161),
.Y(n_10707)
);

AOI22xp33_ASAP7_75t_L g10708 ( 
.A1(n_9975),
.A2(n_9977),
.B1(n_10007),
.B2(n_9909),
.Y(n_10708)
);

NAND2x1p5_ASAP7_75t_L g10709 ( 
.A(n_10059),
.B(n_6612),
.Y(n_10709)
);

NAND2xp5_ASAP7_75t_L g10710 ( 
.A(n_9968),
.B(n_7026),
.Y(n_10710)
);

INVx2_ASAP7_75t_L g10711 ( 
.A(n_9945),
.Y(n_10711)
);

INVx2_ASAP7_75t_L g10712 ( 
.A(n_9963),
.Y(n_10712)
);

INVx3_ASAP7_75t_L g10713 ( 
.A(n_10071),
.Y(n_10713)
);

INVx3_ASAP7_75t_L g10714 ( 
.A(n_10072),
.Y(n_10714)
);

INVx2_ASAP7_75t_L g10715 ( 
.A(n_9966),
.Y(n_10715)
);

INVx5_ASAP7_75t_L g10716 ( 
.A(n_10218),
.Y(n_10716)
);

NAND2xp5_ASAP7_75t_L g10717 ( 
.A(n_9969),
.B(n_7031),
.Y(n_10717)
);

NAND2xp5_ASAP7_75t_L g10718 ( 
.A(n_9970),
.B(n_7033),
.Y(n_10718)
);

INVx4_ASAP7_75t_L g10719 ( 
.A(n_10218),
.Y(n_10719)
);

NAND2xp5_ASAP7_75t_L g10720 ( 
.A(n_9973),
.B(n_7037),
.Y(n_10720)
);

AND2x2_ASAP7_75t_L g10721 ( 
.A(n_10245),
.B(n_7039),
.Y(n_10721)
);

INVx2_ASAP7_75t_L g10722 ( 
.A(n_9978),
.Y(n_10722)
);

NAND2xp5_ASAP7_75t_L g10723 ( 
.A(n_9982),
.B(n_7040),
.Y(n_10723)
);

INVx1_ASAP7_75t_L g10724 ( 
.A(n_10113),
.Y(n_10724)
);

BUFx4f_ASAP7_75t_L g10725 ( 
.A(n_10007),
.Y(n_10725)
);

OAI21xp33_ASAP7_75t_L g10726 ( 
.A1(n_10190),
.A2(n_7050),
.B(n_7047),
.Y(n_10726)
);

NOR2xp33_ASAP7_75t_L g10727 ( 
.A(n_10185),
.B(n_7052),
.Y(n_10727)
);

INVx4_ASAP7_75t_L g10728 ( 
.A(n_10007),
.Y(n_10728)
);

AND2x4_ASAP7_75t_L g10729 ( 
.A(n_10138),
.B(n_6617),
.Y(n_10729)
);

INVx2_ASAP7_75t_L g10730 ( 
.A(n_9983),
.Y(n_10730)
);

NAND2xp5_ASAP7_75t_SL g10731 ( 
.A(n_10089),
.B(n_7055),
.Y(n_10731)
);

INVx2_ASAP7_75t_L g10732 ( 
.A(n_9984),
.Y(n_10732)
);

INVx2_ASAP7_75t_SL g10733 ( 
.A(n_10075),
.Y(n_10733)
);

AND2x4_ASAP7_75t_L g10734 ( 
.A(n_10142),
.B(n_6621),
.Y(n_10734)
);

INVx1_ASAP7_75t_L g10735 ( 
.A(n_10121),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_10125),
.Y(n_10736)
);

INVx2_ASAP7_75t_L g10737 ( 
.A(n_9985),
.Y(n_10737)
);

AND2x4_ASAP7_75t_L g10738 ( 
.A(n_10144),
.B(n_10148),
.Y(n_10738)
);

AND2x2_ASAP7_75t_L g10739 ( 
.A(n_9862),
.B(n_7057),
.Y(n_10739)
);

AND2x4_ASAP7_75t_L g10740 ( 
.A(n_10150),
.B(n_6623),
.Y(n_10740)
);

NAND2xp5_ASAP7_75t_L g10741 ( 
.A(n_10003),
.B(n_7058),
.Y(n_10741)
);

INVx1_ASAP7_75t_L g10742 ( 
.A(n_10127),
.Y(n_10742)
);

INVx4_ASAP7_75t_L g10743 ( 
.A(n_10076),
.Y(n_10743)
);

AND2x6_ASAP7_75t_L g10744 ( 
.A(n_10216),
.B(n_6624),
.Y(n_10744)
);

INVx1_ASAP7_75t_L g10745 ( 
.A(n_10004),
.Y(n_10745)
);

INVx1_ASAP7_75t_L g10746 ( 
.A(n_10087),
.Y(n_10746)
);

INVx4_ASAP7_75t_L g10747 ( 
.A(n_10095),
.Y(n_10747)
);

INVx2_ASAP7_75t_L g10748 ( 
.A(n_10187),
.Y(n_10748)
);

HB1xp67_ASAP7_75t_L g10749 ( 
.A(n_10069),
.Y(n_10749)
);

CKINVDCx5p33_ASAP7_75t_R g10750 ( 
.A(n_10247),
.Y(n_10750)
);

AOI22xp33_ASAP7_75t_L g10751 ( 
.A1(n_10208),
.A2(n_7242),
.B1(n_7302),
.B2(n_7154),
.Y(n_10751)
);

INVx2_ASAP7_75t_L g10752 ( 
.A(n_10189),
.Y(n_10752)
);

AND2x6_ASAP7_75t_L g10753 ( 
.A(n_10170),
.B(n_10078),
.Y(n_10753)
);

NAND2xp5_ASAP7_75t_L g10754 ( 
.A(n_10183),
.B(n_7059),
.Y(n_10754)
);

INVx1_ASAP7_75t_L g10755 ( 
.A(n_10099),
.Y(n_10755)
);

NAND2xp5_ASAP7_75t_L g10756 ( 
.A(n_10157),
.B(n_7060),
.Y(n_10756)
);

INVx2_ASAP7_75t_SL g10757 ( 
.A(n_10164),
.Y(n_10757)
);

NAND2xp33_ASAP7_75t_L g10758 ( 
.A(n_10191),
.B(n_7065),
.Y(n_10758)
);

NAND2xp5_ASAP7_75t_SL g10759 ( 
.A(n_10220),
.B(n_7066),
.Y(n_10759)
);

INVx3_ASAP7_75t_L g10760 ( 
.A(n_10079),
.Y(n_10760)
);

NAND2xp5_ASAP7_75t_L g10761 ( 
.A(n_10134),
.B(n_7067),
.Y(n_10761)
);

AND2x6_ASAP7_75t_L g10762 ( 
.A(n_10081),
.B(n_6628),
.Y(n_10762)
);

AND2x2_ASAP7_75t_L g10763 ( 
.A(n_9803),
.B(n_7071),
.Y(n_10763)
);

NAND2xp5_ASAP7_75t_SL g10764 ( 
.A(n_10640),
.B(n_10096),
.Y(n_10764)
);

OAI22xp5_ASAP7_75t_L g10765 ( 
.A1(n_10499),
.A2(n_10202),
.B1(n_10153),
.B2(n_10082),
.Y(n_10765)
);

NAND2xp5_ASAP7_75t_L g10766 ( 
.A(n_10467),
.B(n_9836),
.Y(n_10766)
);

INVx1_ASAP7_75t_L g10767 ( 
.A(n_10255),
.Y(n_10767)
);

NOR2xp67_ASAP7_75t_L g10768 ( 
.A(n_10254),
.B(n_10100),
.Y(n_10768)
);

OR2x2_ASAP7_75t_L g10769 ( 
.A(n_10445),
.B(n_9771),
.Y(n_10769)
);

NAND2xp33_ASAP7_75t_SL g10770 ( 
.A(n_10407),
.B(n_10399),
.Y(n_10770)
);

BUFx6f_ASAP7_75t_L g10771 ( 
.A(n_10375),
.Y(n_10771)
);

BUFx8_ASAP7_75t_L g10772 ( 
.A(n_10257),
.Y(n_10772)
);

NAND2xp5_ASAP7_75t_SL g10773 ( 
.A(n_10646),
.B(n_10167),
.Y(n_10773)
);

AOI22xp33_ASAP7_75t_L g10774 ( 
.A1(n_10426),
.A2(n_9747),
.B1(n_9725),
.B2(n_10173),
.Y(n_10774)
);

NAND2xp5_ASAP7_75t_L g10775 ( 
.A(n_10492),
.B(n_9972),
.Y(n_10775)
);

OR2x2_ASAP7_75t_L g10776 ( 
.A(n_10324),
.B(n_10424),
.Y(n_10776)
);

INVx1_ASAP7_75t_L g10777 ( 
.A(n_10258),
.Y(n_10777)
);

NAND2xp33_ASAP7_75t_L g10778 ( 
.A(n_10750),
.B(n_10175),
.Y(n_10778)
);

AOI22xp5_ASAP7_75t_L g10779 ( 
.A1(n_10360),
.A2(n_10126),
.B1(n_9925),
.B2(n_9980),
.Y(n_10779)
);

INVx1_ASAP7_75t_L g10780 ( 
.A(n_10272),
.Y(n_10780)
);

NAND2xp5_ASAP7_75t_L g10781 ( 
.A(n_10494),
.B(n_9976),
.Y(n_10781)
);

NAND2xp5_ASAP7_75t_L g10782 ( 
.A(n_10444),
.B(n_10036),
.Y(n_10782)
);

NAND2xp5_ASAP7_75t_L g10783 ( 
.A(n_10265),
.B(n_9828),
.Y(n_10783)
);

NAND2xp5_ASAP7_75t_SL g10784 ( 
.A(n_10517),
.B(n_10253),
.Y(n_10784)
);

AND2x2_ASAP7_75t_L g10785 ( 
.A(n_10548),
.B(n_9857),
.Y(n_10785)
);

NAND2xp5_ASAP7_75t_L g10786 ( 
.A(n_10287),
.B(n_9962),
.Y(n_10786)
);

NOR2xp33_ASAP7_75t_L g10787 ( 
.A(n_10398),
.B(n_10262),
.Y(n_10787)
);

INVx1_ASAP7_75t_L g10788 ( 
.A(n_10273),
.Y(n_10788)
);

INVx2_ASAP7_75t_L g10789 ( 
.A(n_10275),
.Y(n_10789)
);

INVxp67_ASAP7_75t_L g10790 ( 
.A(n_10521),
.Y(n_10790)
);

INVx2_ASAP7_75t_L g10791 ( 
.A(n_10281),
.Y(n_10791)
);

NAND2x1p5_ASAP7_75t_L g10792 ( 
.A(n_10389),
.B(n_10086),
.Y(n_10792)
);

INVxp67_ASAP7_75t_R g10793 ( 
.A(n_10269),
.Y(n_10793)
);

NAND2xp5_ASAP7_75t_SL g10794 ( 
.A(n_10579),
.B(n_10615),
.Y(n_10794)
);

INVx2_ASAP7_75t_L g10795 ( 
.A(n_10284),
.Y(n_10795)
);

NAND2xp5_ASAP7_75t_L g10796 ( 
.A(n_10287),
.B(n_10184),
.Y(n_10796)
);

NOR2xp33_ASAP7_75t_L g10797 ( 
.A(n_10302),
.B(n_10217),
.Y(n_10797)
);

NAND2xp5_ASAP7_75t_SL g10798 ( 
.A(n_10615),
.B(n_9881),
.Y(n_10798)
);

NAND2xp5_ASAP7_75t_L g10799 ( 
.A(n_10317),
.B(n_10186),
.Y(n_10799)
);

NAND2xp5_ASAP7_75t_L g10800 ( 
.A(n_10304),
.B(n_10188),
.Y(n_10800)
);

NOR3xp33_ASAP7_75t_L g10801 ( 
.A(n_10666),
.B(n_10678),
.C(n_10507),
.Y(n_10801)
);

INVx1_ASAP7_75t_L g10802 ( 
.A(n_10286),
.Y(n_10802)
);

INVxp67_ASAP7_75t_L g10803 ( 
.A(n_10553),
.Y(n_10803)
);

INVx2_ASAP7_75t_SL g10804 ( 
.A(n_10433),
.Y(n_10804)
);

INVx2_ASAP7_75t_L g10805 ( 
.A(n_10307),
.Y(n_10805)
);

AOI22xp5_ASAP7_75t_L g10806 ( 
.A1(n_10364),
.A2(n_10097),
.B1(n_10039),
.B2(n_10064),
.Y(n_10806)
);

NAND2xp5_ASAP7_75t_L g10807 ( 
.A(n_10280),
.B(n_10068),
.Y(n_10807)
);

AND2x4_ASAP7_75t_SL g10808 ( 
.A(n_10259),
.B(n_10285),
.Y(n_10808)
);

INVx2_ASAP7_75t_L g10809 ( 
.A(n_10310),
.Y(n_10809)
);

NAND2xp5_ASAP7_75t_L g10810 ( 
.A(n_10495),
.B(n_10090),
.Y(n_10810)
);

OAI22xp5_ASAP7_75t_L g10811 ( 
.A1(n_10361),
.A2(n_10094),
.B1(n_10102),
.B2(n_10214),
.Y(n_10811)
);

AND2x2_ASAP7_75t_L g10812 ( 
.A(n_10374),
.B(n_10558),
.Y(n_10812)
);

NOR2xp33_ASAP7_75t_L g10813 ( 
.A(n_10458),
.B(n_10093),
.Y(n_10813)
);

NAND2xp5_ASAP7_75t_SL g10814 ( 
.A(n_10716),
.B(n_10234),
.Y(n_10814)
);

INVx1_ASAP7_75t_L g10815 ( 
.A(n_10313),
.Y(n_10815)
);

NAND2xp5_ASAP7_75t_L g10816 ( 
.A(n_10271),
.B(n_10026),
.Y(n_10816)
);

INVx1_ASAP7_75t_SL g10817 ( 
.A(n_10466),
.Y(n_10817)
);

NAND2xp5_ASAP7_75t_L g10818 ( 
.A(n_10369),
.B(n_10101),
.Y(n_10818)
);

INVxp67_ASAP7_75t_L g10819 ( 
.A(n_10279),
.Y(n_10819)
);

NAND2xp5_ASAP7_75t_L g10820 ( 
.A(n_10378),
.B(n_10104),
.Y(n_10820)
);

AND2x2_ASAP7_75t_L g10821 ( 
.A(n_10446),
.B(n_10009),
.Y(n_10821)
);

AND2x2_ASAP7_75t_L g10822 ( 
.A(n_10464),
.B(n_10155),
.Y(n_10822)
);

NOR2xp33_ASAP7_75t_L g10823 ( 
.A(n_10266),
.B(n_9799),
.Y(n_10823)
);

AND2x2_ASAP7_75t_L g10824 ( 
.A(n_10509),
.B(n_9981),
.Y(n_10824)
);

INVx1_ASAP7_75t_L g10825 ( 
.A(n_10315),
.Y(n_10825)
);

NOR2xp67_ASAP7_75t_L g10826 ( 
.A(n_10288),
.B(n_10109),
.Y(n_10826)
);

INVx1_ASAP7_75t_L g10827 ( 
.A(n_10323),
.Y(n_10827)
);

CKINVDCx20_ASAP7_75t_R g10828 ( 
.A(n_10263),
.Y(n_10828)
);

NAND2xp5_ASAP7_75t_L g10829 ( 
.A(n_10754),
.B(n_10098),
.Y(n_10829)
);

AOI22xp33_ASAP7_75t_L g10830 ( 
.A1(n_10693),
.A2(n_9805),
.B1(n_10116),
.B2(n_9899),
.Y(n_10830)
);

NAND2xp5_ASAP7_75t_SL g10831 ( 
.A(n_10716),
.B(n_10088),
.Y(n_10831)
);

NAND2xp5_ASAP7_75t_SL g10832 ( 
.A(n_10278),
.B(n_10122),
.Y(n_10832)
);

INVx2_ASAP7_75t_L g10833 ( 
.A(n_10329),
.Y(n_10833)
);

NAND2xp5_ASAP7_75t_SL g10834 ( 
.A(n_10550),
.B(n_10128),
.Y(n_10834)
);

NAND2xp5_ASAP7_75t_L g10835 ( 
.A(n_10283),
.B(n_10043),
.Y(n_10835)
);

INVx2_ASAP7_75t_SL g10836 ( 
.A(n_10433),
.Y(n_10836)
);

NOR2xp33_ASAP7_75t_L g10837 ( 
.A(n_10581),
.B(n_10152),
.Y(n_10837)
);

INVx2_ASAP7_75t_L g10838 ( 
.A(n_10333),
.Y(n_10838)
);

NAND2xp5_ASAP7_75t_L g10839 ( 
.A(n_10504),
.B(n_10195),
.Y(n_10839)
);

NAND2xp5_ASAP7_75t_L g10840 ( 
.A(n_10519),
.B(n_10197),
.Y(n_10840)
);

O2A1O1Ixp33_ASAP7_75t_L g10841 ( 
.A1(n_10554),
.A2(n_6647),
.B(n_6651),
.C(n_6640),
.Y(n_10841)
);

NAND2xp5_ASAP7_75t_L g10842 ( 
.A(n_10534),
.B(n_10210),
.Y(n_10842)
);

NAND2xp5_ASAP7_75t_L g10843 ( 
.A(n_10545),
.B(n_10198),
.Y(n_10843)
);

INVx2_ASAP7_75t_L g10844 ( 
.A(n_10335),
.Y(n_10844)
);

INVx1_ASAP7_75t_L g10845 ( 
.A(n_10344),
.Y(n_10845)
);

NAND2xp5_ASAP7_75t_L g10846 ( 
.A(n_10577),
.B(n_6654),
.Y(n_10846)
);

AND2x4_ASAP7_75t_SL g10847 ( 
.A(n_10268),
.B(n_6657),
.Y(n_10847)
);

NAND2xp5_ASAP7_75t_SL g10848 ( 
.A(n_10520),
.B(n_7074),
.Y(n_10848)
);

BUFx6f_ASAP7_75t_L g10849 ( 
.A(n_10292),
.Y(n_10849)
);

OR2x2_ASAP7_75t_L g10850 ( 
.A(n_10400),
.B(n_10028),
.Y(n_10850)
);

NAND2xp5_ASAP7_75t_L g10851 ( 
.A(n_10584),
.B(n_6663),
.Y(n_10851)
);

NAND2xp5_ASAP7_75t_SL g10852 ( 
.A(n_10597),
.B(n_7077),
.Y(n_10852)
);

INVx2_ASAP7_75t_L g10853 ( 
.A(n_10347),
.Y(n_10853)
);

NAND2xp5_ASAP7_75t_SL g10854 ( 
.A(n_10572),
.B(n_7078),
.Y(n_10854)
);

OAI22xp5_ASAP7_75t_L g10855 ( 
.A1(n_10760),
.A2(n_10168),
.B1(n_7090),
.B2(n_7091),
.Y(n_10855)
);

BUFx3_ASAP7_75t_L g10856 ( 
.A(n_10389),
.Y(n_10856)
);

NAND2xp5_ASAP7_75t_SL g10857 ( 
.A(n_10298),
.B(n_7084),
.Y(n_10857)
);

NAND2xp5_ASAP7_75t_SL g10858 ( 
.A(n_10497),
.B(n_7092),
.Y(n_10858)
);

INVx1_ASAP7_75t_L g10859 ( 
.A(n_10350),
.Y(n_10859)
);

NAND2xp5_ASAP7_75t_L g10860 ( 
.A(n_10355),
.B(n_6679),
.Y(n_10860)
);

NAND2xp5_ASAP7_75t_L g10861 ( 
.A(n_10356),
.B(n_6681),
.Y(n_10861)
);

OAI221xp5_ASAP7_75t_L g10862 ( 
.A1(n_10573),
.A2(n_6700),
.B1(n_6701),
.B2(n_6689),
.C(n_6682),
.Y(n_10862)
);

AOI22xp33_ASAP7_75t_L g10863 ( 
.A1(n_10658),
.A2(n_6709),
.B1(n_6717),
.B2(n_6705),
.Y(n_10863)
);

A2O1A1Ixp33_ASAP7_75t_L g10864 ( 
.A1(n_10649),
.A2(n_9732),
.B(n_6720),
.C(n_6724),
.Y(n_10864)
);

INVx1_ASAP7_75t_L g10865 ( 
.A(n_10359),
.Y(n_10865)
);

INVx1_ASAP7_75t_L g10866 ( 
.A(n_10363),
.Y(n_10866)
);

INVx2_ASAP7_75t_L g10867 ( 
.A(n_10365),
.Y(n_10867)
);

NAND2xp5_ASAP7_75t_L g10868 ( 
.A(n_10368),
.B(n_6719),
.Y(n_10868)
);

AOI22xp33_ASAP7_75t_L g10869 ( 
.A1(n_10671),
.A2(n_6728),
.B1(n_6732),
.B2(n_6725),
.Y(n_10869)
);

AND2x4_ASAP7_75t_L g10870 ( 
.A(n_10260),
.B(n_6736),
.Y(n_10870)
);

NOR2xp33_ASAP7_75t_L g10871 ( 
.A(n_10477),
.B(n_7094),
.Y(n_10871)
);

NAND2xp5_ASAP7_75t_SL g10872 ( 
.A(n_10358),
.B(n_7096),
.Y(n_10872)
);

INVx1_ASAP7_75t_L g10873 ( 
.A(n_10372),
.Y(n_10873)
);

NAND2xp5_ASAP7_75t_L g10874 ( 
.A(n_10377),
.B(n_6744),
.Y(n_10874)
);

NAND2xp5_ASAP7_75t_SL g10875 ( 
.A(n_10680),
.B(n_7099),
.Y(n_10875)
);

NAND2xp5_ASAP7_75t_L g10876 ( 
.A(n_10667),
.B(n_6748),
.Y(n_10876)
);

NAND2xp5_ASAP7_75t_L g10877 ( 
.A(n_10411),
.B(n_6755),
.Y(n_10877)
);

NAND2xp5_ASAP7_75t_L g10878 ( 
.A(n_10756),
.B(n_10761),
.Y(n_10878)
);

NAND2xp5_ASAP7_75t_L g10879 ( 
.A(n_10618),
.B(n_6776),
.Y(n_10879)
);

NAND2xp5_ASAP7_75t_SL g10880 ( 
.A(n_10513),
.B(n_7102),
.Y(n_10880)
);

NAND2xp5_ASAP7_75t_L g10881 ( 
.A(n_10624),
.B(n_6784),
.Y(n_10881)
);

AND2x2_ASAP7_75t_L g10882 ( 
.A(n_10524),
.B(n_10533),
.Y(n_10882)
);

NAND2xp5_ASAP7_75t_SL g10883 ( 
.A(n_10518),
.B(n_7103),
.Y(n_10883)
);

NAND2xp33_ASAP7_75t_L g10884 ( 
.A(n_10753),
.B(n_7107),
.Y(n_10884)
);

AND2x2_ASAP7_75t_L g10885 ( 
.A(n_10471),
.B(n_7119),
.Y(n_10885)
);

NAND2xp5_ASAP7_75t_L g10886 ( 
.A(n_10634),
.B(n_6789),
.Y(n_10886)
);

NAND2xp5_ASAP7_75t_L g10887 ( 
.A(n_10638),
.B(n_6792),
.Y(n_10887)
);

INVx2_ASAP7_75t_L g10888 ( 
.A(n_10745),
.Y(n_10888)
);

AND2x2_ASAP7_75t_L g10889 ( 
.A(n_10488),
.B(n_10566),
.Y(n_10889)
);

NOR2xp67_ASAP7_75t_L g10890 ( 
.A(n_10455),
.B(n_10478),
.Y(n_10890)
);

NAND2xp5_ASAP7_75t_SL g10891 ( 
.A(n_10306),
.B(n_7121),
.Y(n_10891)
);

NAND2xp5_ASAP7_75t_L g10892 ( 
.A(n_10645),
.B(n_6793),
.Y(n_10892)
);

INVx1_ASAP7_75t_SL g10893 ( 
.A(n_10332),
.Y(n_10893)
);

INVx1_ASAP7_75t_L g10894 ( 
.A(n_10448),
.Y(n_10894)
);

INVx1_ASAP7_75t_L g10895 ( 
.A(n_10451),
.Y(n_10895)
);

INVx1_ASAP7_75t_L g10896 ( 
.A(n_10453),
.Y(n_10896)
);

BUFx5_ASAP7_75t_L g10897 ( 
.A(n_10753),
.Y(n_10897)
);

NAND2xp5_ASAP7_75t_L g10898 ( 
.A(n_10653),
.B(n_6797),
.Y(n_10898)
);

INVx1_ASAP7_75t_L g10899 ( 
.A(n_10461),
.Y(n_10899)
);

INVx2_ASAP7_75t_L g10900 ( 
.A(n_10722),
.Y(n_10900)
);

AOI221xp5_ASAP7_75t_L g10901 ( 
.A1(n_10663),
.A2(n_6826),
.B1(n_6830),
.B2(n_6819),
.C(n_6813),
.Y(n_10901)
);

INVx2_ASAP7_75t_L g10902 ( 
.A(n_10730),
.Y(n_10902)
);

INVxp67_ASAP7_75t_L g10903 ( 
.A(n_10582),
.Y(n_10903)
);

OAI22xp5_ASAP7_75t_L g10904 ( 
.A1(n_10463),
.A2(n_7124),
.B1(n_7128),
.B2(n_7123),
.Y(n_10904)
);

NAND2xp5_ASAP7_75t_L g10905 ( 
.A(n_10724),
.B(n_6834),
.Y(n_10905)
);

NAND2xp5_ASAP7_75t_SL g10906 ( 
.A(n_10437),
.B(n_7131),
.Y(n_10906)
);

NAND2xp5_ASAP7_75t_SL g10907 ( 
.A(n_10437),
.B(n_7132),
.Y(n_10907)
);

NOR2xp33_ASAP7_75t_L g10908 ( 
.A(n_10294),
.B(n_7134),
.Y(n_10908)
);

NOR2xp33_ASAP7_75t_L g10909 ( 
.A(n_10546),
.B(n_7137),
.Y(n_10909)
);

HB1xp67_ASAP7_75t_L g10910 ( 
.A(n_10516),
.Y(n_10910)
);

AOI22xp33_ASAP7_75t_L g10911 ( 
.A1(n_10679),
.A2(n_6837),
.B1(n_6850),
.B2(n_6835),
.Y(n_10911)
);

NAND3xp33_ASAP7_75t_L g10912 ( 
.A(n_10661),
.B(n_7142),
.C(n_7139),
.Y(n_10912)
);

INVx2_ASAP7_75t_L g10913 ( 
.A(n_10732),
.Y(n_10913)
);

NAND2xp5_ASAP7_75t_SL g10914 ( 
.A(n_10516),
.B(n_7152),
.Y(n_10914)
);

AND2x2_ASAP7_75t_SL g10915 ( 
.A(n_10725),
.B(n_6863),
.Y(n_10915)
);

INVx2_ASAP7_75t_L g10916 ( 
.A(n_10737),
.Y(n_10916)
);

NAND2xp5_ASAP7_75t_SL g10917 ( 
.A(n_10528),
.B(n_7155),
.Y(n_10917)
);

O2A1O1Ixp5_ASAP7_75t_L g10918 ( 
.A1(n_10706),
.A2(n_6881),
.B(n_6883),
.C(n_6865),
.Y(n_10918)
);

INVx1_ASAP7_75t_L g10919 ( 
.A(n_10469),
.Y(n_10919)
);

INVx2_ASAP7_75t_L g10920 ( 
.A(n_10480),
.Y(n_10920)
);

NAND2xp5_ASAP7_75t_L g10921 ( 
.A(n_10735),
.B(n_6888),
.Y(n_10921)
);

INVx1_ASAP7_75t_SL g10922 ( 
.A(n_10530),
.Y(n_10922)
);

INVx1_ASAP7_75t_L g10923 ( 
.A(n_10482),
.Y(n_10923)
);

NAND2xp5_ASAP7_75t_SL g10924 ( 
.A(n_10528),
.B(n_7157),
.Y(n_10924)
);

INVx1_ASAP7_75t_L g10925 ( 
.A(n_10484),
.Y(n_10925)
);

NAND2xp5_ASAP7_75t_L g10926 ( 
.A(n_10736),
.B(n_10742),
.Y(n_10926)
);

NAND2xp5_ASAP7_75t_SL g10927 ( 
.A(n_10371),
.B(n_7165),
.Y(n_10927)
);

NAND2xp5_ASAP7_75t_L g10928 ( 
.A(n_10379),
.B(n_6889),
.Y(n_10928)
);

NAND2xp5_ASAP7_75t_L g10929 ( 
.A(n_10405),
.B(n_6890),
.Y(n_10929)
);

NAND2xp5_ASAP7_75t_L g10930 ( 
.A(n_10409),
.B(n_6892),
.Y(n_10930)
);

NOR2xp33_ASAP7_75t_L g10931 ( 
.A(n_10270),
.B(n_10392),
.Y(n_10931)
);

NAND2xp5_ASAP7_75t_L g10932 ( 
.A(n_10410),
.B(n_6895),
.Y(n_10932)
);

INVx2_ASAP7_75t_SL g10933 ( 
.A(n_10267),
.Y(n_10933)
);

NAND2xp5_ASAP7_75t_L g10934 ( 
.A(n_10414),
.B(n_6901),
.Y(n_10934)
);

NOR2xp33_ASAP7_75t_SL g10935 ( 
.A(n_10338),
.B(n_7166),
.Y(n_10935)
);

INVx2_ASAP7_75t_L g10936 ( 
.A(n_10485),
.Y(n_10936)
);

INVx2_ASAP7_75t_SL g10937 ( 
.A(n_10292),
.Y(n_10937)
);

INVx2_ASAP7_75t_L g10938 ( 
.A(n_10493),
.Y(n_10938)
);

NOR2xp67_ASAP7_75t_L g10939 ( 
.A(n_10428),
.B(n_4554),
.Y(n_10939)
);

INVx2_ASAP7_75t_L g10940 ( 
.A(n_10500),
.Y(n_10940)
);

INVx2_ASAP7_75t_L g10941 ( 
.A(n_10502),
.Y(n_10941)
);

NAND2xp5_ASAP7_75t_SL g10942 ( 
.A(n_10538),
.B(n_7168),
.Y(n_10942)
);

NOR2xp33_ASAP7_75t_L g10943 ( 
.A(n_10420),
.B(n_7173),
.Y(n_10943)
);

INVx2_ASAP7_75t_L g10944 ( 
.A(n_10510),
.Y(n_10944)
);

NAND2xp5_ASAP7_75t_L g10945 ( 
.A(n_10421),
.B(n_6908),
.Y(n_10945)
);

INVx1_ASAP7_75t_L g10946 ( 
.A(n_10511),
.Y(n_10946)
);

INVx2_ASAP7_75t_L g10947 ( 
.A(n_10523),
.Y(n_10947)
);

NAND2xp5_ASAP7_75t_SL g10948 ( 
.A(n_10636),
.B(n_7176),
.Y(n_10948)
);

INVx1_ASAP7_75t_L g10949 ( 
.A(n_10526),
.Y(n_10949)
);

INVx3_ASAP7_75t_L g10950 ( 
.A(n_10542),
.Y(n_10950)
);

OAI22xp5_ASAP7_75t_L g10951 ( 
.A1(n_10541),
.A2(n_7178),
.B1(n_7179),
.B2(n_7177),
.Y(n_10951)
);

NAND2xp5_ASAP7_75t_SL g10952 ( 
.A(n_10636),
.B(n_7180),
.Y(n_10952)
);

NAND2xp33_ASAP7_75t_L g10953 ( 
.A(n_10708),
.B(n_7182),
.Y(n_10953)
);

INVx2_ASAP7_75t_L g10954 ( 
.A(n_10557),
.Y(n_10954)
);

INVx1_ASAP7_75t_L g10955 ( 
.A(n_10562),
.Y(n_10955)
);

INVx1_ASAP7_75t_L g10956 ( 
.A(n_10564),
.Y(n_10956)
);

INVx1_ASAP7_75t_L g10957 ( 
.A(n_10567),
.Y(n_10957)
);

INVxp67_ASAP7_75t_L g10958 ( 
.A(n_10449),
.Y(n_10958)
);

AOI22xp33_ASAP7_75t_L g10959 ( 
.A1(n_10763),
.A2(n_6913),
.B1(n_6929),
.B2(n_6911),
.Y(n_10959)
);

INVx6_ASAP7_75t_L g10960 ( 
.A(n_10543),
.Y(n_10960)
);

INVxp67_ASAP7_75t_L g10961 ( 
.A(n_10481),
.Y(n_10961)
);

INVx2_ASAP7_75t_L g10962 ( 
.A(n_10576),
.Y(n_10962)
);

NAND2xp33_ASAP7_75t_SL g10963 ( 
.A(n_10689),
.B(n_7184),
.Y(n_10963)
);

NOR2xp33_ASAP7_75t_L g10964 ( 
.A(n_10300),
.B(n_7185),
.Y(n_10964)
);

INVx2_ASAP7_75t_L g10965 ( 
.A(n_10585),
.Y(n_10965)
);

INVx2_ASAP7_75t_SL g10966 ( 
.A(n_10293),
.Y(n_10966)
);

INVx2_ASAP7_75t_L g10967 ( 
.A(n_10587),
.Y(n_10967)
);

INVx2_ASAP7_75t_L g10968 ( 
.A(n_10592),
.Y(n_10968)
);

NOR2xp33_ASAP7_75t_L g10969 ( 
.A(n_10588),
.B(n_7186),
.Y(n_10969)
);

OAI21xp5_ASAP7_75t_L g10970 ( 
.A1(n_10452),
.A2(n_6933),
.B(n_6930),
.Y(n_10970)
);

INVx1_ASAP7_75t_L g10971 ( 
.A(n_10594),
.Y(n_10971)
);

NAND2xp5_ASAP7_75t_L g10972 ( 
.A(n_10601),
.B(n_6939),
.Y(n_10972)
);

INVx1_ASAP7_75t_L g10973 ( 
.A(n_10602),
.Y(n_10973)
);

NAND2xp5_ASAP7_75t_L g10974 ( 
.A(n_10604),
.B(n_6947),
.Y(n_10974)
);

BUFx5_ASAP7_75t_L g10975 ( 
.A(n_10609),
.Y(n_10975)
);

NAND2xp5_ASAP7_75t_SL g10976 ( 
.A(n_10345),
.B(n_7188),
.Y(n_10976)
);

INVx2_ASAP7_75t_L g10977 ( 
.A(n_10290),
.Y(n_10977)
);

NAND2xp5_ASAP7_75t_L g10978 ( 
.A(n_10321),
.B(n_6948),
.Y(n_10978)
);

INVx1_ASAP7_75t_L g10979 ( 
.A(n_10297),
.Y(n_10979)
);

NAND3xp33_ASAP7_75t_L g10980 ( 
.A(n_10529),
.B(n_7200),
.C(n_7190),
.Y(n_10980)
);

NAND2xp5_ASAP7_75t_L g10981 ( 
.A(n_10322),
.B(n_6954),
.Y(n_10981)
);

AND2x4_ASAP7_75t_L g10982 ( 
.A(n_10698),
.B(n_6960),
.Y(n_10982)
);

AND2x2_ASAP7_75t_L g10983 ( 
.A(n_10721),
.B(n_7201),
.Y(n_10983)
);

INVx1_ASAP7_75t_L g10984 ( 
.A(n_10309),
.Y(n_10984)
);

NOR2xp33_ASAP7_75t_L g10985 ( 
.A(n_10468),
.B(n_7202),
.Y(n_10985)
);

INVx1_ASAP7_75t_L g10986 ( 
.A(n_10436),
.Y(n_10986)
);

NAND2xp5_ASAP7_75t_L g10987 ( 
.A(n_10337),
.B(n_6968),
.Y(n_10987)
);

AOI22xp5_ASAP7_75t_L g10988 ( 
.A1(n_10367),
.A2(n_7206),
.B1(n_7212),
.B2(n_7204),
.Y(n_10988)
);

INVx1_ASAP7_75t_L g10989 ( 
.A(n_10441),
.Y(n_10989)
);

INVxp67_ASAP7_75t_L g10990 ( 
.A(n_10370),
.Y(n_10990)
);

NOR2xp33_ASAP7_75t_L g10991 ( 
.A(n_10490),
.B(n_7214),
.Y(n_10991)
);

AOI22xp5_ASAP7_75t_L g10992 ( 
.A1(n_10727),
.A2(n_7217),
.B1(n_7219),
.B2(n_7216),
.Y(n_10992)
);

INVx1_ASAP7_75t_L g10993 ( 
.A(n_10442),
.Y(n_10993)
);

NOR2xp33_ASAP7_75t_L g10994 ( 
.A(n_10388),
.B(n_7220),
.Y(n_10994)
);

AND2x2_ASAP7_75t_L g10995 ( 
.A(n_10575),
.B(n_7223),
.Y(n_10995)
);

NOR3xp33_ASAP7_75t_L g10996 ( 
.A(n_10261),
.B(n_6973),
.C(n_6972),
.Y(n_10996)
);

OAI22xp5_ASAP7_75t_SL g10997 ( 
.A1(n_10383),
.A2(n_7226),
.B1(n_7228),
.B2(n_7225),
.Y(n_10997)
);

NAND2xp5_ASAP7_75t_L g10998 ( 
.A(n_10341),
.B(n_6974),
.Y(n_10998)
);

INVx8_ASAP7_75t_L g10999 ( 
.A(n_10293),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_10443),
.Y(n_11000)
);

NAND2xp5_ASAP7_75t_SL g11001 ( 
.A(n_10719),
.B(n_7229),
.Y(n_11001)
);

INVx1_ASAP7_75t_L g11002 ( 
.A(n_10454),
.Y(n_11002)
);

NAND2xp33_ASAP7_75t_L g11003 ( 
.A(n_10690),
.B(n_7230),
.Y(n_11003)
);

INVx1_ASAP7_75t_L g11004 ( 
.A(n_10535),
.Y(n_11004)
);

NAND2xp5_ASAP7_75t_SL g11005 ( 
.A(n_10651),
.B(n_7232),
.Y(n_11005)
);

INVx2_ASAP7_75t_L g11006 ( 
.A(n_10256),
.Y(n_11006)
);

NOR2xp33_ASAP7_75t_SL g11007 ( 
.A(n_10264),
.B(n_7237),
.Y(n_11007)
);

AOI22xp5_ASAP7_75t_L g11008 ( 
.A1(n_10611),
.A2(n_7241),
.B1(n_7243),
.B2(n_7240),
.Y(n_11008)
);

NAND2xp5_ASAP7_75t_L g11009 ( 
.A(n_10348),
.B(n_6976),
.Y(n_11009)
);

NOR2xp33_ASAP7_75t_L g11010 ( 
.A(n_10626),
.B(n_7246),
.Y(n_11010)
);

AOI22xp33_ASAP7_75t_L g11011 ( 
.A1(n_10739),
.A2(n_6984),
.B1(n_6993),
.B2(n_6980),
.Y(n_11011)
);

INVx1_ASAP7_75t_L g11012 ( 
.A(n_10276),
.Y(n_11012)
);

INVx2_ASAP7_75t_L g11013 ( 
.A(n_10277),
.Y(n_11013)
);

NAND2xp5_ASAP7_75t_L g11014 ( 
.A(n_10349),
.B(n_7000),
.Y(n_11014)
);

NAND2xp5_ASAP7_75t_L g11015 ( 
.A(n_10352),
.B(n_7007),
.Y(n_11015)
);

OAI22xp33_ASAP7_75t_L g11016 ( 
.A1(n_10705),
.A2(n_7255),
.B1(n_7258),
.B2(n_7247),
.Y(n_11016)
);

NAND2xp5_ASAP7_75t_L g11017 ( 
.A(n_10366),
.B(n_7017),
.Y(n_11017)
);

O2A1O1Ixp33_ASAP7_75t_L g11018 ( 
.A1(n_10473),
.A2(n_7023),
.B(n_7030),
.C(n_7020),
.Y(n_11018)
);

INVx2_ASAP7_75t_SL g11019 ( 
.A(n_10299),
.Y(n_11019)
);

BUFx5_ASAP7_75t_L g11020 ( 
.A(n_10657),
.Y(n_11020)
);

OAI22xp33_ASAP7_75t_L g11021 ( 
.A1(n_10401),
.A2(n_7260),
.B1(n_7261),
.B2(n_7259),
.Y(n_11021)
);

NAND3xp33_ASAP7_75t_L g11022 ( 
.A(n_10629),
.B(n_7264),
.C(n_7262),
.Y(n_11022)
);

BUFx6f_ASAP7_75t_L g11023 ( 
.A(n_10299),
.Y(n_11023)
);

NAND2xp5_ASAP7_75t_L g11024 ( 
.A(n_10380),
.B(n_7035),
.Y(n_11024)
);

A2O1A1Ixp33_ASAP7_75t_L g11025 ( 
.A1(n_10635),
.A2(n_7061),
.B(n_7070),
.C(n_7056),
.Y(n_11025)
);

HB1xp67_ASAP7_75t_L g11026 ( 
.A(n_10274),
.Y(n_11026)
);

BUFx6f_ASAP7_75t_SL g11027 ( 
.A(n_10483),
.Y(n_11027)
);

OAI22xp5_ASAP7_75t_L g11028 ( 
.A1(n_10394),
.A2(n_7269),
.B1(n_7271),
.B2(n_7268),
.Y(n_11028)
);

NAND2xp5_ASAP7_75t_L g11029 ( 
.A(n_10403),
.B(n_7072),
.Y(n_11029)
);

INVxp33_ASAP7_75t_L g11030 ( 
.A(n_10417),
.Y(n_11030)
);

INVx3_ASAP7_75t_L g11031 ( 
.A(n_10291),
.Y(n_11031)
);

NOR2xp33_ASAP7_75t_L g11032 ( 
.A(n_10647),
.B(n_10691),
.Y(n_11032)
);

NAND2xp5_ASAP7_75t_L g11033 ( 
.A(n_10404),
.B(n_7081),
.Y(n_11033)
);

NAND2xp5_ASAP7_75t_L g11034 ( 
.A(n_10427),
.B(n_7082),
.Y(n_11034)
);

NOR2xp33_ASAP7_75t_L g11035 ( 
.A(n_10749),
.B(n_7272),
.Y(n_11035)
);

INVx1_ASAP7_75t_L g11036 ( 
.A(n_10660),
.Y(n_11036)
);

NAND2xp5_ASAP7_75t_SL g11037 ( 
.A(n_10651),
.B(n_10665),
.Y(n_11037)
);

AOI22xp33_ASAP7_75t_SL g11038 ( 
.A1(n_10662),
.A2(n_7275),
.B1(n_7278),
.B2(n_7274),
.Y(n_11038)
);

NAND2xp5_ASAP7_75t_L g11039 ( 
.A(n_10674),
.B(n_10701),
.Y(n_11039)
);

NAND2xp5_ASAP7_75t_L g11040 ( 
.A(n_10670),
.B(n_10683),
.Y(n_11040)
);

INVx1_ASAP7_75t_L g11041 ( 
.A(n_10684),
.Y(n_11041)
);

INVxp67_ASAP7_75t_SL g11042 ( 
.A(n_10357),
.Y(n_11042)
);

BUFx6f_ASAP7_75t_L g11043 ( 
.A(n_10314),
.Y(n_11043)
);

AND2x4_ASAP7_75t_SL g11044 ( 
.A(n_10296),
.B(n_10354),
.Y(n_11044)
);

INVx1_ASAP7_75t_L g11045 ( 
.A(n_10702),
.Y(n_11045)
);

INVx1_ASAP7_75t_L g11046 ( 
.A(n_10659),
.Y(n_11046)
);

NAND2xp5_ASAP7_75t_L g11047 ( 
.A(n_10316),
.B(n_7085),
.Y(n_11047)
);

AOI22xp33_ASAP7_75t_L g11048 ( 
.A1(n_10726),
.A2(n_7088),
.B1(n_7095),
.B2(n_7087),
.Y(n_11048)
);

NOR2xp67_ASAP7_75t_L g11049 ( 
.A(n_10688),
.B(n_10694),
.Y(n_11049)
);

INVx2_ASAP7_75t_L g11050 ( 
.A(n_10459),
.Y(n_11050)
);

BUFx6f_ASAP7_75t_L g11051 ( 
.A(n_10314),
.Y(n_11051)
);

NAND2xp5_ASAP7_75t_SL g11052 ( 
.A(n_10665),
.B(n_7279),
.Y(n_11052)
);

INVx1_ASAP7_75t_L g11053 ( 
.A(n_10755),
.Y(n_11053)
);

INVx2_ASAP7_75t_L g11054 ( 
.A(n_10460),
.Y(n_11054)
);

INVx2_ASAP7_75t_L g11055 ( 
.A(n_10474),
.Y(n_11055)
);

NOR2xp67_ASAP7_75t_L g11056 ( 
.A(n_10641),
.B(n_4555),
.Y(n_11056)
);

NAND2xp5_ASAP7_75t_L g11057 ( 
.A(n_10328),
.B(n_7101),
.Y(n_11057)
);

AO22x2_ASAP7_75t_L g11058 ( 
.A1(n_10552),
.A2(n_7113),
.B1(n_7114),
.B2(n_7105),
.Y(n_11058)
);

NAND2xp5_ASAP7_75t_L g11059 ( 
.A(n_10343),
.B(n_7116),
.Y(n_11059)
);

AOI22xp5_ASAP7_75t_L g11060 ( 
.A1(n_10644),
.A2(n_7282),
.B1(n_7283),
.B2(n_7281),
.Y(n_11060)
);

NAND2xp5_ASAP7_75t_L g11061 ( 
.A(n_10346),
.B(n_10353),
.Y(n_11061)
);

NAND2xp5_ASAP7_75t_L g11062 ( 
.A(n_10376),
.B(n_7118),
.Y(n_11062)
);

INVx2_ASAP7_75t_L g11063 ( 
.A(n_10496),
.Y(n_11063)
);

NOR3xp33_ASAP7_75t_L g11064 ( 
.A(n_10450),
.B(n_7129),
.C(n_7127),
.Y(n_11064)
);

NAND2xp5_ASAP7_75t_L g11065 ( 
.A(n_10387),
.B(n_7133),
.Y(n_11065)
);

INVx2_ASAP7_75t_L g11066 ( 
.A(n_10505),
.Y(n_11066)
);

INVx1_ASAP7_75t_L g11067 ( 
.A(n_10457),
.Y(n_11067)
);

INVx3_ASAP7_75t_L g11068 ( 
.A(n_10381),
.Y(n_11068)
);

NAND2xp5_ASAP7_75t_SL g11069 ( 
.A(n_10682),
.B(n_7285),
.Y(n_11069)
);

NOR2xp33_ASAP7_75t_L g11070 ( 
.A(n_10583),
.B(n_7291),
.Y(n_11070)
);

NAND2xp5_ASAP7_75t_L g11071 ( 
.A(n_10425),
.B(n_7138),
.Y(n_11071)
);

INVx2_ASAP7_75t_SL g11072 ( 
.A(n_10340),
.Y(n_11072)
);

NAND2xp5_ASAP7_75t_L g11073 ( 
.A(n_10623),
.B(n_7140),
.Y(n_11073)
);

AND2x2_ASAP7_75t_L g11074 ( 
.A(n_10590),
.B(n_7293),
.Y(n_11074)
);

NAND2xp5_ASAP7_75t_SL g11075 ( 
.A(n_10682),
.B(n_7296),
.Y(n_11075)
);

INVx8_ASAP7_75t_L g11076 ( 
.A(n_10340),
.Y(n_11076)
);

INVx2_ASAP7_75t_L g11077 ( 
.A(n_10506),
.Y(n_11077)
);

NAND2xp5_ASAP7_75t_L g11078 ( 
.A(n_10525),
.B(n_7141),
.Y(n_11078)
);

NAND2xp33_ASAP7_75t_L g11079 ( 
.A(n_10690),
.B(n_7297),
.Y(n_11079)
);

INVx1_ASAP7_75t_L g11080 ( 
.A(n_10532),
.Y(n_11080)
);

NAND2xp5_ASAP7_75t_SL g11081 ( 
.A(n_10336),
.B(n_7299),
.Y(n_11081)
);

BUFx3_ASAP7_75t_L g11082 ( 
.A(n_10305),
.Y(n_11082)
);

INVx1_ASAP7_75t_L g11083 ( 
.A(n_10547),
.Y(n_11083)
);

NAND2xp5_ASAP7_75t_L g11084 ( 
.A(n_10563),
.B(n_7145),
.Y(n_11084)
);

AND2x4_ASAP7_75t_L g11085 ( 
.A(n_10544),
.B(n_7147),
.Y(n_11085)
);

INVx2_ASAP7_75t_L g11086 ( 
.A(n_10580),
.Y(n_11086)
);

AOI221xp5_ASAP7_75t_L g11087 ( 
.A1(n_10475),
.A2(n_7159),
.B1(n_7163),
.B2(n_7156),
.C(n_7148),
.Y(n_11087)
);

BUFx3_ASAP7_75t_L g11088 ( 
.A(n_10308),
.Y(n_11088)
);

NAND2xp5_ASAP7_75t_SL g11089 ( 
.A(n_10686),
.B(n_7303),
.Y(n_11089)
);

NOR2xp33_ASAP7_75t_L g11090 ( 
.A(n_10501),
.B(n_7304),
.Y(n_11090)
);

OAI22xp33_ASAP7_75t_L g11091 ( 
.A1(n_10568),
.A2(n_7308),
.B1(n_7316),
.B2(n_7306),
.Y(n_11091)
);

AOI22xp33_ASAP7_75t_L g11092 ( 
.A1(n_10703),
.A2(n_7170),
.B1(n_7172),
.B2(n_7169),
.Y(n_11092)
);

NAND2xp5_ASAP7_75t_L g11093 ( 
.A(n_10586),
.B(n_7174),
.Y(n_11093)
);

NAND2xp5_ASAP7_75t_L g11094 ( 
.A(n_10589),
.B(n_7175),
.Y(n_11094)
);

INVx1_ASAP7_75t_L g11095 ( 
.A(n_10600),
.Y(n_11095)
);

INVx2_ASAP7_75t_L g11096 ( 
.A(n_10603),
.Y(n_11096)
);

NAND2xp5_ASAP7_75t_L g11097 ( 
.A(n_10606),
.B(n_7181),
.Y(n_11097)
);

INVx1_ASAP7_75t_L g11098 ( 
.A(n_10607),
.Y(n_11098)
);

NOR2xp33_ASAP7_75t_L g11099 ( 
.A(n_10643),
.B(n_7318),
.Y(n_11099)
);

INVx1_ASAP7_75t_SL g11100 ( 
.A(n_10318),
.Y(n_11100)
);

INVxp67_ASAP7_75t_SL g11101 ( 
.A(n_10386),
.Y(n_11101)
);

NAND2xp5_ASAP7_75t_L g11102 ( 
.A(n_10614),
.B(n_7187),
.Y(n_11102)
);

AND2x4_ASAP7_75t_SL g11103 ( 
.A(n_10416),
.B(n_7193),
.Y(n_11103)
);

NAND2xp5_ASAP7_75t_SL g11104 ( 
.A(n_10686),
.B(n_7323),
.Y(n_11104)
);

INVx2_ASAP7_75t_L g11105 ( 
.A(n_10617),
.Y(n_11105)
);

AOI22xp5_ASAP7_75t_L g11106 ( 
.A1(n_10331),
.A2(n_7338),
.B1(n_7339),
.B2(n_7334),
.Y(n_11106)
);

NOR3xp33_ASAP7_75t_L g11107 ( 
.A(n_10465),
.B(n_7196),
.C(n_7195),
.Y(n_11107)
);

AOI22xp33_ASAP7_75t_L g11108 ( 
.A1(n_10729),
.A2(n_7210),
.B1(n_7211),
.B2(n_7209),
.Y(n_11108)
);

INVx2_ASAP7_75t_L g11109 ( 
.A(n_10621),
.Y(n_11109)
);

NAND2xp33_ASAP7_75t_L g11110 ( 
.A(n_10699),
.B(n_7341),
.Y(n_11110)
);

NAND2xp5_ASAP7_75t_L g11111 ( 
.A(n_10627),
.B(n_7213),
.Y(n_11111)
);

INVx2_ASAP7_75t_L g11112 ( 
.A(n_10633),
.Y(n_11112)
);

NAND2xp5_ASAP7_75t_L g11113 ( 
.A(n_10639),
.B(n_7222),
.Y(n_11113)
);

INVx8_ASAP7_75t_L g11114 ( 
.A(n_10342),
.Y(n_11114)
);

INVx1_ASAP7_75t_L g11115 ( 
.A(n_10652),
.Y(n_11115)
);

NAND2xp5_ASAP7_75t_SL g11116 ( 
.A(n_10743),
.B(n_7348),
.Y(n_11116)
);

NAND2xp5_ASAP7_75t_L g11117 ( 
.A(n_10654),
.B(n_7227),
.Y(n_11117)
);

INVx2_ASAP7_75t_SL g11118 ( 
.A(n_10342),
.Y(n_11118)
);

NAND2xp33_ASAP7_75t_SL g11119 ( 
.A(n_10675),
.B(n_7351),
.Y(n_11119)
);

AND2x2_ASAP7_75t_L g11120 ( 
.A(n_10598),
.B(n_7355),
.Y(n_11120)
);

NAND2xp5_ASAP7_75t_L g11121 ( 
.A(n_10656),
.B(n_10664),
.Y(n_11121)
);

BUFx8_ASAP7_75t_L g11122 ( 
.A(n_10408),
.Y(n_11122)
);

OR2x6_ASAP7_75t_L g11123 ( 
.A(n_10319),
.B(n_7238),
.Y(n_11123)
);

NAND2xp5_ASAP7_75t_SL g11124 ( 
.A(n_10747),
.B(n_7356),
.Y(n_11124)
);

NAND2xp5_ASAP7_75t_SL g11125 ( 
.A(n_10630),
.B(n_7358),
.Y(n_11125)
);

NAND2xp5_ASAP7_75t_SL g11126 ( 
.A(n_10630),
.B(n_7360),
.Y(n_11126)
);

NOR2xp33_ASAP7_75t_L g11127 ( 
.A(n_10462),
.B(n_7362),
.Y(n_11127)
);

NAND2xp5_ASAP7_75t_L g11128 ( 
.A(n_10672),
.B(n_7248),
.Y(n_11128)
);

NAND2xp5_ASAP7_75t_L g11129 ( 
.A(n_10711),
.B(n_7249),
.Y(n_11129)
);

NOR2xp67_ASAP7_75t_L g11130 ( 
.A(n_10687),
.B(n_4556),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_L g11131 ( 
.A(n_10712),
.B(n_7250),
.Y(n_11131)
);

INVxp67_ASAP7_75t_L g11132 ( 
.A(n_10408),
.Y(n_11132)
);

AOI221xp5_ASAP7_75t_L g11133 ( 
.A1(n_10514),
.A2(n_7263),
.B1(n_7276),
.B2(n_7257),
.C(n_7252),
.Y(n_11133)
);

NOR2xp33_ASAP7_75t_L g11134 ( 
.A(n_10733),
.B(n_7364),
.Y(n_11134)
);

NAND2xp5_ASAP7_75t_L g11135 ( 
.A(n_10715),
.B(n_7277),
.Y(n_11135)
);

NAND2xp5_ASAP7_75t_L g11136 ( 
.A(n_10632),
.B(n_7286),
.Y(n_11136)
);

AOI22xp33_ASAP7_75t_L g11137 ( 
.A1(n_10734),
.A2(n_10740),
.B1(n_10762),
.B2(n_10704),
.Y(n_11137)
);

INVx2_ASAP7_75t_L g11138 ( 
.A(n_10536),
.Y(n_11138)
);

NAND2xp33_ASAP7_75t_L g11139 ( 
.A(n_10699),
.B(n_7373),
.Y(n_11139)
);

OR2x6_ASAP7_75t_L g11140 ( 
.A(n_10555),
.B(n_7289),
.Y(n_11140)
);

INVx1_ASAP7_75t_L g11141 ( 
.A(n_10746),
.Y(n_11141)
);

NAND2xp5_ASAP7_75t_L g11142 ( 
.A(n_10637),
.B(n_7300),
.Y(n_11142)
);

INVx1_ASAP7_75t_L g11143 ( 
.A(n_10713),
.Y(n_11143)
);

NOR2xp33_ASAP7_75t_L g11144 ( 
.A(n_10714),
.B(n_7375),
.Y(n_11144)
);

INVx2_ASAP7_75t_SL g11145 ( 
.A(n_10413),
.Y(n_11145)
);

INVx2_ASAP7_75t_L g11146 ( 
.A(n_10748),
.Y(n_11146)
);

NOR2xp33_ASAP7_75t_L g11147 ( 
.A(n_10330),
.B(n_7380),
.Y(n_11147)
);

INVx2_ASAP7_75t_L g11148 ( 
.A(n_10752),
.Y(n_11148)
);

OAI22xp33_ASAP7_75t_L g11149 ( 
.A1(n_10390),
.A2(n_10470),
.B1(n_10556),
.B2(n_10728),
.Y(n_11149)
);

NAND2xp5_ASAP7_75t_SL g11150 ( 
.A(n_10413),
.B(n_10430),
.Y(n_11150)
);

INVx2_ASAP7_75t_SL g11151 ( 
.A(n_10430),
.Y(n_11151)
);

BUFx6f_ASAP7_75t_L g11152 ( 
.A(n_10435),
.Y(n_11152)
);

INVx1_ASAP7_75t_L g11153 ( 
.A(n_10620),
.Y(n_11153)
);

NOR2xp33_ASAP7_75t_L g11154 ( 
.A(n_10479),
.B(n_7383),
.Y(n_11154)
);

NAND2xp5_ASAP7_75t_SL g11155 ( 
.A(n_10435),
.B(n_7389),
.Y(n_11155)
);

INVx2_ASAP7_75t_L g11156 ( 
.A(n_10681),
.Y(n_11156)
);

NAND2xp5_ASAP7_75t_L g11157 ( 
.A(n_10642),
.B(n_7301),
.Y(n_11157)
);

INVx1_ASAP7_75t_L g11158 ( 
.A(n_10655),
.Y(n_11158)
);

NAND2xp33_ASAP7_75t_L g11159 ( 
.A(n_10744),
.B(n_7394),
.Y(n_11159)
);

HB1xp67_ASAP7_75t_L g11160 ( 
.A(n_10373),
.Y(n_11160)
);

INVx2_ASAP7_75t_SL g11161 ( 
.A(n_10472),
.Y(n_11161)
);

BUFx6f_ASAP7_75t_L g11162 ( 
.A(n_10472),
.Y(n_11162)
);

INVx2_ASAP7_75t_L g11163 ( 
.A(n_10757),
.Y(n_11163)
);

INVx2_ASAP7_75t_L g11164 ( 
.A(n_10595),
.Y(n_11164)
);

NAND2xp5_ASAP7_75t_L g11165 ( 
.A(n_10631),
.B(n_7305),
.Y(n_11165)
);

INVx2_ASAP7_75t_L g11166 ( 
.A(n_10605),
.Y(n_11166)
);

NOR2xp33_ASAP7_75t_L g11167 ( 
.A(n_10384),
.B(n_7395),
.Y(n_11167)
);

INVx1_ASAP7_75t_L g11168 ( 
.A(n_10628),
.Y(n_11168)
);

INVx2_ASAP7_75t_SL g11169 ( 
.A(n_10489),
.Y(n_11169)
);

INVx2_ASAP7_75t_L g11170 ( 
.A(n_10612),
.Y(n_11170)
);

INVx1_ASAP7_75t_L g11171 ( 
.A(n_10738),
.Y(n_11171)
);

INVx1_ASAP7_75t_L g11172 ( 
.A(n_10385),
.Y(n_11172)
);

INVx2_ASAP7_75t_L g11173 ( 
.A(n_10612),
.Y(n_11173)
);

BUFx2_ASAP7_75t_L g11174 ( 
.A(n_10402),
.Y(n_11174)
);

INVx2_ASAP7_75t_L g11175 ( 
.A(n_10613),
.Y(n_11175)
);

BUFx3_ASAP7_75t_L g11176 ( 
.A(n_10489),
.Y(n_11176)
);

INVx1_ASAP7_75t_SL g11177 ( 
.A(n_10498),
.Y(n_11177)
);

NAND2xp5_ASAP7_75t_L g11178 ( 
.A(n_10429),
.B(n_7307),
.Y(n_11178)
);

AOI22xp33_ASAP7_75t_L g11179 ( 
.A1(n_10762),
.A2(n_7319),
.B1(n_7321),
.B2(n_7310),
.Y(n_11179)
);

INVx3_ASAP7_75t_L g11180 ( 
.A(n_10422),
.Y(n_11180)
);

OR2x2_ASAP7_75t_L g11181 ( 
.A(n_10676),
.B(n_10677),
.Y(n_11181)
);

NAND2xp5_ASAP7_75t_SL g11182 ( 
.A(n_10498),
.B(n_7396),
.Y(n_11182)
);

NAND2xp5_ASAP7_75t_L g11183 ( 
.A(n_10710),
.B(n_7324),
.Y(n_11183)
);

NAND2xp5_ASAP7_75t_SL g11184 ( 
.A(n_10527),
.B(n_7397),
.Y(n_11184)
);

INVx2_ASAP7_75t_L g11185 ( 
.A(n_10613),
.Y(n_11185)
);

NAND2xp5_ASAP7_75t_L g11186 ( 
.A(n_10717),
.B(n_7328),
.Y(n_11186)
);

INVx1_ASAP7_75t_L g11187 ( 
.A(n_10673),
.Y(n_11187)
);

AOI22xp33_ASAP7_75t_L g11188 ( 
.A1(n_10423),
.A2(n_7329),
.B1(n_7335),
.B2(n_7333),
.Y(n_11188)
);

INVx1_ASAP7_75t_L g11189 ( 
.A(n_10718),
.Y(n_11189)
);

INVx1_ASAP7_75t_L g11190 ( 
.A(n_10720),
.Y(n_11190)
);

AOI22xp33_ASAP7_75t_L g11191 ( 
.A1(n_10438),
.A2(n_7336),
.B1(n_7343),
.B2(n_7340),
.Y(n_11191)
);

NAND2xp5_ASAP7_75t_L g11192 ( 
.A(n_10723),
.B(n_7352),
.Y(n_11192)
);

OAI22xp5_ASAP7_75t_L g11193 ( 
.A1(n_10668),
.A2(n_7406),
.B1(n_7407),
.B2(n_7398),
.Y(n_11193)
);

NAND2xp5_ASAP7_75t_L g11194 ( 
.A(n_10741),
.B(n_10301),
.Y(n_11194)
);

NAND2xp5_ASAP7_75t_L g11195 ( 
.A(n_10759),
.B(n_7354),
.Y(n_11195)
);

BUFx8_ASAP7_75t_L g11196 ( 
.A(n_10527),
.Y(n_11196)
);

NAND2xp5_ASAP7_75t_SL g11197 ( 
.A(n_10540),
.B(n_7410),
.Y(n_11197)
);

INVx1_ASAP7_75t_L g11198 ( 
.A(n_10619),
.Y(n_11198)
);

NOR2xp33_ASAP7_75t_SL g11199 ( 
.A(n_10326),
.B(n_7411),
.Y(n_11199)
);

NAND2xp5_ASAP7_75t_L g11200 ( 
.A(n_10731),
.B(n_7363),
.Y(n_11200)
);

NAND2xp33_ASAP7_75t_L g11201 ( 
.A(n_10744),
.B(n_7412),
.Y(n_11201)
);

INVx4_ASAP7_75t_L g11202 ( 
.A(n_10540),
.Y(n_11202)
);

NOR2xp33_ASAP7_75t_L g11203 ( 
.A(n_10456),
.B(n_7413),
.Y(n_11203)
);

NAND2xp5_ASAP7_75t_L g11204 ( 
.A(n_10751),
.B(n_7368),
.Y(n_11204)
);

INVx2_ASAP7_75t_L g11205 ( 
.A(n_10695),
.Y(n_11205)
);

NOR2xp33_ASAP7_75t_L g11206 ( 
.A(n_10320),
.B(n_7417),
.Y(n_11206)
);

INVx1_ASAP7_75t_L g11207 ( 
.A(n_10707),
.Y(n_11207)
);

OAI221xp5_ASAP7_75t_L g11208 ( 
.A1(n_10412),
.A2(n_7374),
.B1(n_7376),
.B2(n_7370),
.C(n_7369),
.Y(n_11208)
);

INVx3_ASAP7_75t_L g11209 ( 
.A(n_10440),
.Y(n_11209)
);

HB1xp67_ASAP7_75t_L g11210 ( 
.A(n_10303),
.Y(n_11210)
);

BUFx3_ASAP7_75t_L g11211 ( 
.A(n_10282),
.Y(n_11211)
);

NAND2xp5_ASAP7_75t_L g11212 ( 
.A(n_10395),
.B(n_7377),
.Y(n_11212)
);

NOR2xp33_ASAP7_75t_L g11213 ( 
.A(n_10491),
.B(n_7418),
.Y(n_11213)
);

NAND2xp33_ASAP7_75t_L g11214 ( 
.A(n_10697),
.B(n_10700),
.Y(n_11214)
);

INVx1_ASAP7_75t_L g11215 ( 
.A(n_10685),
.Y(n_11215)
);

NAND2xp5_ASAP7_75t_L g11216 ( 
.A(n_10616),
.B(n_7379),
.Y(n_11216)
);

INVx1_ASAP7_75t_L g11217 ( 
.A(n_10685),
.Y(n_11217)
);

BUFx6f_ASAP7_75t_L g11218 ( 
.A(n_10551),
.Y(n_11218)
);

NAND2xp5_ASAP7_75t_L g11219 ( 
.A(n_10758),
.B(n_10439),
.Y(n_11219)
);

INVx1_ASAP7_75t_L g11220 ( 
.A(n_10669),
.Y(n_11220)
);

INVx1_ASAP7_75t_L g11221 ( 
.A(n_10434),
.Y(n_11221)
);

NAND2xp5_ASAP7_75t_L g11222 ( 
.A(n_10625),
.B(n_7381),
.Y(n_11222)
);

INVx1_ASAP7_75t_L g11223 ( 
.A(n_10476),
.Y(n_11223)
);

NAND2xp5_ASAP7_75t_SL g11224 ( 
.A(n_10419),
.B(n_7420),
.Y(n_11224)
);

OAI22xp5_ASAP7_75t_L g11225 ( 
.A1(n_10610),
.A2(n_7422),
.B1(n_7423),
.B2(n_7421),
.Y(n_11225)
);

BUFx6f_ASAP7_75t_L g11226 ( 
.A(n_10551),
.Y(n_11226)
);

INVxp67_ASAP7_75t_SL g11227 ( 
.A(n_10418),
.Y(n_11227)
);

INVx2_ASAP7_75t_L g11228 ( 
.A(n_10608),
.Y(n_11228)
);

INVx2_ASAP7_75t_L g11229 ( 
.A(n_10508),
.Y(n_11229)
);

NAND2xp5_ASAP7_75t_L g11230 ( 
.A(n_10486),
.B(n_7387),
.Y(n_11230)
);

NAND2xp5_ASAP7_75t_L g11231 ( 
.A(n_10503),
.B(n_7390),
.Y(n_11231)
);

NOR3xp33_ASAP7_75t_L g11232 ( 
.A(n_10522),
.B(n_7401),
.C(n_7392),
.Y(n_11232)
);

INVx2_ASAP7_75t_SL g11233 ( 
.A(n_10560),
.Y(n_11233)
);

NAND2xp5_ASAP7_75t_L g11234 ( 
.A(n_10539),
.B(n_7402),
.Y(n_11234)
);

INVx1_ASAP7_75t_L g11235 ( 
.A(n_10515),
.Y(n_11235)
);

INVx2_ASAP7_75t_L g11236 ( 
.A(n_10431),
.Y(n_11236)
);

AOI22xp33_ASAP7_75t_L g11237 ( 
.A1(n_10559),
.A2(n_7405),
.B1(n_7414),
.B2(n_7404),
.Y(n_11237)
);

A2O1A1Ixp33_ASAP7_75t_L g11238 ( 
.A1(n_10512),
.A2(n_7439),
.B(n_7449),
.C(n_7424),
.Y(n_11238)
);

OR2x2_ASAP7_75t_L g11239 ( 
.A(n_10334),
.B(n_7426),
.Y(n_11239)
);

INVx2_ASAP7_75t_L g11240 ( 
.A(n_10560),
.Y(n_11240)
);

INVx1_ASAP7_75t_L g11241 ( 
.A(n_10696),
.Y(n_11241)
);

INVxp67_ASAP7_75t_SL g11242 ( 
.A(n_10570),
.Y(n_11242)
);

NOR2xp33_ASAP7_75t_L g11243 ( 
.A(n_10574),
.B(n_7428),
.Y(n_11243)
);

A2O1A1Ixp33_ASAP7_75t_L g11244 ( 
.A1(n_10593),
.A2(n_7459),
.B(n_7466),
.C(n_7450),
.Y(n_11244)
);

INVx1_ASAP7_75t_L g11245 ( 
.A(n_10709),
.Y(n_11245)
);

NAND2xp5_ASAP7_75t_L g11246 ( 
.A(n_10487),
.B(n_7467),
.Y(n_11246)
);

INVx1_ASAP7_75t_L g11247 ( 
.A(n_10289),
.Y(n_11247)
);

NAND2xp5_ASAP7_75t_L g11248 ( 
.A(n_10559),
.B(n_7468),
.Y(n_11248)
);

INVx1_ASAP7_75t_SL g11249 ( 
.A(n_10295),
.Y(n_11249)
);

NAND2xp5_ASAP7_75t_SL g11250 ( 
.A(n_10432),
.B(n_7431),
.Y(n_11250)
);

NAND2xp5_ASAP7_75t_L g11251 ( 
.A(n_10571),
.B(n_7470),
.Y(n_11251)
);

NOR2xp67_ASAP7_75t_L g11252 ( 
.A(n_10578),
.B(n_4557),
.Y(n_11252)
);

NAND2xp5_ASAP7_75t_L g11253 ( 
.A(n_10571),
.B(n_7471),
.Y(n_11253)
);

AOI22xp5_ASAP7_75t_L g11254 ( 
.A1(n_10351),
.A2(n_7434),
.B1(n_7435),
.B2(n_7433),
.Y(n_11254)
);

OAI22xp5_ASAP7_75t_L g11255 ( 
.A1(n_10622),
.A2(n_7442),
.B1(n_7443),
.B2(n_7441),
.Y(n_11255)
);

NAND2xp5_ASAP7_75t_SL g11256 ( 
.A(n_10549),
.B(n_10570),
.Y(n_11256)
);

NOR2xp67_ASAP7_75t_L g11257 ( 
.A(n_10447),
.B(n_10312),
.Y(n_11257)
);

INVx1_ASAP7_75t_L g11258 ( 
.A(n_10596),
.Y(n_11258)
);

INVx2_ASAP7_75t_SL g11259 ( 
.A(n_10596),
.Y(n_11259)
);

INVx1_ASAP7_75t_L g11260 ( 
.A(n_10311),
.Y(n_11260)
);

INVxp67_ASAP7_75t_L g11261 ( 
.A(n_10561),
.Y(n_11261)
);

INVx2_ASAP7_75t_L g11262 ( 
.A(n_10565),
.Y(n_11262)
);

INVx2_ASAP7_75t_L g11263 ( 
.A(n_10591),
.Y(n_11263)
);

INVx1_ASAP7_75t_L g11264 ( 
.A(n_10362),
.Y(n_11264)
);

OR2x2_ASAP7_75t_L g11265 ( 
.A(n_10415),
.B(n_7444),
.Y(n_11265)
);

NAND2xp5_ASAP7_75t_L g11266 ( 
.A(n_10648),
.B(n_7480),
.Y(n_11266)
);

INVx1_ASAP7_75t_L g11267 ( 
.A(n_10531),
.Y(n_11267)
);

OR2x2_ASAP7_75t_L g11268 ( 
.A(n_10599),
.B(n_7446),
.Y(n_11268)
);

INVx2_ASAP7_75t_L g11269 ( 
.A(n_10692),
.Y(n_11269)
);

NAND2xp5_ASAP7_75t_SL g11270 ( 
.A(n_10325),
.B(n_7447),
.Y(n_11270)
);

NAND2xp5_ASAP7_75t_L g11271 ( 
.A(n_10648),
.B(n_7482),
.Y(n_11271)
);

NOR2xp33_ASAP7_75t_L g11272 ( 
.A(n_10382),
.B(n_7448),
.Y(n_11272)
);

INVx1_ASAP7_75t_L g11273 ( 
.A(n_10569),
.Y(n_11273)
);

INVxp67_ASAP7_75t_L g11274 ( 
.A(n_10650),
.Y(n_11274)
);

NAND2xp5_ASAP7_75t_L g11275 ( 
.A(n_10650),
.B(n_7485),
.Y(n_11275)
);

INVx1_ASAP7_75t_L g11276 ( 
.A(n_10537),
.Y(n_11276)
);

NAND2xp5_ASAP7_75t_L g11277 ( 
.A(n_10406),
.B(n_10397),
.Y(n_11277)
);

NAND2xp5_ASAP7_75t_SL g11278 ( 
.A(n_10396),
.B(n_10391),
.Y(n_11278)
);

NAND2xp5_ASAP7_75t_L g11279 ( 
.A(n_10406),
.B(n_7497),
.Y(n_11279)
);

BUFx12f_ASAP7_75t_L g11280 ( 
.A(n_10339),
.Y(n_11280)
);

INVx2_ASAP7_75t_L g11281 ( 
.A(n_10397),
.Y(n_11281)
);

NAND2xp5_ASAP7_75t_L g11282 ( 
.A(n_10393),
.B(n_7500),
.Y(n_11282)
);

INVx2_ASAP7_75t_L g11283 ( 
.A(n_10327),
.Y(n_11283)
);

NAND2xp5_ASAP7_75t_L g11284 ( 
.A(n_10499),
.B(n_7501),
.Y(n_11284)
);

AND2x6_ASAP7_75t_SL g11285 ( 
.A(n_10266),
.B(n_7509),
.Y(n_11285)
);

INVx1_ASAP7_75t_L g11286 ( 
.A(n_10255),
.Y(n_11286)
);

INVx1_ASAP7_75t_L g11287 ( 
.A(n_10926),
.Y(n_11287)
);

INVxp67_ASAP7_75t_L g11288 ( 
.A(n_10787),
.Y(n_11288)
);

AND2x2_ASAP7_75t_L g11289 ( 
.A(n_10812),
.B(n_7510),
.Y(n_11289)
);

INVx1_ASAP7_75t_L g11290 ( 
.A(n_11040),
.Y(n_11290)
);

INVx1_ASAP7_75t_L g11291 ( 
.A(n_10789),
.Y(n_11291)
);

INVx1_ASAP7_75t_L g11292 ( 
.A(n_10791),
.Y(n_11292)
);

AOI22xp5_ASAP7_75t_L g11293 ( 
.A1(n_11032),
.A2(n_10801),
.B1(n_11010),
.B2(n_10909),
.Y(n_11293)
);

NOR2xp33_ASAP7_75t_L g11294 ( 
.A(n_10775),
.B(n_7452),
.Y(n_11294)
);

AOI22xp5_ASAP7_75t_L g11295 ( 
.A1(n_10823),
.A2(n_7454),
.B1(n_7457),
.B2(n_7453),
.Y(n_11295)
);

INVx1_ASAP7_75t_L g11296 ( 
.A(n_10795),
.Y(n_11296)
);

INVx1_ASAP7_75t_L g11297 ( 
.A(n_10805),
.Y(n_11297)
);

INVx1_ASAP7_75t_L g11298 ( 
.A(n_10809),
.Y(n_11298)
);

AO22x2_ASAP7_75t_L g11299 ( 
.A1(n_10764),
.A2(n_7512),
.B1(n_7342),
.B2(n_7347),
.Y(n_11299)
);

INVx1_ASAP7_75t_L g11300 ( 
.A(n_10833),
.Y(n_11300)
);

INVx1_ASAP7_75t_L g11301 ( 
.A(n_10838),
.Y(n_11301)
);

INVx1_ASAP7_75t_L g11302 ( 
.A(n_10844),
.Y(n_11302)
);

NOR2xp33_ASAP7_75t_L g11303 ( 
.A(n_10781),
.B(n_7465),
.Y(n_11303)
);

OAI22xp5_ASAP7_75t_L g11304 ( 
.A1(n_10774),
.A2(n_7474),
.B1(n_7475),
.B2(n_7472),
.Y(n_11304)
);

INVx1_ASAP7_75t_L g11305 ( 
.A(n_10853),
.Y(n_11305)
);

AOI22xp5_ASAP7_75t_L g11306 ( 
.A1(n_10834),
.A2(n_7484),
.B1(n_7488),
.B2(n_7483),
.Y(n_11306)
);

NAND2xp5_ASAP7_75t_L g11307 ( 
.A(n_11004),
.B(n_7489),
.Y(n_11307)
);

NAND2xp5_ASAP7_75t_L g11308 ( 
.A(n_10931),
.B(n_7492),
.Y(n_11308)
);

AO22x2_ASAP7_75t_L g11309 ( 
.A1(n_10811),
.A2(n_7353),
.B1(n_7427),
.B2(n_7326),
.Y(n_11309)
);

INVx1_ASAP7_75t_L g11310 ( 
.A(n_10867),
.Y(n_11310)
);

INVx2_ASAP7_75t_L g11311 ( 
.A(n_10888),
.Y(n_11311)
);

INVx1_ASAP7_75t_L g11312 ( 
.A(n_10920),
.Y(n_11312)
);

NAND2x1p5_ASAP7_75t_L g11313 ( 
.A(n_10856),
.B(n_7438),
.Y(n_11313)
);

AO22x2_ASAP7_75t_L g11314 ( 
.A1(n_10773),
.A2(n_7514),
.B1(n_7530),
.B2(n_7502),
.Y(n_11314)
);

INVx1_ASAP7_75t_L g11315 ( 
.A(n_10936),
.Y(n_11315)
);

INVx3_ASAP7_75t_L g11316 ( 
.A(n_10960),
.Y(n_11316)
);

AO22x2_ASAP7_75t_L g11317 ( 
.A1(n_11219),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_11317)
);

INVx1_ASAP7_75t_L g11318 ( 
.A(n_10938),
.Y(n_11318)
);

INVx1_ASAP7_75t_L g11319 ( 
.A(n_10940),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_10941),
.Y(n_11320)
);

INVx1_ASAP7_75t_L g11321 ( 
.A(n_10944),
.Y(n_11321)
);

AND2x4_ASAP7_75t_L g11322 ( 
.A(n_10808),
.B(n_4558),
.Y(n_11322)
);

BUFx8_ASAP7_75t_L g11323 ( 
.A(n_11027),
.Y(n_11323)
);

NAND2x1p5_ASAP7_75t_L g11324 ( 
.A(n_10817),
.B(n_4560),
.Y(n_11324)
);

AO22x2_ASAP7_75t_L g11325 ( 
.A1(n_10912),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_11325)
);

NAND2xp5_ASAP7_75t_SL g11326 ( 
.A(n_11181),
.B(n_7498),
.Y(n_11326)
);

INVx1_ASAP7_75t_L g11327 ( 
.A(n_10947),
.Y(n_11327)
);

NAND2xp5_ASAP7_75t_L g11328 ( 
.A(n_10878),
.B(n_7503),
.Y(n_11328)
);

INVx1_ASAP7_75t_L g11329 ( 
.A(n_10954),
.Y(n_11329)
);

INVx2_ASAP7_75t_L g11330 ( 
.A(n_10962),
.Y(n_11330)
);

AND2x4_ASAP7_75t_L g11331 ( 
.A(n_11082),
.B(n_4561),
.Y(n_11331)
);

AO22x2_ASAP7_75t_L g11332 ( 
.A1(n_11236),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_11332)
);

NAND2xp5_ASAP7_75t_L g11333 ( 
.A(n_11189),
.B(n_7504),
.Y(n_11333)
);

AND2x4_ASAP7_75t_L g11334 ( 
.A(n_11088),
.B(n_4562),
.Y(n_11334)
);

NAND2xp5_ASAP7_75t_L g11335 ( 
.A(n_11190),
.B(n_7508),
.Y(n_11335)
);

BUFx8_ASAP7_75t_L g11336 ( 
.A(n_10771),
.Y(n_11336)
);

NAND2xp5_ASAP7_75t_SL g11337 ( 
.A(n_10783),
.B(n_7511),
.Y(n_11337)
);

NAND2xp5_ASAP7_75t_L g11338 ( 
.A(n_11061),
.B(n_11158),
.Y(n_11338)
);

AO22x2_ASAP7_75t_L g11339 ( 
.A1(n_10829),
.A2(n_10782),
.B1(n_11022),
.B2(n_10980),
.Y(n_11339)
);

NAND2x1p5_ASAP7_75t_L g11340 ( 
.A(n_10771),
.B(n_4564),
.Y(n_11340)
);

AO22x2_ASAP7_75t_L g11341 ( 
.A1(n_10850),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_11341)
);

CKINVDCx5p33_ASAP7_75t_R g11342 ( 
.A(n_10828),
.Y(n_11342)
);

NAND2x1p5_ASAP7_75t_L g11343 ( 
.A(n_10776),
.B(n_4565),
.Y(n_11343)
);

INVx1_ASAP7_75t_L g11344 ( 
.A(n_10965),
.Y(n_11344)
);

NAND2x1p5_ASAP7_75t_L g11345 ( 
.A(n_11174),
.B(n_4567),
.Y(n_11345)
);

NAND2xp5_ASAP7_75t_L g11346 ( 
.A(n_10810),
.B(n_10882),
.Y(n_11346)
);

INVx1_ASAP7_75t_L g11347 ( 
.A(n_10967),
.Y(n_11347)
);

INVx1_ASAP7_75t_L g11348 ( 
.A(n_10968),
.Y(n_11348)
);

AO22x2_ASAP7_75t_L g11349 ( 
.A1(n_10799),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_11349)
);

AND2x4_ASAP7_75t_L g11350 ( 
.A(n_10933),
.B(n_4568),
.Y(n_11350)
);

INVxp67_ASAP7_75t_L g11351 ( 
.A(n_11026),
.Y(n_11351)
);

HB1xp67_ASAP7_75t_L g11352 ( 
.A(n_10903),
.Y(n_11352)
);

INVxp67_ASAP7_75t_L g11353 ( 
.A(n_11160),
.Y(n_11353)
);

BUFx2_ASAP7_75t_L g11354 ( 
.A(n_10772),
.Y(n_11354)
);

INVx1_ASAP7_75t_L g11355 ( 
.A(n_10767),
.Y(n_11355)
);

INVx1_ASAP7_75t_L g11356 ( 
.A(n_10777),
.Y(n_11356)
);

INVx1_ASAP7_75t_L g11357 ( 
.A(n_10780),
.Y(n_11357)
);

NAND2xp5_ASAP7_75t_SL g11358 ( 
.A(n_10807),
.B(n_7515),
.Y(n_11358)
);

INVx1_ASAP7_75t_L g11359 ( 
.A(n_10788),
.Y(n_11359)
);

INVx1_ASAP7_75t_L g11360 ( 
.A(n_10802),
.Y(n_11360)
);

CKINVDCx5p33_ASAP7_75t_R g11361 ( 
.A(n_11122),
.Y(n_11361)
);

OR2x2_ASAP7_75t_SL g11362 ( 
.A(n_11277),
.B(n_7519),
.Y(n_11362)
);

NAND2xp5_ASAP7_75t_L g11363 ( 
.A(n_10889),
.B(n_7522),
.Y(n_11363)
);

NAND2x1p5_ASAP7_75t_L g11364 ( 
.A(n_11202),
.B(n_10950),
.Y(n_11364)
);

AND2x2_ASAP7_75t_L g11365 ( 
.A(n_10822),
.B(n_7523),
.Y(n_11365)
);

CKINVDCx5p33_ASAP7_75t_R g11366 ( 
.A(n_11196),
.Y(n_11366)
);

INVx1_ASAP7_75t_L g11367 ( 
.A(n_10815),
.Y(n_11367)
);

NAND2xp5_ASAP7_75t_L g11368 ( 
.A(n_10994),
.B(n_7525),
.Y(n_11368)
);

INVx1_ASAP7_75t_L g11369 ( 
.A(n_10825),
.Y(n_11369)
);

BUFx8_ASAP7_75t_L g11370 ( 
.A(n_11218),
.Y(n_11370)
);

AOI22xp5_ASAP7_75t_L g11371 ( 
.A1(n_10908),
.A2(n_7533),
.B1(n_7539),
.B2(n_7527),
.Y(n_11371)
);

AO22x2_ASAP7_75t_L g11372 ( 
.A1(n_10857),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_11372)
);

NOR2xp33_ASAP7_75t_L g11373 ( 
.A(n_11090),
.B(n_7542),
.Y(n_11373)
);

CKINVDCx5p33_ASAP7_75t_R g11374 ( 
.A(n_11280),
.Y(n_11374)
);

NAND2xp5_ASAP7_75t_L g11375 ( 
.A(n_11284),
.B(n_7543),
.Y(n_11375)
);

INVx1_ASAP7_75t_L g11376 ( 
.A(n_10827),
.Y(n_11376)
);

AO22x2_ASAP7_75t_L g11377 ( 
.A1(n_11138),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_11377)
);

AO22x2_ASAP7_75t_L g11378 ( 
.A1(n_10786),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_11378)
);

OAI221xp5_ASAP7_75t_L g11379 ( 
.A1(n_11011),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.C(n_28),
.Y(n_11379)
);

OAI221xp5_ASAP7_75t_L g11380 ( 
.A1(n_10863),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.C(n_31),
.Y(n_11380)
);

AO22x2_ASAP7_75t_L g11381 ( 
.A1(n_11215),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_11381)
);

CKINVDCx5p33_ASAP7_75t_R g11382 ( 
.A(n_10770),
.Y(n_11382)
);

INVx1_ASAP7_75t_L g11383 ( 
.A(n_10845),
.Y(n_11383)
);

AOI22xp5_ASAP7_75t_SL g11384 ( 
.A1(n_10837),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_11384)
);

CKINVDCx5p33_ASAP7_75t_R g11385 ( 
.A(n_10999),
.Y(n_11385)
);

INVx2_ASAP7_75t_L g11386 ( 
.A(n_10900),
.Y(n_11386)
);

INVx1_ASAP7_75t_L g11387 ( 
.A(n_10859),
.Y(n_11387)
);

NAND2x1p5_ASAP7_75t_L g11388 ( 
.A(n_11031),
.B(n_4569),
.Y(n_11388)
);

INVxp67_ASAP7_75t_L g11389 ( 
.A(n_11210),
.Y(n_11389)
);

INVx2_ASAP7_75t_L g11390 ( 
.A(n_10902),
.Y(n_11390)
);

AOI22xp5_ASAP7_75t_L g11391 ( 
.A1(n_11213),
.A2(n_10964),
.B1(n_11149),
.B2(n_10991),
.Y(n_11391)
);

AND2x2_ASAP7_75t_L g11392 ( 
.A(n_10983),
.B(n_33),
.Y(n_11392)
);

INVx1_ASAP7_75t_L g11393 ( 
.A(n_10865),
.Y(n_11393)
);

CKINVDCx5p33_ASAP7_75t_R g11394 ( 
.A(n_10999),
.Y(n_11394)
);

INVx2_ASAP7_75t_L g11395 ( 
.A(n_10913),
.Y(n_11395)
);

HB1xp67_ASAP7_75t_L g11396 ( 
.A(n_10790),
.Y(n_11396)
);

INVx1_ASAP7_75t_L g11397 ( 
.A(n_10866),
.Y(n_11397)
);

AO22x2_ASAP7_75t_L g11398 ( 
.A1(n_11217),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_11398)
);

AO22x2_ASAP7_75t_L g11399 ( 
.A1(n_11064),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_11399)
);

INVx1_ASAP7_75t_L g11400 ( 
.A(n_10873),
.Y(n_11400)
);

AO22x2_ASAP7_75t_L g11401 ( 
.A1(n_11107),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_11401)
);

NOR2xp67_ASAP7_75t_L g11402 ( 
.A(n_10803),
.B(n_4571),
.Y(n_11402)
);

INVx2_ASAP7_75t_L g11403 ( 
.A(n_10916),
.Y(n_11403)
);

AO22x2_ASAP7_75t_L g11404 ( 
.A1(n_10765),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_11404)
);

INVx2_ASAP7_75t_L g11405 ( 
.A(n_10977),
.Y(n_11405)
);

AOI22xp5_ASAP7_75t_L g11406 ( 
.A1(n_10943),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_11406)
);

AND2x4_ASAP7_75t_L g11407 ( 
.A(n_11242),
.B(n_11211),
.Y(n_11407)
);

AOI22xp33_ASAP7_75t_L g11408 ( 
.A1(n_11099),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_11408)
);

INVx1_ASAP7_75t_L g11409 ( 
.A(n_10894),
.Y(n_11409)
);

AOI22xp5_ASAP7_75t_L g11410 ( 
.A1(n_10985),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_11410)
);

AOI22xp5_ASAP7_75t_L g11411 ( 
.A1(n_11147),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_11411)
);

INVx1_ASAP7_75t_L g11412 ( 
.A(n_10895),
.Y(n_11412)
);

INVx1_ASAP7_75t_L g11413 ( 
.A(n_10896),
.Y(n_11413)
);

AO22x2_ASAP7_75t_L g11414 ( 
.A1(n_10784),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_11414)
);

INVx1_ASAP7_75t_L g11415 ( 
.A(n_10899),
.Y(n_11415)
);

OAI221xp5_ASAP7_75t_L g11416 ( 
.A1(n_10869),
.A2(n_10911),
.B1(n_10969),
.B2(n_10959),
.C(n_11127),
.Y(n_11416)
);

NOR2xp33_ASAP7_75t_L g11417 ( 
.A(n_10816),
.B(n_4572),
.Y(n_11417)
);

NAND2xp5_ASAP7_75t_L g11418 ( 
.A(n_10818),
.B(n_49),
.Y(n_11418)
);

INVx2_ASAP7_75t_L g11419 ( 
.A(n_11006),
.Y(n_11419)
);

OAI221xp5_ASAP7_75t_L g11420 ( 
.A1(n_11237),
.A2(n_10830),
.B1(n_11070),
.B2(n_11179),
.C(n_11038),
.Y(n_11420)
);

AOI22xp5_ASAP7_75t_L g11421 ( 
.A1(n_10824),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_11421)
);

AND2x2_ASAP7_75t_L g11422 ( 
.A(n_10885),
.B(n_50),
.Y(n_11422)
);

INVx2_ASAP7_75t_L g11423 ( 
.A(n_11013),
.Y(n_11423)
);

INVx2_ASAP7_75t_L g11424 ( 
.A(n_11050),
.Y(n_11424)
);

AOI22xp5_ASAP7_75t_L g11425 ( 
.A1(n_10832),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_11425)
);

AND2x2_ASAP7_75t_L g11426 ( 
.A(n_10995),
.B(n_10793),
.Y(n_11426)
);

AND2x4_ASAP7_75t_L g11427 ( 
.A(n_11262),
.B(n_4573),
.Y(n_11427)
);

AND2x4_ASAP7_75t_L g11428 ( 
.A(n_11263),
.B(n_4574),
.Y(n_11428)
);

BUFx2_ASAP7_75t_L g11429 ( 
.A(n_11132),
.Y(n_11429)
);

AO22x2_ASAP7_75t_L g11430 ( 
.A1(n_10814),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_11430)
);

INVx1_ASAP7_75t_L g11431 ( 
.A(n_10919),
.Y(n_11431)
);

NAND2xp33_ASAP7_75t_L g11432 ( 
.A(n_10897),
.B(n_54),
.Y(n_11432)
);

INVx1_ASAP7_75t_L g11433 ( 
.A(n_10923),
.Y(n_11433)
);

AO22x2_ASAP7_75t_L g11434 ( 
.A1(n_10942),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_11434)
);

INVxp67_ASAP7_75t_L g11435 ( 
.A(n_10769),
.Y(n_11435)
);

NAND2xp5_ASAP7_75t_L g11436 ( 
.A(n_10820),
.B(n_56),
.Y(n_11436)
);

INVx2_ASAP7_75t_L g11437 ( 
.A(n_11054),
.Y(n_11437)
);

AND2x4_ASAP7_75t_L g11438 ( 
.A(n_11233),
.B(n_4575),
.Y(n_11438)
);

NAND2xp5_ASAP7_75t_SL g11439 ( 
.A(n_10915),
.B(n_57),
.Y(n_11439)
);

AO22x2_ASAP7_75t_L g11440 ( 
.A1(n_11273),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_11440)
);

NOR2xp67_ASAP7_75t_L g11441 ( 
.A(n_10990),
.B(n_4576),
.Y(n_11441)
);

NAND2x1p5_ASAP7_75t_L g11442 ( 
.A(n_11068),
.B(n_4577),
.Y(n_11442)
);

INVx1_ASAP7_75t_L g11443 ( 
.A(n_10925),
.Y(n_11443)
);

INVx1_ASAP7_75t_L g11444 ( 
.A(n_10946),
.Y(n_11444)
);

BUFx8_ASAP7_75t_L g11445 ( 
.A(n_11218),
.Y(n_11445)
);

INVx1_ASAP7_75t_L g11446 ( 
.A(n_10949),
.Y(n_11446)
);

AOI22xp5_ASAP7_75t_L g11447 ( 
.A1(n_11272),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_11447)
);

INVx1_ASAP7_75t_L g11448 ( 
.A(n_10955),
.Y(n_11448)
);

INVx2_ASAP7_75t_L g11449 ( 
.A(n_11055),
.Y(n_11449)
);

AO22x2_ASAP7_75t_L g11450 ( 
.A1(n_11212),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_11450)
);

AO22x2_ASAP7_75t_L g11451 ( 
.A1(n_11194),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_11451)
);

INVx1_ASAP7_75t_L g11452 ( 
.A(n_10956),
.Y(n_11452)
);

NAND2x1p5_ASAP7_75t_L g11453 ( 
.A(n_11180),
.B(n_4578),
.Y(n_11453)
);

INVx1_ASAP7_75t_L g11454 ( 
.A(n_10957),
.Y(n_11454)
);

INVx1_ASAP7_75t_L g11455 ( 
.A(n_10971),
.Y(n_11455)
);

INVxp67_ASAP7_75t_L g11456 ( 
.A(n_10871),
.Y(n_11456)
);

AO22x2_ASAP7_75t_L g11457 ( 
.A1(n_10880),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_11457)
);

NAND2xp5_ASAP7_75t_L g11458 ( 
.A(n_10800),
.B(n_64),
.Y(n_11458)
);

INVx2_ASAP7_75t_L g11459 ( 
.A(n_11063),
.Y(n_11459)
);

INVx1_ASAP7_75t_L g11460 ( 
.A(n_10973),
.Y(n_11460)
);

OR2x2_ASAP7_75t_L g11461 ( 
.A(n_10766),
.B(n_65),
.Y(n_11461)
);

NOR2xp33_ASAP7_75t_L g11462 ( 
.A(n_10797),
.B(n_4580),
.Y(n_11462)
);

AO22x2_ASAP7_75t_L g11463 ( 
.A1(n_10883),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_11463)
);

INVx1_ASAP7_75t_L g11464 ( 
.A(n_11286),
.Y(n_11464)
);

AO22x2_ASAP7_75t_L g11465 ( 
.A1(n_11276),
.A2(n_70),
.B1(n_67),
.B2(n_69),
.Y(n_11465)
);

BUFx2_ASAP7_75t_L g11466 ( 
.A(n_10958),
.Y(n_11466)
);

INVx2_ASAP7_75t_L g11467 ( 
.A(n_11066),
.Y(n_11467)
);

AND2x4_ASAP7_75t_L g11468 ( 
.A(n_11259),
.B(n_4582),
.Y(n_11468)
);

INVxp67_ASAP7_75t_L g11469 ( 
.A(n_11265),
.Y(n_11469)
);

AO22x2_ASAP7_75t_L g11470 ( 
.A1(n_10855),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_11470)
);

NOR2xp33_ASAP7_75t_L g11471 ( 
.A(n_10813),
.B(n_4583),
.Y(n_11471)
);

AO22x2_ASAP7_75t_L g11472 ( 
.A1(n_10891),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_11472)
);

INVx1_ASAP7_75t_L g11473 ( 
.A(n_11036),
.Y(n_11473)
);

AO22x2_ASAP7_75t_L g11474 ( 
.A1(n_11041),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_11474)
);

INVxp67_ASAP7_75t_L g11475 ( 
.A(n_11240),
.Y(n_11475)
);

INVx2_ASAP7_75t_L g11476 ( 
.A(n_11077),
.Y(n_11476)
);

INVx2_ASAP7_75t_SL g11477 ( 
.A(n_11076),
.Y(n_11477)
);

INVx1_ASAP7_75t_L g11478 ( 
.A(n_11045),
.Y(n_11478)
);

BUFx8_ASAP7_75t_L g11479 ( 
.A(n_11226),
.Y(n_11479)
);

NAND2x1p5_ASAP7_75t_L g11480 ( 
.A(n_11209),
.B(n_4584),
.Y(n_11480)
);

NAND2xp5_ASAP7_75t_L g11481 ( 
.A(n_10876),
.B(n_74),
.Y(n_11481)
);

INVx1_ASAP7_75t_L g11482 ( 
.A(n_11053),
.Y(n_11482)
);

BUFx8_ASAP7_75t_L g11483 ( 
.A(n_11226),
.Y(n_11483)
);

AOI22xp5_ASAP7_75t_L g11484 ( 
.A1(n_10806),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_11484)
);

AO22x2_ASAP7_75t_L g11485 ( 
.A1(n_11225),
.A2(n_11255),
.B1(n_10831),
.B2(n_10796),
.Y(n_11485)
);

INVx1_ASAP7_75t_L g11486 ( 
.A(n_11046),
.Y(n_11486)
);

AO22x2_ASAP7_75t_L g11487 ( 
.A1(n_11141),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_11487)
);

INVx1_ASAP7_75t_L g11488 ( 
.A(n_11039),
.Y(n_11488)
);

OAI221xp5_ASAP7_75t_L g11489 ( 
.A1(n_11154),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.C(n_83),
.Y(n_11489)
);

INVx2_ASAP7_75t_L g11490 ( 
.A(n_11086),
.Y(n_11490)
);

AO22x2_ASAP7_75t_L g11491 ( 
.A1(n_11281),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_11491)
);

BUFx2_ASAP7_75t_L g11492 ( 
.A(n_10961),
.Y(n_11492)
);

INVx1_ASAP7_75t_L g11493 ( 
.A(n_10979),
.Y(n_11493)
);

NOR2xp67_ASAP7_75t_L g11494 ( 
.A(n_11228),
.B(n_4585),
.Y(n_11494)
);

NAND2xp5_ASAP7_75t_L g11495 ( 
.A(n_10846),
.B(n_83),
.Y(n_11495)
);

OAI22xp33_ASAP7_75t_SL g11496 ( 
.A1(n_11208),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_11496)
);

AND2x4_ASAP7_75t_L g11497 ( 
.A(n_11044),
.B(n_4586),
.Y(n_11497)
);

AO22x2_ASAP7_75t_L g11498 ( 
.A1(n_10843),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_11498)
);

INVx1_ASAP7_75t_L g11499 ( 
.A(n_10984),
.Y(n_11499)
);

CKINVDCx5p33_ASAP7_75t_R g11500 ( 
.A(n_11076),
.Y(n_11500)
);

NAND2xp5_ASAP7_75t_L g11501 ( 
.A(n_10851),
.B(n_87),
.Y(n_11501)
);

AND2x4_ASAP7_75t_L g11502 ( 
.A(n_10893),
.B(n_4587),
.Y(n_11502)
);

INVx1_ASAP7_75t_L g11503 ( 
.A(n_10986),
.Y(n_11503)
);

AO22x2_ASAP7_75t_L g11504 ( 
.A1(n_11156),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_11504)
);

INVx2_ASAP7_75t_L g11505 ( 
.A(n_11096),
.Y(n_11505)
);

INVx1_ASAP7_75t_L g11506 ( 
.A(n_10989),
.Y(n_11506)
);

A2O1A1Ixp33_ASAP7_75t_L g11507 ( 
.A1(n_11167),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_11507)
);

INVx1_ASAP7_75t_L g11508 ( 
.A(n_10993),
.Y(n_11508)
);

BUFx8_ASAP7_75t_L g11509 ( 
.A(n_11283),
.Y(n_11509)
);

INVx1_ASAP7_75t_L g11510 ( 
.A(n_11000),
.Y(n_11510)
);

INVx1_ASAP7_75t_L g11511 ( 
.A(n_11002),
.Y(n_11511)
);

OA22x2_ASAP7_75t_L g11512 ( 
.A1(n_10997),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_11512)
);

AOI22xp5_ASAP7_75t_SL g11513 ( 
.A1(n_11274),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_11513)
);

AND2x2_ASAP7_75t_L g11514 ( 
.A(n_11074),
.B(n_94),
.Y(n_11514)
);

INVx1_ASAP7_75t_L g11515 ( 
.A(n_11012),
.Y(n_11515)
);

INVx1_ASAP7_75t_L g11516 ( 
.A(n_11067),
.Y(n_11516)
);

AO22x2_ASAP7_75t_L g11517 ( 
.A1(n_10996),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_11517)
);

AND2x2_ASAP7_75t_SL g11518 ( 
.A(n_10778),
.B(n_95),
.Y(n_11518)
);

OAI221xp5_ASAP7_75t_L g11519 ( 
.A1(n_11203),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.C(n_99),
.Y(n_11519)
);

INVx1_ASAP7_75t_L g11520 ( 
.A(n_11080),
.Y(n_11520)
);

AND2x4_ASAP7_75t_L g11521 ( 
.A(n_10922),
.B(n_4588),
.Y(n_11521)
);

INVxp67_ASAP7_75t_L g11522 ( 
.A(n_11198),
.Y(n_11522)
);

BUFx8_ASAP7_75t_L g11523 ( 
.A(n_10849),
.Y(n_11523)
);

INVx1_ASAP7_75t_L g11524 ( 
.A(n_11083),
.Y(n_11524)
);

OAI221xp5_ASAP7_75t_L g11525 ( 
.A1(n_10992),
.A2(n_11008),
.B1(n_10862),
.B2(n_11025),
.C(n_11165),
.Y(n_11525)
);

BUFx8_ASAP7_75t_L g11526 ( 
.A(n_10849),
.Y(n_11526)
);

INVx1_ASAP7_75t_L g11527 ( 
.A(n_11095),
.Y(n_11527)
);

INVx1_ASAP7_75t_L g11528 ( 
.A(n_11098),
.Y(n_11528)
);

OAI22xp5_ASAP7_75t_L g11529 ( 
.A1(n_10779),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_11529)
);

NAND2xp5_ASAP7_75t_L g11530 ( 
.A(n_11035),
.B(n_100),
.Y(n_11530)
);

INVx1_ASAP7_75t_L g11531 ( 
.A(n_11115),
.Y(n_11531)
);

INVx1_ASAP7_75t_L g11532 ( 
.A(n_11121),
.Y(n_11532)
);

INVx1_ASAP7_75t_L g11533 ( 
.A(n_11105),
.Y(n_11533)
);

INVx1_ASAP7_75t_L g11534 ( 
.A(n_11109),
.Y(n_11534)
);

NAND2xp5_ASAP7_75t_L g11535 ( 
.A(n_11047),
.B(n_101),
.Y(n_11535)
);

AND2x2_ASAP7_75t_L g11536 ( 
.A(n_11120),
.B(n_102),
.Y(n_11536)
);

INVx1_ASAP7_75t_L g11537 ( 
.A(n_11112),
.Y(n_11537)
);

INVx1_ASAP7_75t_SL g11538 ( 
.A(n_11100),
.Y(n_11538)
);

AO22x2_ASAP7_75t_L g11539 ( 
.A1(n_11269),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_11539)
);

INVx1_ASAP7_75t_L g11540 ( 
.A(n_11146),
.Y(n_11540)
);

BUFx6f_ASAP7_75t_L g11541 ( 
.A(n_11023),
.Y(n_11541)
);

NAND2x1p5_ASAP7_75t_L g11542 ( 
.A(n_11176),
.B(n_4589),
.Y(n_11542)
);

AND2x4_ASAP7_75t_L g11543 ( 
.A(n_11261),
.B(n_4590),
.Y(n_11543)
);

AO22x2_ASAP7_75t_L g11544 ( 
.A1(n_10842),
.A2(n_106),
.B1(n_103),
.B2(n_104),
.Y(n_11544)
);

INVx1_ASAP7_75t_L g11545 ( 
.A(n_11148),
.Y(n_11545)
);

INVx1_ASAP7_75t_L g11546 ( 
.A(n_11078),
.Y(n_11546)
);

INVx1_ASAP7_75t_L g11547 ( 
.A(n_11084),
.Y(n_11547)
);

INVx2_ASAP7_75t_SL g11548 ( 
.A(n_11114),
.Y(n_11548)
);

INVx2_ASAP7_75t_L g11549 ( 
.A(n_10975),
.Y(n_11549)
);

INVx2_ASAP7_75t_L g11550 ( 
.A(n_10975),
.Y(n_11550)
);

HB1xp67_ASAP7_75t_L g11551 ( 
.A(n_10819),
.Y(n_11551)
);

OAI221xp5_ASAP7_75t_L g11552 ( 
.A1(n_10877),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_11552)
);

NAND2x1p5_ASAP7_75t_L g11553 ( 
.A(n_10804),
.B(n_4591),
.Y(n_11553)
);

NAND2xp5_ASAP7_75t_L g11554 ( 
.A(n_11057),
.B(n_108),
.Y(n_11554)
);

HB1xp67_ASAP7_75t_L g11555 ( 
.A(n_11177),
.Y(n_11555)
);

INVx1_ASAP7_75t_L g11556 ( 
.A(n_11093),
.Y(n_11556)
);

NAND2x1p5_ASAP7_75t_L g11557 ( 
.A(n_10836),
.B(n_4592),
.Y(n_11557)
);

INVx1_ASAP7_75t_L g11558 ( 
.A(n_11094),
.Y(n_11558)
);

CKINVDCx16_ASAP7_75t_R g11559 ( 
.A(n_10935),
.Y(n_11559)
);

CKINVDCx5p33_ASAP7_75t_R g11560 ( 
.A(n_11114),
.Y(n_11560)
);

OAI22xp5_ASAP7_75t_L g11561 ( 
.A1(n_11137),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_11561)
);

NAND2xp5_ASAP7_75t_L g11562 ( 
.A(n_11059),
.B(n_110),
.Y(n_11562)
);

INVx1_ASAP7_75t_L g11563 ( 
.A(n_11097),
.Y(n_11563)
);

OAI22xp5_ASAP7_75t_L g11564 ( 
.A1(n_11207),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_11564)
);

NAND2xp5_ASAP7_75t_L g11565 ( 
.A(n_11062),
.B(n_113),
.Y(n_11565)
);

INVx2_ASAP7_75t_L g11566 ( 
.A(n_10975),
.Y(n_11566)
);

INVx1_ASAP7_75t_L g11567 ( 
.A(n_11102),
.Y(n_11567)
);

OAI221xp5_ASAP7_75t_L g11568 ( 
.A1(n_11183),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.C(n_117),
.Y(n_11568)
);

INVx1_ASAP7_75t_L g11569 ( 
.A(n_11111),
.Y(n_11569)
);

INVx1_ASAP7_75t_L g11570 ( 
.A(n_11113),
.Y(n_11570)
);

NAND2xp5_ASAP7_75t_L g11571 ( 
.A(n_11186),
.B(n_114),
.Y(n_11571)
);

AND2x4_ASAP7_75t_L g11572 ( 
.A(n_10890),
.B(n_4593),
.Y(n_11572)
);

INVx2_ASAP7_75t_SL g11573 ( 
.A(n_10960),
.Y(n_11573)
);

AOI22xp5_ASAP7_75t_L g11574 ( 
.A1(n_11206),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_11574)
);

INVx1_ASAP7_75t_L g11575 ( 
.A(n_11117),
.Y(n_11575)
);

NAND2xp5_ASAP7_75t_L g11576 ( 
.A(n_11192),
.B(n_118),
.Y(n_11576)
);

NAND2x1p5_ASAP7_75t_L g11577 ( 
.A(n_11023),
.B(n_4596),
.Y(n_11577)
);

AND2x4_ASAP7_75t_L g11578 ( 
.A(n_11257),
.B(n_4597),
.Y(n_11578)
);

INVx2_ASAP7_75t_L g11579 ( 
.A(n_10975),
.Y(n_11579)
);

AO22x2_ASAP7_75t_L g11580 ( 
.A1(n_10835),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_11580)
);

INVx1_ASAP7_75t_L g11581 ( 
.A(n_11128),
.Y(n_11581)
);

AND2x2_ASAP7_75t_L g11582 ( 
.A(n_11058),
.B(n_119),
.Y(n_11582)
);

INVx1_ASAP7_75t_L g11583 ( 
.A(n_11129),
.Y(n_11583)
);

OAI221xp5_ASAP7_75t_L g11584 ( 
.A1(n_10927),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_124),
.Y(n_11584)
);

INVx2_ASAP7_75t_L g11585 ( 
.A(n_11020),
.Y(n_11585)
);

NAND2xp5_ASAP7_75t_L g11586 ( 
.A(n_11065),
.B(n_121),
.Y(n_11586)
);

NOR2xp67_ASAP7_75t_L g11587 ( 
.A(n_11205),
.B(n_4599),
.Y(n_11587)
);

BUFx8_ASAP7_75t_L g11588 ( 
.A(n_11043),
.Y(n_11588)
);

INVx1_ASAP7_75t_L g11589 ( 
.A(n_11131),
.Y(n_11589)
);

NAND2xp5_ASAP7_75t_SL g11590 ( 
.A(n_11245),
.B(n_122),
.Y(n_11590)
);

INVx1_ASAP7_75t_L g11591 ( 
.A(n_11135),
.Y(n_11591)
);

INVx1_ASAP7_75t_L g11592 ( 
.A(n_10978),
.Y(n_11592)
);

INVx2_ASAP7_75t_L g11593 ( 
.A(n_11020),
.Y(n_11593)
);

AO22x2_ASAP7_75t_L g11594 ( 
.A1(n_11241),
.A2(n_126),
.B1(n_123),
.B2(n_125),
.Y(n_11594)
);

OAI221xp5_ASAP7_75t_L g11595 ( 
.A1(n_11248),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_11595)
);

INVx2_ASAP7_75t_L g11596 ( 
.A(n_11020),
.Y(n_11596)
);

INVx2_ASAP7_75t_L g11597 ( 
.A(n_11020),
.Y(n_11597)
);

AND2x2_ASAP7_75t_L g11598 ( 
.A(n_11058),
.B(n_10785),
.Y(n_11598)
);

NAND2xp5_ASAP7_75t_L g11599 ( 
.A(n_11071),
.B(n_127),
.Y(n_11599)
);

AND2x6_ASAP7_75t_L g11600 ( 
.A(n_10839),
.B(n_4600),
.Y(n_11600)
);

INVx1_ASAP7_75t_L g11601 ( 
.A(n_10981),
.Y(n_11601)
);

INVx1_ASAP7_75t_L g11602 ( 
.A(n_10987),
.Y(n_11602)
);

INVx1_ASAP7_75t_L g11603 ( 
.A(n_10998),
.Y(n_11603)
);

INVx2_ASAP7_75t_L g11604 ( 
.A(n_11163),
.Y(n_11604)
);

AOI22xp33_ASAP7_75t_L g11605 ( 
.A1(n_11232),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_11605)
);

INVx1_ASAP7_75t_L g11606 ( 
.A(n_11009),
.Y(n_11606)
);

AND2x4_ASAP7_75t_L g11607 ( 
.A(n_11171),
.B(n_4602),
.Y(n_11607)
);

NAND2xp5_ASAP7_75t_L g11608 ( 
.A(n_11073),
.B(n_11136),
.Y(n_11608)
);

AO22x2_ASAP7_75t_L g11609 ( 
.A1(n_10798),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_11609)
);

NAND2xp5_ASAP7_75t_L g11610 ( 
.A(n_11142),
.B(n_132),
.Y(n_11610)
);

AO22x2_ASAP7_75t_L g11611 ( 
.A1(n_11220),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_11611)
);

INVx4_ASAP7_75t_L g11612 ( 
.A(n_11043),
.Y(n_11612)
);

INVx1_ASAP7_75t_L g11613 ( 
.A(n_11014),
.Y(n_11613)
);

INVx6_ASAP7_75t_L g11614 ( 
.A(n_11051),
.Y(n_11614)
);

INVx1_ASAP7_75t_L g11615 ( 
.A(n_11015),
.Y(n_11615)
);

INVx1_ASAP7_75t_L g11616 ( 
.A(n_11017),
.Y(n_11616)
);

AO22x2_ASAP7_75t_L g11617 ( 
.A1(n_10840),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_11617)
);

AO22x2_ASAP7_75t_L g11618 ( 
.A1(n_10794),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_11618)
);

NOR2xp33_ASAP7_75t_L g11619 ( 
.A(n_10821),
.B(n_4603),
.Y(n_11619)
);

INVx1_ASAP7_75t_L g11620 ( 
.A(n_11024),
.Y(n_11620)
);

AO22x2_ASAP7_75t_L g11621 ( 
.A1(n_11193),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_11621)
);

INVx1_ASAP7_75t_L g11622 ( 
.A(n_11029),
.Y(n_11622)
);

INVx2_ASAP7_75t_L g11623 ( 
.A(n_11143),
.Y(n_11623)
);

AOI22xp33_ASAP7_75t_L g11624 ( 
.A1(n_11048),
.A2(n_10953),
.B1(n_10970),
.B2(n_10901),
.Y(n_11624)
);

NOR2xp67_ASAP7_75t_L g11625 ( 
.A(n_11157),
.B(n_11243),
.Y(n_11625)
);

AO22x2_ASAP7_75t_L g11626 ( 
.A1(n_10854),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_11626)
);

AO22x2_ASAP7_75t_L g11627 ( 
.A1(n_11282),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_11627)
);

INVx2_ASAP7_75t_L g11628 ( 
.A(n_11164),
.Y(n_11628)
);

CKINVDCx5p33_ASAP7_75t_R g11629 ( 
.A(n_11285),
.Y(n_11629)
);

OAI21xp33_ASAP7_75t_L g11630 ( 
.A1(n_10988),
.A2(n_141),
.B(n_142),
.Y(n_11630)
);

INVx1_ASAP7_75t_L g11631 ( 
.A(n_11033),
.Y(n_11631)
);

INVx2_ASAP7_75t_L g11632 ( 
.A(n_11166),
.Y(n_11632)
);

A2O1A1Ixp33_ASAP7_75t_L g11633 ( 
.A1(n_10918),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_11633)
);

AO22x2_ASAP7_75t_L g11634 ( 
.A1(n_10872),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_11634)
);

NAND3x1_ASAP7_75t_L g11635 ( 
.A(n_11251),
.B(n_145),
.C(n_146),
.Y(n_11635)
);

INVx1_ASAP7_75t_L g11636 ( 
.A(n_11034),
.Y(n_11636)
);

NAND2xp5_ASAP7_75t_L g11637 ( 
.A(n_11134),
.B(n_146),
.Y(n_11637)
);

NAND2xp5_ASAP7_75t_L g11638 ( 
.A(n_11144),
.B(n_147),
.Y(n_11638)
);

INVx2_ASAP7_75t_L g11639 ( 
.A(n_11153),
.Y(n_11639)
);

OAI22xp5_ASAP7_75t_SL g11640 ( 
.A1(n_11140),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_11640)
);

INVx2_ASAP7_75t_L g11641 ( 
.A(n_11168),
.Y(n_11641)
);

NOR2xp33_ASAP7_75t_L g11642 ( 
.A(n_10858),
.B(n_4604),
.Y(n_11642)
);

NAND2x1p5_ASAP7_75t_L g11643 ( 
.A(n_11051),
.B(n_4605),
.Y(n_11643)
);

AO22x2_ASAP7_75t_L g11644 ( 
.A1(n_11239),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_11644)
);

NOR2xp33_ASAP7_75t_L g11645 ( 
.A(n_10848),
.B(n_4606),
.Y(n_11645)
);

INVx1_ASAP7_75t_L g11646 ( 
.A(n_10928),
.Y(n_11646)
);

AO22x2_ASAP7_75t_L g11647 ( 
.A1(n_11270),
.A2(n_11253),
.B1(n_11271),
.B2(n_11266),
.Y(n_11647)
);

NAND2x1p5_ASAP7_75t_L g11648 ( 
.A(n_11152),
.B(n_11162),
.Y(n_11648)
);

OAI22xp5_ASAP7_75t_L g11649 ( 
.A1(n_11042),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_11649)
);

OR2x2_ASAP7_75t_SL g11650 ( 
.A(n_11229),
.B(n_151),
.Y(n_11650)
);

HB1xp67_ASAP7_75t_L g11651 ( 
.A(n_11249),
.Y(n_11651)
);

OAI22xp5_ASAP7_75t_L g11652 ( 
.A1(n_11101),
.A2(n_11227),
.B1(n_10768),
.B2(n_10792),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_10929),
.Y(n_11653)
);

A2O1A1Ixp33_ASAP7_75t_L g11654 ( 
.A1(n_10864),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_11654)
);

INVx2_ASAP7_75t_L g11655 ( 
.A(n_11170),
.Y(n_11655)
);

NAND2xp5_ASAP7_75t_L g11656 ( 
.A(n_11172),
.B(n_154),
.Y(n_11656)
);

INVx1_ASAP7_75t_SL g11657 ( 
.A(n_11268),
.Y(n_11657)
);

NAND2xp5_ASAP7_75t_L g11658 ( 
.A(n_11187),
.B(n_155),
.Y(n_11658)
);

INVx1_ASAP7_75t_L g11659 ( 
.A(n_10930),
.Y(n_11659)
);

AO22x2_ASAP7_75t_L g11660 ( 
.A1(n_11275),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_11660)
);

INVx1_ASAP7_75t_L g11661 ( 
.A(n_10932),
.Y(n_11661)
);

CKINVDCx5p33_ASAP7_75t_R g11662 ( 
.A(n_11140),
.Y(n_11662)
);

INVx1_ASAP7_75t_L g11663 ( 
.A(n_10934),
.Y(n_11663)
);

AO22x2_ASAP7_75t_L g11664 ( 
.A1(n_11279),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_11664)
);

XOR2x2_ASAP7_75t_L g11665 ( 
.A(n_11278),
.B(n_159),
.Y(n_11665)
);

OR2x6_ASAP7_75t_L g11666 ( 
.A(n_11256),
.B(n_4607),
.Y(n_11666)
);

INVx1_ASAP7_75t_L g11667 ( 
.A(n_10945),
.Y(n_11667)
);

AOI22xp5_ASAP7_75t_L g11668 ( 
.A1(n_11110),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_11668)
);

AND2x6_ASAP7_75t_SL g11669 ( 
.A(n_11123),
.B(n_160),
.Y(n_11669)
);

INVx1_ASAP7_75t_L g11670 ( 
.A(n_10860),
.Y(n_11670)
);

NAND2xp5_ASAP7_75t_L g11671 ( 
.A(n_11222),
.B(n_162),
.Y(n_11671)
);

NAND2xp5_ASAP7_75t_L g11672 ( 
.A(n_11221),
.B(n_163),
.Y(n_11672)
);

AND2x2_ASAP7_75t_L g11673 ( 
.A(n_10982),
.B(n_164),
.Y(n_11673)
);

AO22x2_ASAP7_75t_L g11674 ( 
.A1(n_11200),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_11674)
);

INVx2_ASAP7_75t_L g11675 ( 
.A(n_11173),
.Y(n_11675)
);

AOI22xp5_ASAP7_75t_L g11676 ( 
.A1(n_11139),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_11676)
);

NAND2xp5_ASAP7_75t_L g11677 ( 
.A(n_11223),
.B(n_11235),
.Y(n_11677)
);

INVxp67_ASAP7_75t_L g11678 ( 
.A(n_11260),
.Y(n_11678)
);

INVx1_ASAP7_75t_L g11679 ( 
.A(n_10861),
.Y(n_11679)
);

NAND2xp5_ASAP7_75t_L g11680 ( 
.A(n_10868),
.B(n_167),
.Y(n_11680)
);

AND2x2_ASAP7_75t_L g11681 ( 
.A(n_11175),
.B(n_168),
.Y(n_11681)
);

INVx2_ASAP7_75t_L g11682 ( 
.A(n_11185),
.Y(n_11682)
);

NAND2x1p5_ASAP7_75t_L g11683 ( 
.A(n_11152),
.B(n_4608),
.Y(n_11683)
);

OAI221xp5_ASAP7_75t_L g11684 ( 
.A1(n_11092),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_11684)
);

NOR2xp33_ASAP7_75t_L g11685 ( 
.A(n_10852),
.B(n_4609),
.Y(n_11685)
);

INVx1_ASAP7_75t_L g11686 ( 
.A(n_10874),
.Y(n_11686)
);

NAND2xp5_ASAP7_75t_L g11687 ( 
.A(n_10879),
.B(n_10881),
.Y(n_11687)
);

AND2x4_ASAP7_75t_L g11688 ( 
.A(n_11258),
.B(n_4610),
.Y(n_11688)
);

HB1xp67_ASAP7_75t_L g11689 ( 
.A(n_10937),
.Y(n_11689)
);

INVx1_ASAP7_75t_L g11690 ( 
.A(n_10886),
.Y(n_11690)
);

INVx1_ASAP7_75t_L g11691 ( 
.A(n_10887),
.Y(n_11691)
);

BUFx3_ASAP7_75t_L g11692 ( 
.A(n_11162),
.Y(n_11692)
);

AOI22xp33_ASAP7_75t_L g11693 ( 
.A1(n_11159),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_11693)
);

INVx1_ASAP7_75t_L g11694 ( 
.A(n_10892),
.Y(n_11694)
);

NAND2xp5_ASAP7_75t_L g11695 ( 
.A(n_10898),
.B(n_172),
.Y(n_11695)
);

AO22x2_ASAP7_75t_L g11696 ( 
.A1(n_11195),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_11696)
);

BUFx8_ASAP7_75t_L g11697 ( 
.A(n_10966),
.Y(n_11697)
);

BUFx2_ASAP7_75t_L g11698 ( 
.A(n_11019),
.Y(n_11698)
);

BUFx6f_ASAP7_75t_L g11699 ( 
.A(n_11072),
.Y(n_11699)
);

AO22x2_ASAP7_75t_L g11700 ( 
.A1(n_11001),
.A2(n_177),
.B1(n_173),
.B2(n_176),
.Y(n_11700)
);

INVx1_ASAP7_75t_L g11701 ( 
.A(n_10905),
.Y(n_11701)
);

AO22x2_ASAP7_75t_L g11702 ( 
.A1(n_11230),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_11702)
);

NAND2xp5_ASAP7_75t_L g11703 ( 
.A(n_10921),
.B(n_179),
.Y(n_11703)
);

INVx1_ASAP7_75t_L g11704 ( 
.A(n_10972),
.Y(n_11704)
);

AO22x2_ASAP7_75t_L g11705 ( 
.A1(n_11231),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_11705)
);

INVxp67_ASAP7_75t_L g11706 ( 
.A(n_11264),
.Y(n_11706)
);

NAND2x1p5_ASAP7_75t_L g11707 ( 
.A(n_11037),
.B(n_4611),
.Y(n_11707)
);

INVx1_ASAP7_75t_L g11708 ( 
.A(n_10974),
.Y(n_11708)
);

AO22x2_ASAP7_75t_L g11709 ( 
.A1(n_11234),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_11709)
);

CKINVDCx20_ASAP7_75t_R g11710 ( 
.A(n_11119),
.Y(n_11710)
);

INVxp67_ASAP7_75t_L g11711 ( 
.A(n_11267),
.Y(n_11711)
);

INVx1_ASAP7_75t_L g11712 ( 
.A(n_10841),
.Y(n_11712)
);

INVx1_ASAP7_75t_L g11713 ( 
.A(n_11018),
.Y(n_11713)
);

AOI22xp33_ASAP7_75t_L g11714 ( 
.A1(n_11201),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_11714)
);

NOR2xp33_ASAP7_75t_L g11715 ( 
.A(n_11224),
.B(n_4614),
.Y(n_11715)
);

INVx1_ASAP7_75t_L g11716 ( 
.A(n_11178),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_11246),
.B(n_184),
.Y(n_11717)
);

INVx1_ASAP7_75t_L g11718 ( 
.A(n_10897),
.Y(n_11718)
);

AO22x2_ASAP7_75t_L g11719 ( 
.A1(n_11155),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_11719)
);

OAI221xp5_ASAP7_75t_L g11720 ( 
.A1(n_11108),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_11720)
);

AO22x2_ASAP7_75t_L g11721 ( 
.A1(n_11182),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_11721)
);

AOI22xp5_ASAP7_75t_L g11722 ( 
.A1(n_11214),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_11722)
);

INVx1_ASAP7_75t_L g11723 ( 
.A(n_10897),
.Y(n_11723)
);

BUFx6f_ASAP7_75t_SL g11724 ( 
.A(n_10870),
.Y(n_11724)
);

INVxp67_ASAP7_75t_L g11725 ( 
.A(n_10910),
.Y(n_11725)
);

INVx1_ASAP7_75t_L g11726 ( 
.A(n_10897),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_11204),
.Y(n_11727)
);

NAND2x1p5_ASAP7_75t_L g11728 ( 
.A(n_11150),
.B(n_4615),
.Y(n_11728)
);

AO22x2_ASAP7_75t_L g11729 ( 
.A1(n_11184),
.A2(n_11197),
.B1(n_11089),
.B2(n_11104),
.Y(n_11729)
);

AND2x4_ASAP7_75t_L g11730 ( 
.A(n_11118),
.B(n_4616),
.Y(n_11730)
);

AO22x2_ASAP7_75t_L g11731 ( 
.A1(n_11081),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_11731)
);

INVx1_ASAP7_75t_L g11732 ( 
.A(n_11216),
.Y(n_11732)
);

INVx2_ASAP7_75t_L g11733 ( 
.A(n_11247),
.Y(n_11733)
);

CKINVDCx14_ASAP7_75t_R g11734 ( 
.A(n_11123),
.Y(n_11734)
);

INVxp67_ASAP7_75t_SL g11735 ( 
.A(n_11049),
.Y(n_11735)
);

OAI221xp5_ASAP7_75t_L g11736 ( 
.A1(n_11188),
.A2(n_195),
.B1(n_192),
.B2(n_194),
.C(n_196),
.Y(n_11736)
);

CKINVDCx5p33_ASAP7_75t_R g11737 ( 
.A(n_11145),
.Y(n_11737)
);

INVx1_ASAP7_75t_L g11738 ( 
.A(n_11056),
.Y(n_11738)
);

NAND2x1p5_ASAP7_75t_L g11739 ( 
.A(n_11151),
.B(n_4617),
.Y(n_11739)
);

BUFx8_ASAP7_75t_L g11740 ( 
.A(n_11161),
.Y(n_11740)
);

INVxp67_ASAP7_75t_L g11741 ( 
.A(n_11169),
.Y(n_11741)
);

INVx2_ASAP7_75t_L g11742 ( 
.A(n_11085),
.Y(n_11742)
);

NAND2xp5_ASAP7_75t_L g11743 ( 
.A(n_10826),
.B(n_11016),
.Y(n_11743)
);

INVx1_ASAP7_75t_L g11744 ( 
.A(n_11130),
.Y(n_11744)
);

NAND2xp5_ASAP7_75t_L g11745 ( 
.A(n_11106),
.B(n_196),
.Y(n_11745)
);

OR2x6_ASAP7_75t_L g11746 ( 
.A(n_11252),
.B(n_4618),
.Y(n_11746)
);

INVx2_ASAP7_75t_SL g11747 ( 
.A(n_10847),
.Y(n_11747)
);

AO22x2_ASAP7_75t_L g11748 ( 
.A1(n_10948),
.A2(n_10952),
.B1(n_11052),
.B2(n_11005),
.Y(n_11748)
);

NOR2xp33_ASAP7_75t_L g11749 ( 
.A(n_10875),
.B(n_4619),
.Y(n_11749)
);

INVx1_ASAP7_75t_L g11750 ( 
.A(n_11238),
.Y(n_11750)
);

INVx1_ASAP7_75t_L g11751 ( 
.A(n_11244),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_10939),
.Y(n_11752)
);

INVx1_ASAP7_75t_L g11753 ( 
.A(n_11087),
.Y(n_11753)
);

HB1xp67_ASAP7_75t_L g11754 ( 
.A(n_11069),
.Y(n_11754)
);

INVxp67_ASAP7_75t_L g11755 ( 
.A(n_10976),
.Y(n_11755)
);

INVx2_ASAP7_75t_L g11756 ( 
.A(n_11116),
.Y(n_11756)
);

AO22x2_ASAP7_75t_L g11757 ( 
.A1(n_11075),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_11757)
);

NAND2xp5_ASAP7_75t_SL g11758 ( 
.A(n_11007),
.B(n_197),
.Y(n_11758)
);

BUFx2_ASAP7_75t_L g11759 ( 
.A(n_10963),
.Y(n_11759)
);

INVx1_ASAP7_75t_L g11760 ( 
.A(n_11133),
.Y(n_11760)
);

INVxp67_ASAP7_75t_L g11761 ( 
.A(n_11199),
.Y(n_11761)
);

AO22x2_ASAP7_75t_L g11762 ( 
.A1(n_11125),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_11762)
);

AND2x4_ASAP7_75t_L g11763 ( 
.A(n_11126),
.B(n_4621),
.Y(n_11763)
);

INVx1_ASAP7_75t_L g11764 ( 
.A(n_10884),
.Y(n_11764)
);

CKINVDCx5p33_ASAP7_75t_R g11765 ( 
.A(n_11103),
.Y(n_11765)
);

INVx1_ASAP7_75t_L g11766 ( 
.A(n_11124),
.Y(n_11766)
);

XNOR2xp5_ASAP7_75t_L g11767 ( 
.A(n_11030),
.B(n_4622),
.Y(n_11767)
);

AOI22xp5_ASAP7_75t_L g11768 ( 
.A1(n_11003),
.A2(n_11079),
.B1(n_10906),
.B2(n_10914),
.Y(n_11768)
);

INVx1_ASAP7_75t_L g11769 ( 
.A(n_11191),
.Y(n_11769)
);

INVx1_ASAP7_75t_L g11770 ( 
.A(n_11028),
.Y(n_11770)
);

OAI221xp5_ASAP7_75t_L g11771 ( 
.A1(n_11254),
.A2(n_203),
.B1(n_200),
.B2(n_202),
.C(n_204),
.Y(n_11771)
);

NAND2x1p5_ASAP7_75t_L g11772 ( 
.A(n_10907),
.B(n_4625),
.Y(n_11772)
);

AO22x2_ASAP7_75t_L g11773 ( 
.A1(n_10904),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_11773)
);

INVx1_ASAP7_75t_L g11774 ( 
.A(n_10951),
.Y(n_11774)
);

INVx1_ASAP7_75t_L g11775 ( 
.A(n_10917),
.Y(n_11775)
);

NAND2xp5_ASAP7_75t_L g11776 ( 
.A(n_11091),
.B(n_205),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_10924),
.Y(n_11777)
);

AND2x4_ASAP7_75t_L g11778 ( 
.A(n_11250),
.B(n_4627),
.Y(n_11778)
);

CKINVDCx5p33_ASAP7_75t_R g11779 ( 
.A(n_11060),
.Y(n_11779)
);

INVx1_ASAP7_75t_L g11780 ( 
.A(n_11021),
.Y(n_11780)
);

OAI221xp5_ASAP7_75t_L g11781 ( 
.A1(n_11032),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.C(n_208),
.Y(n_11781)
);

INVx1_ASAP7_75t_L g11782 ( 
.A(n_10926),
.Y(n_11782)
);

NAND2xp5_ASAP7_75t_L g11783 ( 
.A(n_11032),
.B(n_207),
.Y(n_11783)
);

NAND2x1p5_ASAP7_75t_L g11784 ( 
.A(n_10856),
.B(n_4628),
.Y(n_11784)
);

AO22x2_ASAP7_75t_L g11785 ( 
.A1(n_10801),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_11785)
);

NAND2x1p5_ASAP7_75t_L g11786 ( 
.A(n_10856),
.B(n_4629),
.Y(n_11786)
);

OAI221xp5_ASAP7_75t_L g11787 ( 
.A1(n_11032),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.C(n_212),
.Y(n_11787)
);

AO22x2_ASAP7_75t_L g11788 ( 
.A1(n_10801),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_11788)
);

NOR2xp33_ASAP7_75t_L g11789 ( 
.A(n_11032),
.B(n_4630),
.Y(n_11789)
);

AO22x2_ASAP7_75t_L g11790 ( 
.A1(n_10801),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_11790)
);

INVx1_ASAP7_75t_L g11791 ( 
.A(n_10926),
.Y(n_11791)
);

INVx1_ASAP7_75t_L g11792 ( 
.A(n_10926),
.Y(n_11792)
);

INVx1_ASAP7_75t_L g11793 ( 
.A(n_10926),
.Y(n_11793)
);

INVx1_ASAP7_75t_L g11794 ( 
.A(n_10926),
.Y(n_11794)
);

INVx1_ASAP7_75t_L g11795 ( 
.A(n_10926),
.Y(n_11795)
);

INVx1_ASAP7_75t_L g11796 ( 
.A(n_10926),
.Y(n_11796)
);

NAND2x1p5_ASAP7_75t_L g11797 ( 
.A(n_10856),
.B(n_4632),
.Y(n_11797)
);

AND2x4_ASAP7_75t_L g11798 ( 
.A(n_10808),
.B(n_4633),
.Y(n_11798)
);

NAND2xp5_ASAP7_75t_L g11799 ( 
.A(n_11032),
.B(n_215),
.Y(n_11799)
);

INVx2_ASAP7_75t_L g11800 ( 
.A(n_10789),
.Y(n_11800)
);

BUFx8_ASAP7_75t_L g11801 ( 
.A(n_11027),
.Y(n_11801)
);

BUFx8_ASAP7_75t_L g11802 ( 
.A(n_11027),
.Y(n_11802)
);

INVx1_ASAP7_75t_L g11803 ( 
.A(n_10926),
.Y(n_11803)
);

INVx1_ASAP7_75t_L g11804 ( 
.A(n_10926),
.Y(n_11804)
);

INVx1_ASAP7_75t_L g11805 ( 
.A(n_10926),
.Y(n_11805)
);

INVx2_ASAP7_75t_L g11806 ( 
.A(n_10789),
.Y(n_11806)
);

AND2x4_ASAP7_75t_L g11807 ( 
.A(n_10808),
.B(n_4634),
.Y(n_11807)
);

INVx1_ASAP7_75t_L g11808 ( 
.A(n_10926),
.Y(n_11808)
);

INVx1_ASAP7_75t_L g11809 ( 
.A(n_10926),
.Y(n_11809)
);

AND2x2_ASAP7_75t_L g11810 ( 
.A(n_10812),
.B(n_216),
.Y(n_11810)
);

NAND2xp5_ASAP7_75t_L g11811 ( 
.A(n_11032),
.B(n_216),
.Y(n_11811)
);

AND2x4_ASAP7_75t_L g11812 ( 
.A(n_10808),
.B(n_4635),
.Y(n_11812)
);

INVx1_ASAP7_75t_L g11813 ( 
.A(n_10926),
.Y(n_11813)
);

AO22x2_ASAP7_75t_L g11814 ( 
.A1(n_10801),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_11814)
);

INVx1_ASAP7_75t_L g11815 ( 
.A(n_10926),
.Y(n_11815)
);

NAND2xp5_ASAP7_75t_L g11816 ( 
.A(n_11032),
.B(n_217),
.Y(n_11816)
);

INVx2_ASAP7_75t_L g11817 ( 
.A(n_10789),
.Y(n_11817)
);

INVx1_ASAP7_75t_L g11818 ( 
.A(n_10926),
.Y(n_11818)
);

INVx1_ASAP7_75t_L g11819 ( 
.A(n_10926),
.Y(n_11819)
);

INVx2_ASAP7_75t_L g11820 ( 
.A(n_10789),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_10926),
.Y(n_11821)
);

BUFx6f_ASAP7_75t_SL g11822 ( 
.A(n_10771),
.Y(n_11822)
);

INVx1_ASAP7_75t_L g11823 ( 
.A(n_10926),
.Y(n_11823)
);

INVx1_ASAP7_75t_L g11824 ( 
.A(n_10926),
.Y(n_11824)
);

AOI22xp33_ASAP7_75t_L g11825 ( 
.A1(n_11032),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_11825)
);

INVx1_ASAP7_75t_L g11826 ( 
.A(n_10926),
.Y(n_11826)
);

AO22x2_ASAP7_75t_L g11827 ( 
.A1(n_10801),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_11827)
);

INVx1_ASAP7_75t_L g11828 ( 
.A(n_10926),
.Y(n_11828)
);

INVx2_ASAP7_75t_L g11829 ( 
.A(n_10789),
.Y(n_11829)
);

INVx1_ASAP7_75t_L g11830 ( 
.A(n_10926),
.Y(n_11830)
);

NAND2x1p5_ASAP7_75t_L g11831 ( 
.A(n_10856),
.B(n_4636),
.Y(n_11831)
);

AOI22xp5_ASAP7_75t_SL g11832 ( 
.A1(n_11032),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_11832)
);

AO22x2_ASAP7_75t_L g11833 ( 
.A1(n_10801),
.A2(n_226),
.B1(n_223),
.B2(n_225),
.Y(n_11833)
);

AO22x2_ASAP7_75t_L g11834 ( 
.A1(n_10801),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_11834)
);

NAND2xp5_ASAP7_75t_L g11835 ( 
.A(n_11032),
.B(n_227),
.Y(n_11835)
);

NOR2xp67_ASAP7_75t_L g11836 ( 
.A(n_11189),
.B(n_4637),
.Y(n_11836)
);

INVx3_ASAP7_75t_L g11837 ( 
.A(n_10960),
.Y(n_11837)
);

HB1xp67_ASAP7_75t_L g11838 ( 
.A(n_10776),
.Y(n_11838)
);

INVx1_ASAP7_75t_L g11839 ( 
.A(n_10926),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_10926),
.Y(n_11840)
);

INVx2_ASAP7_75t_L g11841 ( 
.A(n_10789),
.Y(n_11841)
);

NAND2xp5_ASAP7_75t_SL g11842 ( 
.A(n_11032),
.B(n_228),
.Y(n_11842)
);

INVx1_ASAP7_75t_L g11843 ( 
.A(n_10926),
.Y(n_11843)
);

NAND2xp5_ASAP7_75t_L g11844 ( 
.A(n_11032),
.B(n_229),
.Y(n_11844)
);

INVx1_ASAP7_75t_L g11845 ( 
.A(n_10926),
.Y(n_11845)
);

AND2x2_ASAP7_75t_L g11846 ( 
.A(n_10812),
.B(n_230),
.Y(n_11846)
);

INVx2_ASAP7_75t_L g11847 ( 
.A(n_10789),
.Y(n_11847)
);

AOI22xp5_ASAP7_75t_L g11848 ( 
.A1(n_11032),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_11848)
);

NAND2xp5_ASAP7_75t_L g11849 ( 
.A(n_11032),
.B(n_231),
.Y(n_11849)
);

INVx1_ASAP7_75t_L g11850 ( 
.A(n_10926),
.Y(n_11850)
);

INVx1_ASAP7_75t_L g11851 ( 
.A(n_10926),
.Y(n_11851)
);

AOI22xp5_ASAP7_75t_L g11852 ( 
.A1(n_11032),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_11852)
);

INVx1_ASAP7_75t_L g11853 ( 
.A(n_10926),
.Y(n_11853)
);

AND2x2_ASAP7_75t_L g11854 ( 
.A(n_10812),
.B(n_233),
.Y(n_11854)
);

INVx1_ASAP7_75t_L g11855 ( 
.A(n_10926),
.Y(n_11855)
);

AND2x2_ASAP7_75t_L g11856 ( 
.A(n_10812),
.B(n_234),
.Y(n_11856)
);

INVx1_ASAP7_75t_L g11857 ( 
.A(n_10926),
.Y(n_11857)
);

INVx1_ASAP7_75t_L g11858 ( 
.A(n_10926),
.Y(n_11858)
);

NAND2x1p5_ASAP7_75t_L g11859 ( 
.A(n_10856),
.B(n_4638),
.Y(n_11859)
);

AND2x2_ASAP7_75t_L g11860 ( 
.A(n_10812),
.B(n_235),
.Y(n_11860)
);

NAND2xp5_ASAP7_75t_L g11861 ( 
.A(n_11032),
.B(n_236),
.Y(n_11861)
);

INVx1_ASAP7_75t_L g11862 ( 
.A(n_10926),
.Y(n_11862)
);

INVx1_ASAP7_75t_L g11863 ( 
.A(n_10926),
.Y(n_11863)
);

AND2x4_ASAP7_75t_L g11864 ( 
.A(n_10808),
.B(n_4640),
.Y(n_11864)
);

INVx2_ASAP7_75t_L g11865 ( 
.A(n_10789),
.Y(n_11865)
);

AO22x2_ASAP7_75t_L g11866 ( 
.A1(n_10801),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_11866)
);

INVx1_ASAP7_75t_L g11867 ( 
.A(n_10926),
.Y(n_11867)
);

INVx1_ASAP7_75t_L g11868 ( 
.A(n_10926),
.Y(n_11868)
);

BUFx3_ASAP7_75t_L g11869 ( 
.A(n_11122),
.Y(n_11869)
);

NAND3xp33_ASAP7_75t_L g11870 ( 
.A(n_11032),
.B(n_237),
.C(n_238),
.Y(n_11870)
);

AO22x2_ASAP7_75t_L g11871 ( 
.A1(n_10801),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_11871)
);

NAND2xp5_ASAP7_75t_L g11872 ( 
.A(n_11032),
.B(n_240),
.Y(n_11872)
);

OAI221xp5_ASAP7_75t_L g11873 ( 
.A1(n_11032),
.A2(n_244),
.B1(n_241),
.B2(n_242),
.C(n_245),
.Y(n_11873)
);

INVx1_ASAP7_75t_L g11874 ( 
.A(n_10926),
.Y(n_11874)
);

INVx1_ASAP7_75t_L g11875 ( 
.A(n_10926),
.Y(n_11875)
);

INVx1_ASAP7_75t_L g11876 ( 
.A(n_10926),
.Y(n_11876)
);

INVx2_ASAP7_75t_L g11877 ( 
.A(n_10789),
.Y(n_11877)
);

AOI22xp5_ASAP7_75t_L g11878 ( 
.A1(n_11032),
.A2(n_246),
.B1(n_242),
.B2(n_245),
.Y(n_11878)
);

AND2x2_ASAP7_75t_L g11879 ( 
.A(n_10812),
.B(n_246),
.Y(n_11879)
);

NAND2xp5_ASAP7_75t_SL g11880 ( 
.A(n_11032),
.B(n_247),
.Y(n_11880)
);

AND2x2_ASAP7_75t_L g11881 ( 
.A(n_10812),
.B(n_247),
.Y(n_11881)
);

NOR2xp33_ASAP7_75t_L g11882 ( 
.A(n_11032),
.B(n_4641),
.Y(n_11882)
);

INVx1_ASAP7_75t_L g11883 ( 
.A(n_10926),
.Y(n_11883)
);

NAND2xp5_ASAP7_75t_L g11884 ( 
.A(n_11032),
.B(n_248),
.Y(n_11884)
);

INVx2_ASAP7_75t_L g11885 ( 
.A(n_10789),
.Y(n_11885)
);

INVx1_ASAP7_75t_L g11886 ( 
.A(n_10926),
.Y(n_11886)
);

AO22x2_ASAP7_75t_L g11887 ( 
.A1(n_10801),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_11887)
);

AO22x2_ASAP7_75t_L g11888 ( 
.A1(n_10801),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_11888)
);

INVx1_ASAP7_75t_L g11889 ( 
.A(n_10926),
.Y(n_11889)
);

OR2x2_ASAP7_75t_L g11890 ( 
.A(n_10776),
.B(n_252),
.Y(n_11890)
);

BUFx3_ASAP7_75t_L g11891 ( 
.A(n_11122),
.Y(n_11891)
);

INVx2_ASAP7_75t_L g11892 ( 
.A(n_10789),
.Y(n_11892)
);

BUFx2_ASAP7_75t_SL g11893 ( 
.A(n_10856),
.Y(n_11893)
);

INVx1_ASAP7_75t_L g11894 ( 
.A(n_10926),
.Y(n_11894)
);

INVx1_ASAP7_75t_L g11895 ( 
.A(n_10926),
.Y(n_11895)
);

AND2x4_ASAP7_75t_L g11896 ( 
.A(n_10808),
.B(n_4642),
.Y(n_11896)
);

AND2x6_ASAP7_75t_L g11897 ( 
.A(n_11158),
.B(n_4643),
.Y(n_11897)
);

INVx1_ASAP7_75t_L g11898 ( 
.A(n_10926),
.Y(n_11898)
);

INVx1_ASAP7_75t_L g11899 ( 
.A(n_10926),
.Y(n_11899)
);

AND2x6_ASAP7_75t_L g11900 ( 
.A(n_11158),
.B(n_4644),
.Y(n_11900)
);

INVx1_ASAP7_75t_L g11901 ( 
.A(n_10926),
.Y(n_11901)
);

AO22x2_ASAP7_75t_L g11902 ( 
.A1(n_10801),
.A2(n_255),
.B1(n_252),
.B2(n_254),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_10926),
.Y(n_11903)
);

AND2x2_ASAP7_75t_L g11904 ( 
.A(n_10812),
.B(n_254),
.Y(n_11904)
);

AO22x2_ASAP7_75t_L g11905 ( 
.A1(n_10801),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_11905)
);

AOI22xp5_ASAP7_75t_L g11906 ( 
.A1(n_11032),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_11906)
);

INVx1_ASAP7_75t_SL g11907 ( 
.A(n_10817),
.Y(n_11907)
);

CKINVDCx20_ASAP7_75t_R g11908 ( 
.A(n_10828),
.Y(n_11908)
);

AO22x2_ASAP7_75t_L g11909 ( 
.A1(n_10801),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_11909)
);

INVx1_ASAP7_75t_L g11910 ( 
.A(n_10926),
.Y(n_11910)
);

OAI221xp5_ASAP7_75t_L g11911 ( 
.A1(n_11032),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.C(n_262),
.Y(n_11911)
);

INVx2_ASAP7_75t_SL g11912 ( 
.A(n_10999),
.Y(n_11912)
);

INVx1_ASAP7_75t_L g11913 ( 
.A(n_10926),
.Y(n_11913)
);

NAND2x1p5_ASAP7_75t_L g11914 ( 
.A(n_10856),
.B(n_4645),
.Y(n_11914)
);

INVxp67_ASAP7_75t_L g11915 ( 
.A(n_10787),
.Y(n_11915)
);

NAND2x1p5_ASAP7_75t_L g11916 ( 
.A(n_10856),
.B(n_4647),
.Y(n_11916)
);

OAI22xp33_ASAP7_75t_SL g11917 ( 
.A1(n_11032),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_11917)
);

INVx1_ASAP7_75t_L g11918 ( 
.A(n_10926),
.Y(n_11918)
);

AND2x6_ASAP7_75t_L g11919 ( 
.A(n_11158),
.B(n_4649),
.Y(n_11919)
);

NAND2xp33_ASAP7_75t_L g11920 ( 
.A(n_10801),
.B(n_263),
.Y(n_11920)
);

NAND2xp33_ASAP7_75t_L g11921 ( 
.A(n_10801),
.B(n_265),
.Y(n_11921)
);

NAND2xp5_ASAP7_75t_L g11922 ( 
.A(n_11032),
.B(n_266),
.Y(n_11922)
);

INVxp67_ASAP7_75t_L g11923 ( 
.A(n_10787),
.Y(n_11923)
);

OAI22xp5_ASAP7_75t_L g11924 ( 
.A1(n_11032),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_11924)
);

INVx1_ASAP7_75t_L g11925 ( 
.A(n_10926),
.Y(n_11925)
);

AND2x2_ASAP7_75t_L g11926 ( 
.A(n_10812),
.B(n_267),
.Y(n_11926)
);

INVx1_ASAP7_75t_L g11927 ( 
.A(n_10926),
.Y(n_11927)
);

INVx2_ASAP7_75t_L g11928 ( 
.A(n_10789),
.Y(n_11928)
);

INVx1_ASAP7_75t_L g11929 ( 
.A(n_10926),
.Y(n_11929)
);

A2O1A1Ixp33_ASAP7_75t_L g11930 ( 
.A1(n_11293),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_11930)
);

INVx1_ASAP7_75t_L g11931 ( 
.A(n_11355),
.Y(n_11931)
);

NOR2xp33_ASAP7_75t_L g11932 ( 
.A(n_11288),
.B(n_4650),
.Y(n_11932)
);

INVx1_ASAP7_75t_L g11933 ( 
.A(n_11356),
.Y(n_11933)
);

AOI21xp5_ASAP7_75t_L g11934 ( 
.A1(n_11432),
.A2(n_4654),
.B(n_4651),
.Y(n_11934)
);

NAND2xp5_ASAP7_75t_SL g11935 ( 
.A(n_11391),
.B(n_4655),
.Y(n_11935)
);

AOI21xp5_ASAP7_75t_L g11936 ( 
.A1(n_11338),
.A2(n_4657),
.B(n_4656),
.Y(n_11936)
);

AOI21xp5_ASAP7_75t_L g11937 ( 
.A1(n_11920),
.A2(n_11921),
.B(n_11417),
.Y(n_11937)
);

NAND2xp5_ASAP7_75t_L g11938 ( 
.A(n_11346),
.B(n_11838),
.Y(n_11938)
);

INVx3_ASAP7_75t_L g11939 ( 
.A(n_11316),
.Y(n_11939)
);

CKINVDCx5p33_ASAP7_75t_R g11940 ( 
.A(n_11342),
.Y(n_11940)
);

AO32x2_ASAP7_75t_L g11941 ( 
.A1(n_11529),
.A2(n_271),
.A3(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_11941)
);

AOI22xp33_ASAP7_75t_L g11942 ( 
.A1(n_11416),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_11942)
);

BUFx6f_ASAP7_75t_L g11943 ( 
.A(n_11541),
.Y(n_11943)
);

AOI21xp5_ASAP7_75t_L g11944 ( 
.A1(n_11624),
.A2(n_4660),
.B(n_4659),
.Y(n_11944)
);

AOI21xp5_ASAP7_75t_L g11945 ( 
.A1(n_11608),
.A2(n_4664),
.B(n_4662),
.Y(n_11945)
);

OAI21xp5_ASAP7_75t_L g11946 ( 
.A1(n_11294),
.A2(n_273),
.B(n_274),
.Y(n_11946)
);

AOI21xp5_ASAP7_75t_L g11947 ( 
.A1(n_11687),
.A2(n_4666),
.B(n_4665),
.Y(n_11947)
);

AOI21xp5_ASAP7_75t_L g11948 ( 
.A1(n_11789),
.A2(n_4668),
.B(n_4667),
.Y(n_11948)
);

O2A1O1Ixp5_ASAP7_75t_L g11949 ( 
.A1(n_11654),
.A2(n_11880),
.B(n_11842),
.C(n_11882),
.Y(n_11949)
);

AO22x1_ASAP7_75t_L g11950 ( 
.A1(n_11897),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_11950)
);

NAND2xp5_ASAP7_75t_L g11951 ( 
.A(n_11670),
.B(n_275),
.Y(n_11951)
);

AOI21xp5_ASAP7_75t_L g11952 ( 
.A1(n_11339),
.A2(n_11525),
.B(n_11337),
.Y(n_11952)
);

NAND2xp5_ASAP7_75t_L g11953 ( 
.A(n_11679),
.B(n_11686),
.Y(n_11953)
);

NAND2xp5_ASAP7_75t_L g11954 ( 
.A(n_11690),
.B(n_276),
.Y(n_11954)
);

A2O1A1Ixp33_ASAP7_75t_L g11955 ( 
.A1(n_11420),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_11955)
);

OAI21xp33_ASAP7_75t_L g11956 ( 
.A1(n_11303),
.A2(n_278),
.B(n_279),
.Y(n_11956)
);

A2O1A1Ixp33_ASAP7_75t_L g11957 ( 
.A1(n_11625),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_11957)
);

CKINVDCx10_ASAP7_75t_R g11958 ( 
.A(n_11822),
.Y(n_11958)
);

AOI21x1_ASAP7_75t_L g11959 ( 
.A1(n_11647),
.A2(n_4675),
.B(n_4669),
.Y(n_11959)
);

AND2x4_ASAP7_75t_L g11960 ( 
.A(n_11407),
.B(n_4676),
.Y(n_11960)
);

NAND2xp5_ASAP7_75t_L g11961 ( 
.A(n_11691),
.B(n_280),
.Y(n_11961)
);

AOI21xp5_ASAP7_75t_L g11962 ( 
.A1(n_11287),
.A2(n_4679),
.B(n_4678),
.Y(n_11962)
);

AOI21xp5_ASAP7_75t_L g11963 ( 
.A1(n_11290),
.A2(n_4682),
.B(n_4681),
.Y(n_11963)
);

INVx2_ASAP7_75t_L g11964 ( 
.A(n_11311),
.Y(n_11964)
);

AOI21xp5_ASAP7_75t_L g11965 ( 
.A1(n_11782),
.A2(n_4684),
.B(n_4683),
.Y(n_11965)
);

BUFx6f_ASAP7_75t_L g11966 ( 
.A(n_11541),
.Y(n_11966)
);

NAND2xp5_ASAP7_75t_L g11967 ( 
.A(n_11694),
.B(n_11701),
.Y(n_11967)
);

BUFx6f_ASAP7_75t_L g11968 ( 
.A(n_11692),
.Y(n_11968)
);

INVx2_ASAP7_75t_L g11969 ( 
.A(n_11330),
.Y(n_11969)
);

OR2x6_ASAP7_75t_L g11970 ( 
.A(n_11893),
.B(n_4686),
.Y(n_11970)
);

AOI21xp5_ASAP7_75t_L g11971 ( 
.A1(n_11791),
.A2(n_4688),
.B(n_4687),
.Y(n_11971)
);

NAND2x1_ASAP7_75t_L g11972 ( 
.A(n_11752),
.B(n_4689),
.Y(n_11972)
);

NOR2xp33_ASAP7_75t_R g11973 ( 
.A(n_11908),
.B(n_4690),
.Y(n_11973)
);

AOI21xp5_ASAP7_75t_L g11974 ( 
.A1(n_11792),
.A2(n_4692),
.B(n_4691),
.Y(n_11974)
);

NOR2x1_ASAP7_75t_L g11975 ( 
.A(n_11870),
.B(n_282),
.Y(n_11975)
);

NOR2xp33_ASAP7_75t_SL g11976 ( 
.A(n_11361),
.B(n_4693),
.Y(n_11976)
);

NAND2xp5_ASAP7_75t_SL g11977 ( 
.A(n_11646),
.B(n_4694),
.Y(n_11977)
);

NAND2xp5_ASAP7_75t_L g11978 ( 
.A(n_11704),
.B(n_283),
.Y(n_11978)
);

AOI21xp5_ASAP7_75t_L g11979 ( 
.A1(n_11793),
.A2(n_4696),
.B(n_4695),
.Y(n_11979)
);

AOI21xp5_ASAP7_75t_L g11980 ( 
.A1(n_11794),
.A2(n_4698),
.B(n_4697),
.Y(n_11980)
);

OAI321xp33_ASAP7_75t_L g11981 ( 
.A1(n_11781),
.A2(n_285),
.A3(n_287),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_11981)
);

AOI21xp5_ASAP7_75t_L g11982 ( 
.A1(n_11795),
.A2(n_4701),
.B(n_4699),
.Y(n_11982)
);

AOI21x1_ASAP7_75t_L g11983 ( 
.A1(n_11299),
.A2(n_4704),
.B(n_4703),
.Y(n_11983)
);

NOR2xp33_ASAP7_75t_L g11984 ( 
.A(n_11915),
.B(n_4707),
.Y(n_11984)
);

BUFx2_ASAP7_75t_L g11985 ( 
.A(n_11435),
.Y(n_11985)
);

AND2x4_ASAP7_75t_L g11986 ( 
.A(n_11555),
.B(n_11651),
.Y(n_11986)
);

NAND2xp5_ASAP7_75t_SL g11987 ( 
.A(n_11653),
.B(n_4708),
.Y(n_11987)
);

AND2x2_ASAP7_75t_L g11988 ( 
.A(n_11598),
.B(n_4709),
.Y(n_11988)
);

NAND2xp5_ASAP7_75t_L g11989 ( 
.A(n_11708),
.B(n_284),
.Y(n_11989)
);

OAI21xp5_ASAP7_75t_L g11990 ( 
.A1(n_11368),
.A2(n_285),
.B(n_286),
.Y(n_11990)
);

INVx1_ASAP7_75t_L g11991 ( 
.A(n_11357),
.Y(n_11991)
);

NAND2xp5_ASAP7_75t_SL g11992 ( 
.A(n_11659),
.B(n_4710),
.Y(n_11992)
);

AOI21xp5_ASAP7_75t_L g11993 ( 
.A1(n_11796),
.A2(n_11804),
.B(n_11803),
.Y(n_11993)
);

AND2x2_ASAP7_75t_L g11994 ( 
.A(n_11780),
.B(n_4711),
.Y(n_11994)
);

OAI22xp5_ASAP7_75t_L g11995 ( 
.A1(n_11753),
.A2(n_11779),
.B1(n_11456),
.B2(n_11518),
.Y(n_11995)
);

O2A1O1Ixp5_ASAP7_75t_L g11996 ( 
.A1(n_11507),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_11996)
);

AOI21xp5_ASAP7_75t_L g11997 ( 
.A1(n_11805),
.A2(n_4713),
.B(n_4712),
.Y(n_11997)
);

NAND2xp5_ASAP7_75t_L g11998 ( 
.A(n_11808),
.B(n_290),
.Y(n_11998)
);

BUFx4f_ASAP7_75t_L g11999 ( 
.A(n_11614),
.Y(n_11999)
);

AOI21xp5_ASAP7_75t_L g12000 ( 
.A1(n_11809),
.A2(n_4718),
.B(n_4716),
.Y(n_12000)
);

NOR2xp33_ASAP7_75t_L g12001 ( 
.A(n_11923),
.B(n_4719),
.Y(n_12001)
);

OAI21xp5_ASAP7_75t_L g12002 ( 
.A1(n_11373),
.A2(n_290),
.B(n_291),
.Y(n_12002)
);

INVx2_ASAP7_75t_L g12003 ( 
.A(n_11800),
.Y(n_12003)
);

BUFx4f_ASAP7_75t_L g12004 ( 
.A(n_11648),
.Y(n_12004)
);

AOI22xp5_ASAP7_75t_L g12005 ( 
.A1(n_11471),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_12005)
);

AOI21xp5_ASAP7_75t_L g12006 ( 
.A1(n_11813),
.A2(n_4722),
.B(n_4721),
.Y(n_12006)
);

NOR2xp33_ASAP7_75t_L g12007 ( 
.A(n_11907),
.B(n_11538),
.Y(n_12007)
);

AOI22xp5_ASAP7_75t_L g12008 ( 
.A1(n_11462),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_12008)
);

AOI21xp5_ASAP7_75t_L g12009 ( 
.A1(n_11815),
.A2(n_4724),
.B(n_4723),
.Y(n_12009)
);

AOI21xp5_ASAP7_75t_L g12010 ( 
.A1(n_11818),
.A2(n_11821),
.B(n_11819),
.Y(n_12010)
);

O2A1O1Ixp33_ASAP7_75t_L g12011 ( 
.A1(n_11783),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_12011)
);

AOI22xp5_ASAP7_75t_L g12012 ( 
.A1(n_11748),
.A2(n_11729),
.B1(n_11630),
.B2(n_11358),
.Y(n_12012)
);

OAI21xp5_ASAP7_75t_L g12013 ( 
.A1(n_11308),
.A2(n_295),
.B(n_296),
.Y(n_12013)
);

BUFx8_ASAP7_75t_L g12014 ( 
.A(n_11724),
.Y(n_12014)
);

INVx1_ASAP7_75t_L g12015 ( 
.A(n_11359),
.Y(n_12015)
);

NOR3xp33_ASAP7_75t_L g12016 ( 
.A(n_11489),
.B(n_11519),
.C(n_11771),
.Y(n_12016)
);

AOI21xp5_ASAP7_75t_L g12017 ( 
.A1(n_11823),
.A2(n_11826),
.B(n_11824),
.Y(n_12017)
);

OAI22xp5_ASAP7_75t_L g12018 ( 
.A1(n_11799),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_12018)
);

AOI21xp5_ASAP7_75t_L g12019 ( 
.A1(n_11828),
.A2(n_4726),
.B(n_4725),
.Y(n_12019)
);

NOR2xp33_ASAP7_75t_L g12020 ( 
.A(n_11657),
.B(n_4727),
.Y(n_12020)
);

AOI21xp5_ASAP7_75t_L g12021 ( 
.A1(n_11830),
.A2(n_4729),
.B(n_4728),
.Y(n_12021)
);

NAND2xp5_ASAP7_75t_L g12022 ( 
.A(n_11839),
.B(n_297),
.Y(n_12022)
);

AND2x2_ASAP7_75t_L g12023 ( 
.A(n_11582),
.B(n_4730),
.Y(n_12023)
);

O2A1O1Ixp5_ASAP7_75t_SL g12024 ( 
.A1(n_11924),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_12024)
);

NOR2xp33_ASAP7_75t_L g12025 ( 
.A(n_11755),
.B(n_4731),
.Y(n_12025)
);

NOR2xp33_ASAP7_75t_L g12026 ( 
.A(n_11559),
.B(n_4733),
.Y(n_12026)
);

NAND2xp5_ASAP7_75t_L g12027 ( 
.A(n_11840),
.B(n_300),
.Y(n_12027)
);

OAI22xp5_ASAP7_75t_L g12028 ( 
.A1(n_11811),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_12028)
);

AOI21xp5_ASAP7_75t_L g12029 ( 
.A1(n_11843),
.A2(n_4735),
.B(n_4734),
.Y(n_12029)
);

INVxp67_ASAP7_75t_L g12030 ( 
.A(n_11352),
.Y(n_12030)
);

NAND2xp5_ASAP7_75t_L g12031 ( 
.A(n_11845),
.B(n_301),
.Y(n_12031)
);

INVx1_ASAP7_75t_L g12032 ( 
.A(n_11360),
.Y(n_12032)
);

AOI21xp5_ASAP7_75t_L g12033 ( 
.A1(n_11850),
.A2(n_4738),
.B(n_4737),
.Y(n_12033)
);

AOI21x1_ASAP7_75t_L g12034 ( 
.A1(n_11309),
.A2(n_4740),
.B(n_4739),
.Y(n_12034)
);

O2A1O1Ixp33_ASAP7_75t_L g12035 ( 
.A1(n_11816),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_12035)
);

A2O1A1Ixp33_ASAP7_75t_L g12036 ( 
.A1(n_11760),
.A2(n_306),
.B(n_304),
.C(n_305),
.Y(n_12036)
);

INVx2_ASAP7_75t_L g12037 ( 
.A(n_11806),
.Y(n_12037)
);

AOI21xp5_ASAP7_75t_L g12038 ( 
.A1(n_11851),
.A2(n_4743),
.B(n_4741),
.Y(n_12038)
);

OAI22xp5_ASAP7_75t_L g12039 ( 
.A1(n_11835),
.A2(n_309),
.B1(n_306),
.B2(n_308),
.Y(n_12039)
);

NOR3xp33_ASAP7_75t_L g12040 ( 
.A(n_11787),
.B(n_308),
.C(n_309),
.Y(n_12040)
);

NOR2x1_ASAP7_75t_L g12041 ( 
.A(n_11759),
.B(n_310),
.Y(n_12041)
);

AOI21xp5_ASAP7_75t_L g12042 ( 
.A1(n_11853),
.A2(n_11857),
.B(n_11855),
.Y(n_12042)
);

NOR2x1_ASAP7_75t_L g12043 ( 
.A(n_11661),
.B(n_310),
.Y(n_12043)
);

OAI21xp5_ASAP7_75t_L g12044 ( 
.A1(n_11328),
.A2(n_11638),
.B(n_11371),
.Y(n_12044)
);

NOR2xp33_ASAP7_75t_L g12045 ( 
.A(n_11426),
.B(n_4744),
.Y(n_12045)
);

OAI321xp33_ASAP7_75t_L g12046 ( 
.A1(n_11873),
.A2(n_313),
.A3(n_315),
.B1(n_311),
.B2(n_312),
.C(n_314),
.Y(n_12046)
);

AOI22xp5_ASAP7_75t_L g12047 ( 
.A1(n_11485),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_12047)
);

OAI21xp5_ASAP7_75t_L g12048 ( 
.A1(n_11375),
.A2(n_315),
.B(n_316),
.Y(n_12048)
);

OAI21xp5_ASAP7_75t_L g12049 ( 
.A1(n_11663),
.A2(n_11667),
.B(n_11844),
.Y(n_12049)
);

INVx1_ASAP7_75t_SL g12050 ( 
.A(n_11466),
.Y(n_12050)
);

NAND2xp5_ASAP7_75t_L g12051 ( 
.A(n_11858),
.B(n_11862),
.Y(n_12051)
);

NAND2xp5_ASAP7_75t_SL g12052 ( 
.A(n_11546),
.B(n_4745),
.Y(n_12052)
);

AOI21xp5_ASAP7_75t_L g12053 ( 
.A1(n_11863),
.A2(n_4747),
.B(n_4746),
.Y(n_12053)
);

AOI21xp33_ASAP7_75t_L g12054 ( 
.A1(n_11713),
.A2(n_316),
.B(n_317),
.Y(n_12054)
);

AOI21xp5_ASAP7_75t_L g12055 ( 
.A1(n_11867),
.A2(n_4749),
.B(n_4748),
.Y(n_12055)
);

AND2x4_ASAP7_75t_L g12056 ( 
.A(n_11429),
.B(n_4750),
.Y(n_12056)
);

A2O1A1Ixp33_ASAP7_75t_L g12057 ( 
.A1(n_11849),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_12057)
);

AOI21xp5_ASAP7_75t_L g12058 ( 
.A1(n_11868),
.A2(n_4753),
.B(n_4752),
.Y(n_12058)
);

A2O1A1Ixp33_ASAP7_75t_L g12059 ( 
.A1(n_11861),
.A2(n_321),
.B(n_318),
.C(n_320),
.Y(n_12059)
);

AO21x1_ASAP7_75t_L g12060 ( 
.A1(n_11917),
.A2(n_321),
.B(n_322),
.Y(n_12060)
);

NAND2xp5_ASAP7_75t_L g12061 ( 
.A(n_11874),
.B(n_322),
.Y(n_12061)
);

AOI21xp5_ASAP7_75t_L g12062 ( 
.A1(n_11875),
.A2(n_4755),
.B(n_4754),
.Y(n_12062)
);

INVx2_ASAP7_75t_L g12063 ( 
.A(n_11817),
.Y(n_12063)
);

A2O1A1Ixp33_ASAP7_75t_L g12064 ( 
.A1(n_11872),
.A2(n_325),
.B(n_323),
.C(n_324),
.Y(n_12064)
);

NAND2xp5_ASAP7_75t_L g12065 ( 
.A(n_11876),
.B(n_323),
.Y(n_12065)
);

INVx2_ASAP7_75t_L g12066 ( 
.A(n_11820),
.Y(n_12066)
);

NAND2xp5_ASAP7_75t_L g12067 ( 
.A(n_11883),
.B(n_324),
.Y(n_12067)
);

BUFx2_ASAP7_75t_L g12068 ( 
.A(n_11492),
.Y(n_12068)
);

AOI22xp5_ASAP7_75t_L g12069 ( 
.A1(n_11326),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_12069)
);

O2A1O1Ixp33_ASAP7_75t_L g12070 ( 
.A1(n_11884),
.A2(n_328),
.B(n_326),
.C(n_327),
.Y(n_12070)
);

NAND2xp5_ASAP7_75t_SL g12071 ( 
.A(n_11547),
.B(n_4756),
.Y(n_12071)
);

CKINVDCx8_ASAP7_75t_R g12072 ( 
.A(n_11366),
.Y(n_12072)
);

INVx2_ASAP7_75t_L g12073 ( 
.A(n_11829),
.Y(n_12073)
);

AOI22xp33_ASAP7_75t_L g12074 ( 
.A1(n_11911),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_12074)
);

NAND2xp5_ASAP7_75t_L g12075 ( 
.A(n_11886),
.B(n_11889),
.Y(n_12075)
);

NAND2xp5_ASAP7_75t_L g12076 ( 
.A(n_11894),
.B(n_329),
.Y(n_12076)
);

NAND2xp5_ASAP7_75t_L g12077 ( 
.A(n_11895),
.B(n_331),
.Y(n_12077)
);

NAND2xp5_ASAP7_75t_L g12078 ( 
.A(n_11898),
.B(n_331),
.Y(n_12078)
);

BUFx8_ASAP7_75t_L g12079 ( 
.A(n_11354),
.Y(n_12079)
);

INVx1_ASAP7_75t_L g12080 ( 
.A(n_11367),
.Y(n_12080)
);

NAND2xp5_ASAP7_75t_L g12081 ( 
.A(n_11899),
.B(n_332),
.Y(n_12081)
);

INVx2_ASAP7_75t_L g12082 ( 
.A(n_11841),
.Y(n_12082)
);

AOI21xp5_ASAP7_75t_L g12083 ( 
.A1(n_11901),
.A2(n_4758),
.B(n_4757),
.Y(n_12083)
);

AOI21xp5_ASAP7_75t_L g12084 ( 
.A1(n_11903),
.A2(n_4760),
.B(n_4759),
.Y(n_12084)
);

AOI21xp5_ASAP7_75t_L g12085 ( 
.A1(n_11910),
.A2(n_4762),
.B(n_4761),
.Y(n_12085)
);

AOI21xp5_ASAP7_75t_L g12086 ( 
.A1(n_11913),
.A2(n_4764),
.B(n_4763),
.Y(n_12086)
);

AOI21xp5_ASAP7_75t_L g12087 ( 
.A1(n_11918),
.A2(n_4767),
.B(n_4766),
.Y(n_12087)
);

O2A1O1Ixp33_ASAP7_75t_L g12088 ( 
.A1(n_11922),
.A2(n_11758),
.B(n_11439),
.C(n_11568),
.Y(n_12088)
);

INVx4_ASAP7_75t_L g12089 ( 
.A(n_11385),
.Y(n_12089)
);

AOI21xp5_ASAP7_75t_L g12090 ( 
.A1(n_11925),
.A2(n_4770),
.B(n_4769),
.Y(n_12090)
);

AND2x2_ASAP7_75t_L g12091 ( 
.A(n_11810),
.B(n_4772),
.Y(n_12091)
);

AOI21xp5_ASAP7_75t_L g12092 ( 
.A1(n_11927),
.A2(n_4774),
.B(n_4773),
.Y(n_12092)
);

NAND2xp5_ASAP7_75t_L g12093 ( 
.A(n_11929),
.B(n_332),
.Y(n_12093)
);

INVx2_ASAP7_75t_SL g12094 ( 
.A(n_11523),
.Y(n_12094)
);

A2O1A1Ixp33_ASAP7_75t_L g12095 ( 
.A1(n_11484),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_12095)
);

NAND2xp5_ASAP7_75t_SL g12096 ( 
.A(n_11556),
.B(n_4775),
.Y(n_12096)
);

BUFx6f_ASAP7_75t_L g12097 ( 
.A(n_11699),
.Y(n_12097)
);

NOR2xp33_ASAP7_75t_L g12098 ( 
.A(n_11619),
.B(n_11761),
.Y(n_12098)
);

OAI21x1_ASAP7_75t_L g12099 ( 
.A1(n_11549),
.A2(n_4779),
.B(n_4777),
.Y(n_12099)
);

AND2x2_ASAP7_75t_L g12100 ( 
.A(n_11846),
.B(n_4780),
.Y(n_12100)
);

BUFx6f_ASAP7_75t_L g12101 ( 
.A(n_11699),
.Y(n_12101)
);

O2A1O1Ixp33_ASAP7_75t_L g12102 ( 
.A1(n_11776),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_12102)
);

AND2x4_ASAP7_75t_L g12103 ( 
.A(n_11351),
.B(n_4781),
.Y(n_12103)
);

NOR2xp33_ASAP7_75t_L g12104 ( 
.A(n_11743),
.B(n_4782),
.Y(n_12104)
);

O2A1O1Ixp33_ASAP7_75t_L g12105 ( 
.A1(n_11530),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_12105)
);

OAI22xp5_ASAP7_75t_L g12106 ( 
.A1(n_11469),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_12106)
);

OAI22xp5_ASAP7_75t_L g12107 ( 
.A1(n_11768),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_12107)
);

NAND2xp5_ASAP7_75t_L g12108 ( 
.A(n_11488),
.B(n_339),
.Y(n_12108)
);

AOI21x1_ASAP7_75t_L g12109 ( 
.A1(n_11418),
.A2(n_4784),
.B(n_4783),
.Y(n_12109)
);

OAI22xp5_ASAP7_75t_L g12110 ( 
.A1(n_11710),
.A2(n_344),
.B1(n_340),
.B2(n_343),
.Y(n_12110)
);

OAI22xp5_ASAP7_75t_L g12111 ( 
.A1(n_11735),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_12111)
);

NAND2xp5_ASAP7_75t_L g12112 ( 
.A(n_11558),
.B(n_346),
.Y(n_12112)
);

INVxp67_ASAP7_75t_L g12113 ( 
.A(n_11396),
.Y(n_12113)
);

A2O1A1Ixp33_ASAP7_75t_L g12114 ( 
.A1(n_11745),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_12114)
);

NOR2xp33_ASAP7_75t_L g12115 ( 
.A(n_11382),
.B(n_4785),
.Y(n_12115)
);

OAI21xp5_ASAP7_75t_L g12116 ( 
.A1(n_11563),
.A2(n_347),
.B(n_349),
.Y(n_12116)
);

NOR2xp67_ASAP7_75t_L g12117 ( 
.A(n_11837),
.B(n_4786),
.Y(n_12117)
);

INVx1_ASAP7_75t_L g12118 ( 
.A(n_11369),
.Y(n_12118)
);

NOR2x1p5_ASAP7_75t_SL g12119 ( 
.A(n_11550),
.B(n_4787),
.Y(n_12119)
);

AOI22x1_ASAP7_75t_L g12120 ( 
.A1(n_11832),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_12120)
);

BUFx2_ASAP7_75t_L g12121 ( 
.A(n_11551),
.Y(n_12121)
);

NAND3xp33_ASAP7_75t_L g12122 ( 
.A(n_11406),
.B(n_352),
.C(n_353),
.Y(n_12122)
);

NAND2xp5_ASAP7_75t_L g12123 ( 
.A(n_11567),
.B(n_353),
.Y(n_12123)
);

NOR2xp33_ASAP7_75t_L g12124 ( 
.A(n_11436),
.B(n_4788),
.Y(n_12124)
);

NAND2xp5_ASAP7_75t_L g12125 ( 
.A(n_11569),
.B(n_354),
.Y(n_12125)
);

INVx1_ASAP7_75t_L g12126 ( 
.A(n_11376),
.Y(n_12126)
);

NAND2xp5_ASAP7_75t_L g12127 ( 
.A(n_11570),
.B(n_354),
.Y(n_12127)
);

INVx4_ASAP7_75t_L g12128 ( 
.A(n_11394),
.Y(n_12128)
);

OAI21xp5_ASAP7_75t_L g12129 ( 
.A1(n_11575),
.A2(n_355),
.B(n_356),
.Y(n_12129)
);

AOI21xp5_ASAP7_75t_L g12130 ( 
.A1(n_11764),
.A2(n_4791),
.B(n_4789),
.Y(n_12130)
);

OAI22xp5_ASAP7_75t_L g12131 ( 
.A1(n_11295),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_12131)
);

AOI21xp5_ASAP7_75t_L g12132 ( 
.A1(n_11581),
.A2(n_4793),
.B(n_4792),
.Y(n_12132)
);

AOI21xp5_ASAP7_75t_L g12133 ( 
.A1(n_11583),
.A2(n_4796),
.B(n_4795),
.Y(n_12133)
);

A2O1A1Ixp33_ASAP7_75t_L g12134 ( 
.A1(n_11481),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_12134)
);

AOI21xp5_ASAP7_75t_L g12135 ( 
.A1(n_11589),
.A2(n_4798),
.B(n_4797),
.Y(n_12135)
);

AOI21xp5_ASAP7_75t_L g12136 ( 
.A1(n_11591),
.A2(n_4801),
.B(n_4800),
.Y(n_12136)
);

A2O1A1Ixp33_ASAP7_75t_L g12137 ( 
.A1(n_11637),
.A2(n_361),
.B(n_358),
.C(n_360),
.Y(n_12137)
);

NAND2xp5_ASAP7_75t_L g12138 ( 
.A(n_11592),
.B(n_360),
.Y(n_12138)
);

INVx2_ASAP7_75t_L g12139 ( 
.A(n_11847),
.Y(n_12139)
);

NAND2xp5_ASAP7_75t_L g12140 ( 
.A(n_11601),
.B(n_361),
.Y(n_12140)
);

AOI21xp5_ASAP7_75t_L g12141 ( 
.A1(n_11602),
.A2(n_4803),
.B(n_4802),
.Y(n_12141)
);

BUFx6f_ASAP7_75t_L g12142 ( 
.A(n_11500),
.Y(n_12142)
);

AOI21xp5_ASAP7_75t_L g12143 ( 
.A1(n_11603),
.A2(n_4807),
.B(n_4804),
.Y(n_12143)
);

O2A1O1Ixp33_ASAP7_75t_L g12144 ( 
.A1(n_11552),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_12144)
);

NAND2xp5_ASAP7_75t_L g12145 ( 
.A(n_11606),
.B(n_362),
.Y(n_12145)
);

O2A1O1Ixp5_ASAP7_75t_L g12146 ( 
.A1(n_11633),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_12146)
);

NAND2xp5_ASAP7_75t_SL g12147 ( 
.A(n_11613),
.B(n_4808),
.Y(n_12147)
);

A2O1A1Ixp33_ASAP7_75t_L g12148 ( 
.A1(n_11495),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_12148)
);

A2O1A1Ixp33_ASAP7_75t_L g12149 ( 
.A1(n_11501),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_12149)
);

AND2x4_ASAP7_75t_L g12150 ( 
.A(n_11353),
.B(n_4809),
.Y(n_12150)
);

NAND2xp5_ASAP7_75t_L g12151 ( 
.A(n_11615),
.B(n_369),
.Y(n_12151)
);

INVx2_ASAP7_75t_L g12152 ( 
.A(n_11865),
.Y(n_12152)
);

AOI21xp5_ASAP7_75t_L g12153 ( 
.A1(n_11616),
.A2(n_11622),
.B(n_11620),
.Y(n_12153)
);

NAND2xp5_ASAP7_75t_SL g12154 ( 
.A(n_11631),
.B(n_4810),
.Y(n_12154)
);

BUFx4f_ASAP7_75t_L g12155 ( 
.A(n_11666),
.Y(n_12155)
);

NAND3xp33_ASAP7_75t_L g12156 ( 
.A(n_11410),
.B(n_369),
.C(n_370),
.Y(n_12156)
);

OAI22xp5_ASAP7_75t_L g12157 ( 
.A1(n_11775),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_12157)
);

O2A1O1Ixp5_ASAP7_75t_L g12158 ( 
.A1(n_11590),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_12158)
);

NOR2x1_ASAP7_75t_L g12159 ( 
.A(n_11652),
.B(n_373),
.Y(n_12159)
);

NAND2x1p5_ASAP7_75t_L g12160 ( 
.A(n_11869),
.B(n_11891),
.Y(n_12160)
);

AOI21xp5_ASAP7_75t_L g12161 ( 
.A1(n_11636),
.A2(n_4813),
.B(n_4812),
.Y(n_12161)
);

AOI22xp33_ASAP7_75t_L g12162 ( 
.A1(n_11584),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_12162)
);

NAND2xp5_ASAP7_75t_L g12163 ( 
.A(n_11532),
.B(n_374),
.Y(n_12163)
);

AOI22xp33_ASAP7_75t_L g12164 ( 
.A1(n_11595),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_12164)
);

NAND2xp5_ASAP7_75t_L g12165 ( 
.A(n_11458),
.B(n_377),
.Y(n_12165)
);

AOI21x1_ASAP7_75t_L g12166 ( 
.A1(n_11314),
.A2(n_4815),
.B(n_4814),
.Y(n_12166)
);

BUFx8_ASAP7_75t_L g12167 ( 
.A(n_11698),
.Y(n_12167)
);

INVx2_ASAP7_75t_L g12168 ( 
.A(n_11877),
.Y(n_12168)
);

OAI21x1_ASAP7_75t_L g12169 ( 
.A1(n_11566),
.A2(n_4817),
.B(n_4816),
.Y(n_12169)
);

NAND2xp5_ASAP7_75t_L g12170 ( 
.A(n_11461),
.B(n_378),
.Y(n_12170)
);

NOR2xp33_ASAP7_75t_L g12171 ( 
.A(n_11754),
.B(n_4818),
.Y(n_12171)
);

A2O1A1Ixp33_ASAP7_75t_L g12172 ( 
.A1(n_11535),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_12172)
);

A2O1A1Ixp33_ASAP7_75t_L g12173 ( 
.A1(n_11554),
.A2(n_11562),
.B(n_11571),
.C(n_11565),
.Y(n_12173)
);

AOI21xp5_ASAP7_75t_L g12174 ( 
.A1(n_11746),
.A2(n_4820),
.B(n_4819),
.Y(n_12174)
);

AOI221xp5_ASAP7_75t_L g12175 ( 
.A1(n_11496),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.C(n_383),
.Y(n_12175)
);

AOI21xp5_ASAP7_75t_L g12176 ( 
.A1(n_11746),
.A2(n_4822),
.B(n_4821),
.Y(n_12176)
);

OAI21xp5_ASAP7_75t_L g12177 ( 
.A1(n_11304),
.A2(n_381),
.B(n_384),
.Y(n_12177)
);

BUFx2_ASAP7_75t_L g12178 ( 
.A(n_11737),
.Y(n_12178)
);

OAI21xp33_ASAP7_75t_L g12179 ( 
.A1(n_11408),
.A2(n_384),
.B(n_385),
.Y(n_12179)
);

AOI21xp5_ASAP7_75t_L g12180 ( 
.A1(n_11738),
.A2(n_4824),
.B(n_4823),
.Y(n_12180)
);

NOR2xp67_ASAP7_75t_L g12181 ( 
.A(n_11573),
.B(n_4825),
.Y(n_12181)
);

AOI21xp5_ASAP7_75t_L g12182 ( 
.A1(n_11744),
.A2(n_4827),
.B(n_4826),
.Y(n_12182)
);

AOI21xp5_ASAP7_75t_L g12183 ( 
.A1(n_11716),
.A2(n_4829),
.B(n_4828),
.Y(n_12183)
);

NOR2xp33_ASAP7_75t_L g12184 ( 
.A(n_11756),
.B(n_4830),
.Y(n_12184)
);

HB1xp67_ASAP7_75t_L g12185 ( 
.A(n_11383),
.Y(n_12185)
);

OAI21xp33_ASAP7_75t_SL g12186 ( 
.A1(n_11411),
.A2(n_386),
.B(n_387),
.Y(n_12186)
);

AND2x4_ASAP7_75t_L g12187 ( 
.A(n_11607),
.B(n_11389),
.Y(n_12187)
);

INVx2_ASAP7_75t_L g12188 ( 
.A(n_11885),
.Y(n_12188)
);

AOI21xp5_ASAP7_75t_L g12189 ( 
.A1(n_11727),
.A2(n_11732),
.B(n_11593),
.Y(n_12189)
);

AOI21xp5_ASAP7_75t_L g12190 ( 
.A1(n_11585),
.A2(n_4832),
.B(n_4831),
.Y(n_12190)
);

INVxp67_ASAP7_75t_L g12191 ( 
.A(n_11689),
.Y(n_12191)
);

INVx2_ASAP7_75t_SL g12192 ( 
.A(n_11526),
.Y(n_12192)
);

NAND2xp5_ASAP7_75t_L g12193 ( 
.A(n_11774),
.B(n_386),
.Y(n_12193)
);

AOI22xp5_ASAP7_75t_L g12194 ( 
.A1(n_11645),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_12194)
);

AOI21xp5_ASAP7_75t_L g12195 ( 
.A1(n_11596),
.A2(n_4834),
.B(n_4833),
.Y(n_12195)
);

AOI21xp5_ASAP7_75t_L g12196 ( 
.A1(n_11597),
.A2(n_4836),
.B(n_4835),
.Y(n_12196)
);

INVx1_ASAP7_75t_L g12197 ( 
.A(n_11387),
.Y(n_12197)
);

BUFx2_ASAP7_75t_L g12198 ( 
.A(n_11522),
.Y(n_12198)
);

BUFx2_ASAP7_75t_L g12199 ( 
.A(n_11697),
.Y(n_12199)
);

NOR2x1_ASAP7_75t_L g12200 ( 
.A(n_11441),
.B(n_389),
.Y(n_12200)
);

NAND2xp5_ASAP7_75t_L g12201 ( 
.A(n_11770),
.B(n_390),
.Y(n_12201)
);

NOR2xp33_ASAP7_75t_L g12202 ( 
.A(n_11363),
.B(n_4837),
.Y(n_12202)
);

NAND2xp5_ASAP7_75t_L g12203 ( 
.A(n_11892),
.B(n_391),
.Y(n_12203)
);

NAND2xp5_ASAP7_75t_L g12204 ( 
.A(n_11928),
.B(n_391),
.Y(n_12204)
);

BUFx2_ASAP7_75t_L g12205 ( 
.A(n_11740),
.Y(n_12205)
);

A2O1A1Ixp33_ASAP7_75t_L g12206 ( 
.A1(n_11576),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_12206)
);

AOI21xp5_ASAP7_75t_L g12207 ( 
.A1(n_11579),
.A2(n_11751),
.B(n_11750),
.Y(n_12207)
);

NOR2xp33_ASAP7_75t_L g12208 ( 
.A(n_11766),
.B(n_4838),
.Y(n_12208)
);

INVx2_ASAP7_75t_L g12209 ( 
.A(n_11386),
.Y(n_12209)
);

AOI22xp5_ASAP7_75t_L g12210 ( 
.A1(n_11685),
.A2(n_395),
.B1(n_392),
.B2(n_394),
.Y(n_12210)
);

O2A1O1Ixp33_ASAP7_75t_L g12211 ( 
.A1(n_11379),
.A2(n_11380),
.B(n_11720),
.C(n_11684),
.Y(n_12211)
);

AOI21xp5_ASAP7_75t_L g12212 ( 
.A1(n_11718),
.A2(n_4840),
.B(n_4839),
.Y(n_12212)
);

AOI21x1_ASAP7_75t_L g12213 ( 
.A1(n_11712),
.A2(n_4843),
.B(n_4842),
.Y(n_12213)
);

NAND2xp5_ASAP7_75t_L g12214 ( 
.A(n_11533),
.B(n_395),
.Y(n_12214)
);

NAND2xp5_ASAP7_75t_SL g12215 ( 
.A(n_11836),
.B(n_4844),
.Y(n_12215)
);

AOI21xp5_ASAP7_75t_L g12216 ( 
.A1(n_11723),
.A2(n_4847),
.B(n_4846),
.Y(n_12216)
);

AND2x2_ASAP7_75t_L g12217 ( 
.A(n_11854),
.B(n_4848),
.Y(n_12217)
);

NOR2xp33_ASAP7_75t_L g12218 ( 
.A(n_11777),
.B(n_4850),
.Y(n_12218)
);

A2O1A1Ixp33_ASAP7_75t_L g12219 ( 
.A1(n_11586),
.A2(n_398),
.B(n_396),
.C(n_397),
.Y(n_12219)
);

AOI21xp5_ASAP7_75t_L g12220 ( 
.A1(n_11726),
.A2(n_4855),
.B(n_4854),
.Y(n_12220)
);

INVx2_ASAP7_75t_L g12221 ( 
.A(n_11390),
.Y(n_12221)
);

NAND2xp5_ASAP7_75t_L g12222 ( 
.A(n_11534),
.B(n_396),
.Y(n_12222)
);

AOI21xp5_ASAP7_75t_L g12223 ( 
.A1(n_11749),
.A2(n_4857),
.B(n_4856),
.Y(n_12223)
);

OAI21xp33_ASAP7_75t_L g12224 ( 
.A1(n_11447),
.A2(n_397),
.B(n_399),
.Y(n_12224)
);

NAND2xp5_ASAP7_75t_L g12225 ( 
.A(n_11537),
.B(n_11540),
.Y(n_12225)
);

BUFx2_ASAP7_75t_L g12226 ( 
.A(n_11725),
.Y(n_12226)
);

NOR2x1p5_ASAP7_75t_SL g12227 ( 
.A(n_11405),
.B(n_4858),
.Y(n_12227)
);

NAND2x1p5_ASAP7_75t_L g12228 ( 
.A(n_11612),
.B(n_4859),
.Y(n_12228)
);

AOI21xp5_ASAP7_75t_L g12229 ( 
.A1(n_11715),
.A2(n_4861),
.B(n_4860),
.Y(n_12229)
);

O2A1O1Ixp5_ASAP7_75t_L g12230 ( 
.A1(n_11561),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_12230)
);

NAND3xp33_ASAP7_75t_L g12231 ( 
.A(n_11574),
.B(n_400),
.C(n_402),
.Y(n_12231)
);

INVx2_ASAP7_75t_L g12232 ( 
.A(n_11395),
.Y(n_12232)
);

AND2x2_ASAP7_75t_L g12233 ( 
.A(n_11856),
.B(n_4862),
.Y(n_12233)
);

O2A1O1Ixp33_ASAP7_75t_L g12234 ( 
.A1(n_11736),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_12234)
);

NOR3xp33_ASAP7_75t_L g12235 ( 
.A(n_11642),
.B(n_403),
.C(n_404),
.Y(n_12235)
);

OAI21xp5_ASAP7_75t_L g12236 ( 
.A1(n_11599),
.A2(n_405),
.B(n_406),
.Y(n_12236)
);

INVx3_ASAP7_75t_L g12237 ( 
.A(n_11364),
.Y(n_12237)
);

NAND2xp5_ASAP7_75t_L g12238 ( 
.A(n_11545),
.B(n_405),
.Y(n_12238)
);

OAI21xp5_ASAP7_75t_L g12239 ( 
.A1(n_11610),
.A2(n_406),
.B(n_407),
.Y(n_12239)
);

BUFx3_ASAP7_75t_L g12240 ( 
.A(n_11588),
.Y(n_12240)
);

AOI21xp5_ASAP7_75t_L g12241 ( 
.A1(n_11587),
.A2(n_4864),
.B(n_4863),
.Y(n_12241)
);

NAND2xp5_ASAP7_75t_L g12242 ( 
.A(n_11403),
.B(n_11291),
.Y(n_12242)
);

AOI21xp5_ASAP7_75t_L g12243 ( 
.A1(n_11440),
.A2(n_4866),
.B(n_4865),
.Y(n_12243)
);

AO22x1_ASAP7_75t_L g12244 ( 
.A1(n_11897),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_12244)
);

NAND2xp5_ASAP7_75t_L g12245 ( 
.A(n_11292),
.B(n_408),
.Y(n_12245)
);

HB1xp67_ASAP7_75t_L g12246 ( 
.A(n_11393),
.Y(n_12246)
);

OAI22xp5_ASAP7_75t_L g12247 ( 
.A1(n_11425),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_12247)
);

AOI21xp5_ASAP7_75t_L g12248 ( 
.A1(n_11594),
.A2(n_4868),
.B(n_4867),
.Y(n_12248)
);

AOI22xp5_ASAP7_75t_L g12249 ( 
.A1(n_11763),
.A2(n_413),
.B1(n_410),
.B2(n_412),
.Y(n_12249)
);

CKINVDCx10_ASAP7_75t_R g12250 ( 
.A(n_11666),
.Y(n_12250)
);

AOI21xp5_ASAP7_75t_L g12251 ( 
.A1(n_11494),
.A2(n_4871),
.B(n_4870),
.Y(n_12251)
);

O2A1O1Ixp5_ASAP7_75t_L g12252 ( 
.A1(n_11649),
.A2(n_11564),
.B(n_11695),
.C(n_11680),
.Y(n_12252)
);

AOI21xp5_ASAP7_75t_L g12253 ( 
.A1(n_11377),
.A2(n_4874),
.B(n_4872),
.Y(n_12253)
);

BUFx8_ASAP7_75t_L g12254 ( 
.A(n_11860),
.Y(n_12254)
);

INVx1_ASAP7_75t_L g12255 ( 
.A(n_11397),
.Y(n_12255)
);

NAND2xp5_ASAP7_75t_L g12256 ( 
.A(n_11296),
.B(n_412),
.Y(n_12256)
);

AO22x1_ASAP7_75t_L g12257 ( 
.A1(n_11897),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_12257)
);

NAND2xp5_ASAP7_75t_L g12258 ( 
.A(n_11297),
.B(n_414),
.Y(n_12258)
);

INVx3_ASAP7_75t_L g12259 ( 
.A(n_11560),
.Y(n_12259)
);

HB1xp67_ASAP7_75t_L g12260 ( 
.A(n_11400),
.Y(n_12260)
);

NAND2xp5_ASAP7_75t_L g12261 ( 
.A(n_11298),
.B(n_11300),
.Y(n_12261)
);

OAI22xp5_ASAP7_75t_L g12262 ( 
.A1(n_11384),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_12262)
);

AOI22xp5_ASAP7_75t_L g12263 ( 
.A1(n_11778),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_12263)
);

AOI21xp5_ASAP7_75t_L g12264 ( 
.A1(n_11332),
.A2(n_4877),
.B(n_4875),
.Y(n_12264)
);

NOR3xp33_ASAP7_75t_L g12265 ( 
.A(n_11640),
.B(n_418),
.C(n_419),
.Y(n_12265)
);

A2O1A1Ixp33_ASAP7_75t_L g12266 ( 
.A1(n_11668),
.A2(n_422),
.B(n_420),
.C(n_421),
.Y(n_12266)
);

NAND2xp5_ASAP7_75t_L g12267 ( 
.A(n_11301),
.B(n_420),
.Y(n_12267)
);

A2O1A1Ixp33_ASAP7_75t_L g12268 ( 
.A1(n_11676),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_12268)
);

NAND2xp5_ASAP7_75t_L g12269 ( 
.A(n_11302),
.B(n_423),
.Y(n_12269)
);

NAND2xp5_ASAP7_75t_L g12270 ( 
.A(n_11305),
.B(n_424),
.Y(n_12270)
);

NAND2xp5_ASAP7_75t_L g12271 ( 
.A(n_11310),
.B(n_424),
.Y(n_12271)
);

NAND2xp5_ASAP7_75t_L g12272 ( 
.A(n_11312),
.B(n_425),
.Y(n_12272)
);

NOR2xp33_ASAP7_75t_SL g12273 ( 
.A(n_11765),
.B(n_4880),
.Y(n_12273)
);

NAND2xp5_ASAP7_75t_L g12274 ( 
.A(n_11315),
.B(n_425),
.Y(n_12274)
);

NOR3xp33_ASAP7_75t_L g12275 ( 
.A(n_11671),
.B(n_426),
.C(n_427),
.Y(n_12275)
);

AOI21xp5_ASAP7_75t_L g12276 ( 
.A1(n_11404),
.A2(n_4882),
.B(n_4881),
.Y(n_12276)
);

NAND2xp5_ASAP7_75t_L g12277 ( 
.A(n_11318),
.B(n_11319),
.Y(n_12277)
);

NOR2xp33_ASAP7_75t_L g12278 ( 
.A(n_11629),
.B(n_4884),
.Y(n_12278)
);

NOR2xp33_ASAP7_75t_L g12279 ( 
.A(n_11365),
.B(n_4885),
.Y(n_12279)
);

OR2x6_ASAP7_75t_L g12280 ( 
.A(n_11345),
.B(n_4886),
.Y(n_12280)
);

INVx2_ASAP7_75t_L g12281 ( 
.A(n_11419),
.Y(n_12281)
);

NOR2xp67_ASAP7_75t_L g12282 ( 
.A(n_11678),
.B(n_4887),
.Y(n_12282)
);

INVx3_ASAP7_75t_L g12283 ( 
.A(n_11370),
.Y(n_12283)
);

AOI21xp5_ASAP7_75t_L g12284 ( 
.A1(n_11343),
.A2(n_4889),
.B(n_4888),
.Y(n_12284)
);

INVx1_ASAP7_75t_L g12285 ( 
.A(n_11409),
.Y(n_12285)
);

NAND2xp5_ASAP7_75t_SL g12286 ( 
.A(n_11402),
.B(n_4890),
.Y(n_12286)
);

AOI21xp5_ASAP7_75t_L g12287 ( 
.A1(n_11388),
.A2(n_4892),
.B(n_4891),
.Y(n_12287)
);

INVx1_ASAP7_75t_L g12288 ( 
.A(n_11412),
.Y(n_12288)
);

BUFx2_ASAP7_75t_SL g12289 ( 
.A(n_11747),
.Y(n_12289)
);

AND2x2_ASAP7_75t_L g12290 ( 
.A(n_11879),
.B(n_4893),
.Y(n_12290)
);

AOI21xp5_ASAP7_75t_L g12291 ( 
.A1(n_11442),
.A2(n_4896),
.B(n_4894),
.Y(n_12291)
);

NAND2xp5_ASAP7_75t_L g12292 ( 
.A(n_11320),
.B(n_427),
.Y(n_12292)
);

OAI22xp33_ASAP7_75t_L g12293 ( 
.A1(n_11848),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_12293)
);

OAI22xp5_ASAP7_75t_L g12294 ( 
.A1(n_11650),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_12294)
);

NAND2xp5_ASAP7_75t_L g12295 ( 
.A(n_11321),
.B(n_431),
.Y(n_12295)
);

NAND2xp5_ASAP7_75t_L g12296 ( 
.A(n_11327),
.B(n_432),
.Y(n_12296)
);

OAI321xp33_ASAP7_75t_L g12297 ( 
.A1(n_11852),
.A2(n_434),
.A3(n_436),
.B1(n_432),
.B2(n_433),
.C(n_435),
.Y(n_12297)
);

INVx1_ASAP7_75t_SL g12298 ( 
.A(n_11742),
.Y(n_12298)
);

BUFx6f_ASAP7_75t_L g12299 ( 
.A(n_11477),
.Y(n_12299)
);

AOI21xp5_ASAP7_75t_L g12300 ( 
.A1(n_11453),
.A2(n_4898),
.B(n_4897),
.Y(n_12300)
);

INVx1_ASAP7_75t_SL g12301 ( 
.A(n_11289),
.Y(n_12301)
);

BUFx2_ASAP7_75t_L g12302 ( 
.A(n_11641),
.Y(n_12302)
);

BUFx12f_ASAP7_75t_L g12303 ( 
.A(n_11323),
.Y(n_12303)
);

BUFx4f_ASAP7_75t_L g12304 ( 
.A(n_11900),
.Y(n_12304)
);

AO22x1_ASAP7_75t_L g12305 ( 
.A1(n_11900),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_12305)
);

AOI21xp5_ASAP7_75t_L g12306 ( 
.A1(n_11480),
.A2(n_4900),
.B(n_4899),
.Y(n_12306)
);

NOR2xp33_ASAP7_75t_L g12307 ( 
.A(n_11307),
.B(n_4901),
.Y(n_12307)
);

O2A1O1Ixp33_ASAP7_75t_L g12308 ( 
.A1(n_11717),
.A2(n_438),
.B(n_436),
.C(n_437),
.Y(n_12308)
);

AOI21xp5_ASAP7_75t_L g12309 ( 
.A1(n_11707),
.A2(n_11341),
.B(n_11329),
.Y(n_12309)
);

NAND2xp5_ASAP7_75t_L g12310 ( 
.A(n_11344),
.B(n_438),
.Y(n_12310)
);

NAND2xp5_ASAP7_75t_SL g12311 ( 
.A(n_11703),
.B(n_4902),
.Y(n_12311)
);

NAND3xp33_ASAP7_75t_L g12312 ( 
.A(n_11878),
.B(n_439),
.C(n_440),
.Y(n_12312)
);

INVx2_ASAP7_75t_SL g12313 ( 
.A(n_11445),
.Y(n_12313)
);

O2A1O1Ixp33_ASAP7_75t_L g12314 ( 
.A1(n_11656),
.A2(n_442),
.B(n_440),
.C(n_441),
.Y(n_12314)
);

BUFx4f_ASAP7_75t_L g12315 ( 
.A(n_11900),
.Y(n_12315)
);

NAND2xp5_ASAP7_75t_L g12316 ( 
.A(n_11347),
.B(n_11348),
.Y(n_12316)
);

A2O1A1Ixp33_ASAP7_75t_L g12317 ( 
.A1(n_11722),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_12317)
);

NAND2xp5_ASAP7_75t_L g12318 ( 
.A(n_11423),
.B(n_443),
.Y(n_12318)
);

AOI21x1_ASAP7_75t_L g12319 ( 
.A1(n_11486),
.A2(n_4905),
.B(n_4903),
.Y(n_12319)
);

NAND2xp5_ASAP7_75t_L g12320 ( 
.A(n_11424),
.B(n_444),
.Y(n_12320)
);

AOI21xp5_ASAP7_75t_L g12321 ( 
.A1(n_11728),
.A2(n_4907),
.B(n_4906),
.Y(n_12321)
);

AOI21xp5_ASAP7_75t_L g12322 ( 
.A1(n_11470),
.A2(n_4911),
.B(n_4910),
.Y(n_12322)
);

INVxp67_ASAP7_75t_L g12323 ( 
.A(n_11604),
.Y(n_12323)
);

INVx3_ASAP7_75t_L g12324 ( 
.A(n_11479),
.Y(n_12324)
);

INVx1_ASAP7_75t_L g12325 ( 
.A(n_11413),
.Y(n_12325)
);

NAND2xp33_ASAP7_75t_L g12326 ( 
.A(n_11919),
.B(n_444),
.Y(n_12326)
);

AO221x1_ASAP7_75t_L g12327 ( 
.A1(n_11785),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.C(n_448),
.Y(n_12327)
);

OAI321xp33_ASAP7_75t_L g12328 ( 
.A1(n_11906),
.A2(n_447),
.A3(n_449),
.B1(n_445),
.B2(n_446),
.C(n_448),
.Y(n_12328)
);

AOI21xp5_ASAP7_75t_L g12329 ( 
.A1(n_11772),
.A2(n_4913),
.B(n_4912),
.Y(n_12329)
);

AOI21xp5_ASAP7_75t_L g12330 ( 
.A1(n_11542),
.A2(n_4915),
.B(n_4914),
.Y(n_12330)
);

INVx2_ASAP7_75t_L g12331 ( 
.A(n_11437),
.Y(n_12331)
);

NOR2xp33_ASAP7_75t_L g12332 ( 
.A(n_11734),
.B(n_4916),
.Y(n_12332)
);

AOI21xp33_ASAP7_75t_L g12333 ( 
.A1(n_11769),
.A2(n_449),
.B(n_450),
.Y(n_12333)
);

AOI21xp5_ASAP7_75t_L g12334 ( 
.A1(n_11617),
.A2(n_4918),
.B(n_4917),
.Y(n_12334)
);

AND2x6_ASAP7_75t_SL g12335 ( 
.A(n_11881),
.B(n_450),
.Y(n_12335)
);

NAND2xp5_ASAP7_75t_L g12336 ( 
.A(n_11449),
.B(n_451),
.Y(n_12336)
);

INVx4_ASAP7_75t_L g12337 ( 
.A(n_11322),
.Y(n_12337)
);

AOI21xp5_ASAP7_75t_L g12338 ( 
.A1(n_11580),
.A2(n_4920),
.B(n_4919),
.Y(n_12338)
);

NOR2xp33_ASAP7_75t_L g12339 ( 
.A(n_11475),
.B(n_4921),
.Y(n_12339)
);

INVx1_ASAP7_75t_SL g12340 ( 
.A(n_11628),
.Y(n_12340)
);

NAND2xp5_ASAP7_75t_L g12341 ( 
.A(n_11459),
.B(n_11467),
.Y(n_12341)
);

AOI21xp5_ASAP7_75t_L g12342 ( 
.A1(n_11621),
.A2(n_4923),
.B(n_4922),
.Y(n_12342)
);

INVx2_ASAP7_75t_SL g12343 ( 
.A(n_11483),
.Y(n_12343)
);

BUFx3_ASAP7_75t_L g12344 ( 
.A(n_11336),
.Y(n_12344)
);

AOI21xp5_ASAP7_75t_L g12345 ( 
.A1(n_11451),
.A2(n_11474),
.B(n_11317),
.Y(n_12345)
);

NOR2xp33_ASAP7_75t_L g12346 ( 
.A(n_11662),
.B(n_4924),
.Y(n_12346)
);

NOR2xp33_ASAP7_75t_L g12347 ( 
.A(n_11333),
.B(n_4925),
.Y(n_12347)
);

AOI21x1_ASAP7_75t_L g12348 ( 
.A1(n_11415),
.A2(n_4930),
.B(n_4927),
.Y(n_12348)
);

NOR2xp33_ASAP7_75t_L g12349 ( 
.A(n_11335),
.B(n_4931),
.Y(n_12349)
);

NOR2xp67_ASAP7_75t_L g12350 ( 
.A(n_11706),
.B(n_4932),
.Y(n_12350)
);

AOI21x1_ASAP7_75t_L g12351 ( 
.A1(n_11431),
.A2(n_11443),
.B(n_11433),
.Y(n_12351)
);

NOR2xp33_ASAP7_75t_L g12352 ( 
.A(n_11741),
.B(n_4933),
.Y(n_12352)
);

INVx4_ASAP7_75t_L g12353 ( 
.A(n_11798),
.Y(n_12353)
);

AOI21xp5_ASAP7_75t_L g12354 ( 
.A1(n_11577),
.A2(n_4936),
.B(n_4934),
.Y(n_12354)
);

OAI21xp5_ASAP7_75t_L g12355 ( 
.A1(n_11306),
.A2(n_451),
.B(n_452),
.Y(n_12355)
);

INVx2_ASAP7_75t_L g12356 ( 
.A(n_11476),
.Y(n_12356)
);

NAND2xp5_ASAP7_75t_L g12357 ( 
.A(n_11490),
.B(n_11505),
.Y(n_12357)
);

OA21x2_ASAP7_75t_L g12358 ( 
.A1(n_11444),
.A2(n_452),
.B(n_453),
.Y(n_12358)
);

AND2x2_ASAP7_75t_L g12359 ( 
.A(n_11904),
.B(n_4937),
.Y(n_12359)
);

AOI21xp5_ASAP7_75t_L g12360 ( 
.A1(n_11643),
.A2(n_4941),
.B(n_4940),
.Y(n_12360)
);

INVx2_ASAP7_75t_SL g12361 ( 
.A(n_11548),
.Y(n_12361)
);

A2O1A1Ixp33_ASAP7_75t_L g12362 ( 
.A1(n_11421),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_12362)
);

AOI21x1_ASAP7_75t_L g12363 ( 
.A1(n_11446),
.A2(n_4943),
.B(n_4942),
.Y(n_12363)
);

NAND3xp33_ASAP7_75t_L g12364 ( 
.A(n_11693),
.B(n_454),
.C(n_455),
.Y(n_12364)
);

NAND2xp5_ASAP7_75t_SL g12365 ( 
.A(n_11324),
.B(n_4944),
.Y(n_12365)
);

A2O1A1Ixp33_ASAP7_75t_L g12366 ( 
.A1(n_11714),
.A2(n_458),
.B(n_456),
.C(n_457),
.Y(n_12366)
);

AND2x4_ASAP7_75t_L g12367 ( 
.A(n_11912),
.B(n_4945),
.Y(n_12367)
);

INVx4_ASAP7_75t_L g12368 ( 
.A(n_11807),
.Y(n_12368)
);

INVx1_ASAP7_75t_L g12369 ( 
.A(n_11448),
.Y(n_12369)
);

AOI21xp5_ASAP7_75t_L g12370 ( 
.A1(n_11683),
.A2(n_4947),
.B(n_4946),
.Y(n_12370)
);

AOI21xp5_ASAP7_75t_L g12371 ( 
.A1(n_11739),
.A2(n_4950),
.B(n_4948),
.Y(n_12371)
);

NAND2xp5_ASAP7_75t_L g12372 ( 
.A(n_11493),
.B(n_457),
.Y(n_12372)
);

AOI21xp5_ASAP7_75t_L g12373 ( 
.A1(n_11452),
.A2(n_11455),
.B(n_11454),
.Y(n_12373)
);

INVx1_ASAP7_75t_L g12374 ( 
.A(n_11460),
.Y(n_12374)
);

INVx2_ASAP7_75t_L g12375 ( 
.A(n_11623),
.Y(n_12375)
);

BUFx8_ASAP7_75t_L g12376 ( 
.A(n_11926),
.Y(n_12376)
);

NAND2xp5_ASAP7_75t_L g12377 ( 
.A(n_11499),
.B(n_11503),
.Y(n_12377)
);

NAND2xp5_ASAP7_75t_L g12378 ( 
.A(n_11506),
.B(n_458),
.Y(n_12378)
);

NAND2xp5_ASAP7_75t_L g12379 ( 
.A(n_11508),
.B(n_459),
.Y(n_12379)
);

INVx8_ASAP7_75t_L g12380 ( 
.A(n_11331),
.Y(n_12380)
);

NAND2xp5_ASAP7_75t_L g12381 ( 
.A(n_11510),
.B(n_459),
.Y(n_12381)
);

AOI21xp5_ASAP7_75t_L g12382 ( 
.A1(n_11464),
.A2(n_4952),
.B(n_4951),
.Y(n_12382)
);

INVx4_ASAP7_75t_L g12383 ( 
.A(n_11812),
.Y(n_12383)
);

AOI22xp33_ASAP7_75t_L g12384 ( 
.A1(n_11372),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_12384)
);

AOI21xp5_ASAP7_75t_L g12385 ( 
.A1(n_11473),
.A2(n_11482),
.B(n_11478),
.Y(n_12385)
);

NAND2xp5_ASAP7_75t_L g12386 ( 
.A(n_11511),
.B(n_461),
.Y(n_12386)
);

O2A1O1Ixp5_ASAP7_75t_L g12387 ( 
.A1(n_11672),
.A2(n_464),
.B(n_462),
.C(n_463),
.Y(n_12387)
);

HB1xp67_ASAP7_75t_L g12388 ( 
.A(n_11515),
.Y(n_12388)
);

INVx1_ASAP7_75t_L g12389 ( 
.A(n_11516),
.Y(n_12389)
);

AOI21xp5_ASAP7_75t_L g12390 ( 
.A1(n_11487),
.A2(n_11349),
.B(n_11520),
.Y(n_12390)
);

AND2x4_ASAP7_75t_L g12391 ( 
.A(n_11655),
.B(n_4953),
.Y(n_12391)
);

OAI21xp33_ASAP7_75t_L g12392 ( 
.A1(n_11825),
.A2(n_11605),
.B(n_11644),
.Y(n_12392)
);

AND2x2_ASAP7_75t_L g12393 ( 
.A(n_11681),
.B(n_4954),
.Y(n_12393)
);

OAI21xp5_ASAP7_75t_L g12394 ( 
.A1(n_11635),
.A2(n_464),
.B(n_465),
.Y(n_12394)
);

O2A1O1Ixp33_ASAP7_75t_L g12395 ( 
.A1(n_11658),
.A2(n_467),
.B(n_465),
.C(n_466),
.Y(n_12395)
);

CKINVDCx5p33_ASAP7_75t_R g12396 ( 
.A(n_11801),
.Y(n_12396)
);

AOI21xp5_ASAP7_75t_L g12397 ( 
.A1(n_11524),
.A2(n_11528),
.B(n_11527),
.Y(n_12397)
);

INVx1_ASAP7_75t_L g12398 ( 
.A(n_11531),
.Y(n_12398)
);

AOI22xp5_ASAP7_75t_L g12399 ( 
.A1(n_11919),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_12399)
);

INVx1_ASAP7_75t_L g12400 ( 
.A(n_11639),
.Y(n_12400)
);

BUFx6f_ASAP7_75t_L g12401 ( 
.A(n_11334),
.Y(n_12401)
);

INVx3_ASAP7_75t_L g12402 ( 
.A(n_11688),
.Y(n_12402)
);

AOI21xp5_ASAP7_75t_L g12403 ( 
.A1(n_11504),
.A2(n_4957),
.B(n_4955),
.Y(n_12403)
);

INVx2_ASAP7_75t_L g12404 ( 
.A(n_11632),
.Y(n_12404)
);

OAI21x1_ASAP7_75t_L g12405 ( 
.A1(n_11733),
.A2(n_4959),
.B(n_4958),
.Y(n_12405)
);

NAND2xp5_ASAP7_75t_SL g12406 ( 
.A(n_11711),
.B(n_4960),
.Y(n_12406)
);

NAND2xp5_ASAP7_75t_L g12407 ( 
.A(n_11544),
.B(n_469),
.Y(n_12407)
);

AND2x2_ASAP7_75t_L g12408 ( 
.A(n_11392),
.B(n_4961),
.Y(n_12408)
);

AOI22xp5_ASAP7_75t_L g12409 ( 
.A1(n_11919),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_12409)
);

NAND3xp33_ASAP7_75t_L g12410 ( 
.A(n_11513),
.B(n_470),
.C(n_471),
.Y(n_12410)
);

AOI21xp33_ASAP7_75t_L g12411 ( 
.A1(n_11325),
.A2(n_472),
.B(n_473),
.Y(n_12411)
);

HB1xp67_ASAP7_75t_L g12412 ( 
.A(n_11675),
.Y(n_12412)
);

AOI22xp5_ASAP7_75t_L g12413 ( 
.A1(n_11600),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_12413)
);

A2O1A1Ixp33_ASAP7_75t_L g12414 ( 
.A1(n_11422),
.A2(n_477),
.B(n_475),
.C(n_476),
.Y(n_12414)
);

NAND2xp5_ASAP7_75t_L g12415 ( 
.A(n_11890),
.B(n_475),
.Y(n_12415)
);

AOI21xp5_ASAP7_75t_L g12416 ( 
.A1(n_11784),
.A2(n_4963),
.B(n_4962),
.Y(n_12416)
);

AOI21xp5_ASAP7_75t_L g12417 ( 
.A1(n_11786),
.A2(n_4965),
.B(n_4964),
.Y(n_12417)
);

NOR2xp33_ASAP7_75t_L g12418 ( 
.A(n_11427),
.B(n_4966),
.Y(n_12418)
);

NOR2x1_ASAP7_75t_R g12419 ( 
.A(n_11374),
.B(n_4969),
.Y(n_12419)
);

AOI21xp5_ASAP7_75t_L g12420 ( 
.A1(n_11797),
.A2(n_4971),
.B(n_4970),
.Y(n_12420)
);

NAND2xp5_ASAP7_75t_L g12421 ( 
.A(n_11682),
.B(n_476),
.Y(n_12421)
);

OAI21x1_ASAP7_75t_L g12422 ( 
.A1(n_11340),
.A2(n_4973),
.B(n_4972),
.Y(n_12422)
);

INVx2_ASAP7_75t_L g12423 ( 
.A(n_11677),
.Y(n_12423)
);

INVx1_ASAP7_75t_L g12424 ( 
.A(n_11498),
.Y(n_12424)
);

O2A1O1Ixp5_ASAP7_75t_L g12425 ( 
.A1(n_11428),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_12425)
);

NAND2xp5_ASAP7_75t_L g12426 ( 
.A(n_11600),
.B(n_478),
.Y(n_12426)
);

BUFx6f_ASAP7_75t_L g12427 ( 
.A(n_11864),
.Y(n_12427)
);

INVx2_ASAP7_75t_L g12428 ( 
.A(n_11730),
.Y(n_12428)
);

NAND2xp5_ASAP7_75t_L g12429 ( 
.A(n_11600),
.B(n_479),
.Y(n_12429)
);

AOI22xp33_ASAP7_75t_L g12430 ( 
.A1(n_11788),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_12430)
);

INVx1_ASAP7_75t_L g12431 ( 
.A(n_11378),
.Y(n_12431)
);

AOI21xp5_ASAP7_75t_L g12432 ( 
.A1(n_11831),
.A2(n_11914),
.B(n_11859),
.Y(n_12432)
);

AOI22xp5_ASAP7_75t_L g12433 ( 
.A1(n_11514),
.A2(n_483),
.B1(n_480),
.B2(n_481),
.Y(n_12433)
);

AND2x2_ASAP7_75t_L g12434 ( 
.A(n_11434),
.B(n_4974),
.Y(n_12434)
);

AOI21x1_ASAP7_75t_L g12435 ( 
.A1(n_11790),
.A2(n_4976),
.B(n_4975),
.Y(n_12435)
);

INVx2_ASAP7_75t_L g12436 ( 
.A(n_11438),
.Y(n_12436)
);

NAND2xp5_ASAP7_75t_SL g12437 ( 
.A(n_11572),
.B(n_4977),
.Y(n_12437)
);

INVx1_ASAP7_75t_L g12438 ( 
.A(n_11491),
.Y(n_12438)
);

AOI21xp5_ASAP7_75t_L g12439 ( 
.A1(n_11916),
.A2(n_4980),
.B(n_4979),
.Y(n_12439)
);

AOI21xp33_ASAP7_75t_L g12440 ( 
.A1(n_11814),
.A2(n_483),
.B(n_484),
.Y(n_12440)
);

OAI21xp5_ASAP7_75t_L g12441 ( 
.A1(n_11536),
.A2(n_484),
.B(n_485),
.Y(n_12441)
);

NAND2xp5_ASAP7_75t_SL g12442 ( 
.A(n_11578),
.B(n_4981),
.Y(n_12442)
);

AOI21xp5_ASAP7_75t_L g12443 ( 
.A1(n_11773),
.A2(n_11450),
.B(n_11398),
.Y(n_12443)
);

AOI21xp5_ASAP7_75t_L g12444 ( 
.A1(n_11381),
.A2(n_4984),
.B(n_4982),
.Y(n_12444)
);

INVx1_ASAP7_75t_L g12445 ( 
.A(n_11702),
.Y(n_12445)
);

NAND2xp5_ASAP7_75t_L g12446 ( 
.A(n_11705),
.B(n_486),
.Y(n_12446)
);

INVx2_ASAP7_75t_L g12447 ( 
.A(n_11468),
.Y(n_12447)
);

NOR2xp33_ASAP7_75t_SL g12448 ( 
.A(n_11802),
.B(n_4986),
.Y(n_12448)
);

INVx11_ASAP7_75t_L g12449 ( 
.A(n_11509),
.Y(n_12449)
);

BUFx12f_ASAP7_75t_L g12450 ( 
.A(n_11362),
.Y(n_12450)
);

INVx2_ASAP7_75t_L g12451 ( 
.A(n_11350),
.Y(n_12451)
);

NAND2xp5_ASAP7_75t_SL g12452 ( 
.A(n_11553),
.B(n_4987),
.Y(n_12452)
);

AO32x2_ASAP7_75t_L g12453 ( 
.A1(n_11827),
.A2(n_488),
.A3(n_486),
.B1(n_487),
.B2(n_489),
.Y(n_12453)
);

AOI22xp5_ASAP7_75t_L g12454 ( 
.A1(n_11731),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_12454)
);

AND2x2_ASAP7_75t_L g12455 ( 
.A(n_11626),
.B(n_4988),
.Y(n_12455)
);

OAI21xp5_ASAP7_75t_L g12456 ( 
.A1(n_11512),
.A2(n_490),
.B(n_491),
.Y(n_12456)
);

NAND2xp5_ASAP7_75t_L g12457 ( 
.A(n_11709),
.B(n_492),
.Y(n_12457)
);

NOR2xp67_ASAP7_75t_SL g12458 ( 
.A(n_11673),
.B(n_492),
.Y(n_12458)
);

AOI21xp5_ASAP7_75t_L g12459 ( 
.A1(n_11557),
.A2(n_4990),
.B(n_4989),
.Y(n_12459)
);

NOR2xp67_ASAP7_75t_L g12460 ( 
.A(n_11767),
.B(n_4991),
.Y(n_12460)
);

OAI22xp5_ASAP7_75t_L g12461 ( 
.A1(n_11465),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_12461)
);

NAND2xp5_ASAP7_75t_L g12462 ( 
.A(n_11674),
.B(n_493),
.Y(n_12462)
);

INVx3_ASAP7_75t_L g12463 ( 
.A(n_11896),
.Y(n_12463)
);

AOI22xp33_ASAP7_75t_L g12464 ( 
.A1(n_11833),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_12464)
);

NAND2xp5_ASAP7_75t_L g12465 ( 
.A(n_11696),
.B(n_496),
.Y(n_12465)
);

A2O1A1Ixp33_ASAP7_75t_L g12466 ( 
.A1(n_11543),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_12466)
);

HB1xp67_ASAP7_75t_L g12467 ( 
.A(n_11609),
.Y(n_12467)
);

AOI21xp5_ASAP7_75t_L g12468 ( 
.A1(n_11457),
.A2(n_4994),
.B(n_4992),
.Y(n_12468)
);

AOI21xp5_ASAP7_75t_L g12469 ( 
.A1(n_11463),
.A2(n_4996),
.B(n_4995),
.Y(n_12469)
);

OAI21xp5_ASAP7_75t_L g12470 ( 
.A1(n_11313),
.A2(n_497),
.B(n_499),
.Y(n_12470)
);

NAND2xp5_ASAP7_75t_L g12471 ( 
.A(n_11517),
.B(n_11472),
.Y(n_12471)
);

INVx1_ASAP7_75t_L g12472 ( 
.A(n_11834),
.Y(n_12472)
);

AOI21xp5_ASAP7_75t_L g12473 ( 
.A1(n_11611),
.A2(n_4998),
.B(n_4997),
.Y(n_12473)
);

NOR2xp67_ASAP7_75t_L g12474 ( 
.A(n_11502),
.B(n_4999),
.Y(n_12474)
);

INVx2_ASAP7_75t_L g12475 ( 
.A(n_11700),
.Y(n_12475)
);

AOI21xp5_ASAP7_75t_L g12476 ( 
.A1(n_11414),
.A2(n_5001),
.B(n_5000),
.Y(n_12476)
);

NAND2x1_ASAP7_75t_L g12477 ( 
.A(n_11497),
.B(n_5002),
.Y(n_12477)
);

NAND2xp5_ASAP7_75t_SL g12478 ( 
.A(n_11521),
.B(n_5003),
.Y(n_12478)
);

AND2x2_ASAP7_75t_L g12479 ( 
.A(n_11634),
.B(n_5004),
.Y(n_12479)
);

NOR2xp33_ASAP7_75t_L g12480 ( 
.A(n_11669),
.B(n_5005),
.Y(n_12480)
);

INVxp67_ASAP7_75t_L g12481 ( 
.A(n_11539),
.Y(n_12481)
);

INVx1_ASAP7_75t_SL g12482 ( 
.A(n_11665),
.Y(n_12482)
);

OAI21xp5_ASAP7_75t_L g12483 ( 
.A1(n_11399),
.A2(n_500),
.B(n_501),
.Y(n_12483)
);

AOI21xp5_ASAP7_75t_L g12484 ( 
.A1(n_11627),
.A2(n_5007),
.B(n_5006),
.Y(n_12484)
);

OAI22xp5_ASAP7_75t_L g12485 ( 
.A1(n_11757),
.A2(n_503),
.B1(n_500),
.B2(n_502),
.Y(n_12485)
);

AOI21xp5_ASAP7_75t_L g12486 ( 
.A1(n_11660),
.A2(n_5009),
.B(n_5008),
.Y(n_12486)
);

AOI22xp5_ASAP7_75t_L g12487 ( 
.A1(n_11401),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_12487)
);

NAND2xp5_ASAP7_75t_SL g12488 ( 
.A(n_11762),
.B(n_5010),
.Y(n_12488)
);

AOI21xp5_ASAP7_75t_L g12489 ( 
.A1(n_11664),
.A2(n_5012),
.B(n_5011),
.Y(n_12489)
);

CKINVDCx10_ASAP7_75t_R g12490 ( 
.A(n_11430),
.Y(n_12490)
);

OAI22xp5_ASAP7_75t_L g12491 ( 
.A1(n_11866),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_12491)
);

AOI21xp5_ASAP7_75t_L g12492 ( 
.A1(n_11909),
.A2(n_5014),
.B(n_5013),
.Y(n_12492)
);

AOI21x1_ASAP7_75t_L g12493 ( 
.A1(n_11871),
.A2(n_5016),
.B(n_5015),
.Y(n_12493)
);

NAND3xp33_ASAP7_75t_SL g12494 ( 
.A(n_11887),
.B(n_505),
.C(n_506),
.Y(n_12494)
);

NOR3xp33_ASAP7_75t_L g12495 ( 
.A(n_11888),
.B(n_11905),
.C(n_11902),
.Y(n_12495)
);

AOI21xp5_ASAP7_75t_L g12496 ( 
.A1(n_11719),
.A2(n_5020),
.B(n_5018),
.Y(n_12496)
);

INVx3_ASAP7_75t_L g12497 ( 
.A(n_11721),
.Y(n_12497)
);

AOI21x1_ASAP7_75t_L g12498 ( 
.A1(n_11618),
.A2(n_5023),
.B(n_5022),
.Y(n_12498)
);

O2A1O1Ixp33_ASAP7_75t_L g12499 ( 
.A1(n_11920),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_12499)
);

AOI21xp5_ASAP7_75t_L g12500 ( 
.A1(n_11293),
.A2(n_5025),
.B(n_5024),
.Y(n_12500)
);

A2O1A1Ixp33_ASAP7_75t_L g12501 ( 
.A1(n_11293),
.A2(n_510),
.B(n_507),
.C(n_508),
.Y(n_12501)
);

INVx2_ASAP7_75t_L g12502 ( 
.A(n_11311),
.Y(n_12502)
);

INVx2_ASAP7_75t_L g12503 ( 
.A(n_11311),
.Y(n_12503)
);

AOI21xp5_ASAP7_75t_L g12504 ( 
.A1(n_11293),
.A2(n_5027),
.B(n_5026),
.Y(n_12504)
);

NOR2xp67_ASAP7_75t_L g12505 ( 
.A(n_11288),
.B(n_5028),
.Y(n_12505)
);

O2A1O1Ixp33_ASAP7_75t_L g12506 ( 
.A1(n_11920),
.A2(n_512),
.B(n_510),
.C(n_511),
.Y(n_12506)
);

INVx11_ASAP7_75t_L g12507 ( 
.A(n_11336),
.Y(n_12507)
);

INVx1_ASAP7_75t_L g12508 ( 
.A(n_11355),
.Y(n_12508)
);

NAND2xp5_ASAP7_75t_L g12509 ( 
.A(n_11338),
.B(n_511),
.Y(n_12509)
);

AOI21xp5_ASAP7_75t_L g12510 ( 
.A1(n_11293),
.A2(n_5030),
.B(n_5029),
.Y(n_12510)
);

NAND2xp5_ASAP7_75t_L g12511 ( 
.A(n_11338),
.B(n_512),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_11355),
.Y(n_12512)
);

O2A1O1Ixp33_ASAP7_75t_SL g12513 ( 
.A1(n_11507),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_12513)
);

AOI21xp5_ASAP7_75t_L g12514 ( 
.A1(n_11293),
.A2(n_5032),
.B(n_5031),
.Y(n_12514)
);

NAND2xp5_ASAP7_75t_L g12515 ( 
.A(n_11338),
.B(n_513),
.Y(n_12515)
);

INVx2_ASAP7_75t_L g12516 ( 
.A(n_11311),
.Y(n_12516)
);

O2A1O1Ixp33_ASAP7_75t_L g12517 ( 
.A1(n_11920),
.A2(n_516),
.B(n_514),
.C(n_515),
.Y(n_12517)
);

AOI21xp5_ASAP7_75t_L g12518 ( 
.A1(n_11293),
.A2(n_5035),
.B(n_5033),
.Y(n_12518)
);

BUFx3_ASAP7_75t_L g12519 ( 
.A(n_11523),
.Y(n_12519)
);

INVx2_ASAP7_75t_L g12520 ( 
.A(n_11311),
.Y(n_12520)
);

INVx3_ASAP7_75t_L g12521 ( 
.A(n_11316),
.Y(n_12521)
);

AOI21xp5_ASAP7_75t_L g12522 ( 
.A1(n_11293),
.A2(n_5037),
.B(n_5036),
.Y(n_12522)
);

A2O1A1Ixp33_ASAP7_75t_L g12523 ( 
.A1(n_11293),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_12523)
);

NOR2xp67_ASAP7_75t_SL g12524 ( 
.A(n_11416),
.B(n_518),
.Y(n_12524)
);

AND2x2_ASAP7_75t_L g12525 ( 
.A(n_11598),
.B(n_5038),
.Y(n_12525)
);

INVx2_ASAP7_75t_L g12526 ( 
.A(n_11311),
.Y(n_12526)
);

AO21x1_ASAP7_75t_L g12527 ( 
.A1(n_11920),
.A2(n_519),
.B(n_520),
.Y(n_12527)
);

OAI21xp33_ASAP7_75t_L g12528 ( 
.A1(n_11293),
.A2(n_521),
.B(n_522),
.Y(n_12528)
);

INVx1_ASAP7_75t_L g12529 ( 
.A(n_11355),
.Y(n_12529)
);

O2A1O1Ixp33_ASAP7_75t_L g12530 ( 
.A1(n_11920),
.A2(n_523),
.B(n_521),
.C(n_522),
.Y(n_12530)
);

INVx2_ASAP7_75t_L g12531 ( 
.A(n_11311),
.Y(n_12531)
);

A2O1A1Ixp33_ASAP7_75t_L g12532 ( 
.A1(n_11293),
.A2(n_525),
.B(n_523),
.C(n_524),
.Y(n_12532)
);

O2A1O1Ixp5_ASAP7_75t_L g12533 ( 
.A1(n_11529),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_12533)
);

INVx4_ASAP7_75t_L g12534 ( 
.A(n_11385),
.Y(n_12534)
);

O2A1O1Ixp33_ASAP7_75t_SL g12535 ( 
.A1(n_11507),
.A2(n_528),
.B(n_526),
.C(n_527),
.Y(n_12535)
);

INVx2_ASAP7_75t_L g12536 ( 
.A(n_11311),
.Y(n_12536)
);

OAI21xp5_ASAP7_75t_L g12537 ( 
.A1(n_11293),
.A2(n_527),
.B(n_528),
.Y(n_12537)
);

AOI21xp5_ASAP7_75t_L g12538 ( 
.A1(n_11293),
.A2(n_5040),
.B(n_5039),
.Y(n_12538)
);

OAI321xp33_ASAP7_75t_L g12539 ( 
.A1(n_11293),
.A2(n_532),
.A3(n_534),
.B1(n_530),
.B2(n_531),
.C(n_533),
.Y(n_12539)
);

AOI21xp5_ASAP7_75t_L g12540 ( 
.A1(n_11293),
.A2(n_5042),
.B(n_5041),
.Y(n_12540)
);

INVxp67_ASAP7_75t_L g12541 ( 
.A(n_11838),
.Y(n_12541)
);

O2A1O1Ixp5_ASAP7_75t_L g12542 ( 
.A1(n_11529),
.A2(n_532),
.B(n_530),
.C(n_531),
.Y(n_12542)
);

INVx2_ASAP7_75t_L g12543 ( 
.A(n_11311),
.Y(n_12543)
);

AO21x1_ASAP7_75t_L g12544 ( 
.A1(n_11920),
.A2(n_533),
.B(n_535),
.Y(n_12544)
);

NAND2xp5_ASAP7_75t_L g12545 ( 
.A(n_11338),
.B(n_535),
.Y(n_12545)
);

NAND2xp5_ASAP7_75t_SL g12546 ( 
.A(n_11293),
.B(n_5044),
.Y(n_12546)
);

A2O1A1Ixp33_ASAP7_75t_L g12547 ( 
.A1(n_11293),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_12547)
);

INVx1_ASAP7_75t_SL g12548 ( 
.A(n_11907),
.Y(n_12548)
);

O2A1O1Ixp33_ASAP7_75t_L g12549 ( 
.A1(n_11920),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_12549)
);

INVx2_ASAP7_75t_L g12550 ( 
.A(n_11311),
.Y(n_12550)
);

INVxp67_ASAP7_75t_SL g12551 ( 
.A(n_11551),
.Y(n_12551)
);

NOR2xp33_ASAP7_75t_L g12552 ( 
.A(n_11293),
.B(n_5045),
.Y(n_12552)
);

O2A1O1Ixp33_ASAP7_75t_L g12553 ( 
.A1(n_11920),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_12553)
);

NAND2xp5_ASAP7_75t_SL g12554 ( 
.A(n_11293),
.B(n_5046),
.Y(n_12554)
);

A2O1A1Ixp33_ASAP7_75t_L g12555 ( 
.A1(n_11293),
.A2(n_542),
.B(n_539),
.C(n_540),
.Y(n_12555)
);

O2A1O1Ixp33_ASAP7_75t_L g12556 ( 
.A1(n_11920),
.A2(n_544),
.B(n_542),
.C(n_543),
.Y(n_12556)
);

NAND2xp5_ASAP7_75t_L g12557 ( 
.A(n_11338),
.B(n_543),
.Y(n_12557)
);

BUFx12f_ASAP7_75t_L g12558 ( 
.A(n_11323),
.Y(n_12558)
);

AOI21xp5_ASAP7_75t_L g12559 ( 
.A1(n_11293),
.A2(n_5048),
.B(n_5047),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_11338),
.B(n_544),
.Y(n_12560)
);

NOR3xp33_ASAP7_75t_L g12561 ( 
.A(n_11416),
.B(n_545),
.C(n_546),
.Y(n_12561)
);

NAND2xp5_ASAP7_75t_L g12562 ( 
.A(n_11338),
.B(n_545),
.Y(n_12562)
);

AOI22xp33_ASAP7_75t_L g12563 ( 
.A1(n_11920),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_12563)
);

NAND2xp5_ASAP7_75t_L g12564 ( 
.A(n_11338),
.B(n_547),
.Y(n_12564)
);

AOI21xp5_ASAP7_75t_L g12565 ( 
.A1(n_11293),
.A2(n_5050),
.B(n_5049),
.Y(n_12565)
);

NAND2xp5_ASAP7_75t_L g12566 ( 
.A(n_11338),
.B(n_549),
.Y(n_12566)
);

NAND2xp5_ASAP7_75t_L g12567 ( 
.A(n_11338),
.B(n_549),
.Y(n_12567)
);

AOI211xp5_ASAP7_75t_L g12568 ( 
.A1(n_11920),
.A2(n_552),
.B(n_550),
.C(n_551),
.Y(n_12568)
);

INVx2_ASAP7_75t_L g12569 ( 
.A(n_11311),
.Y(n_12569)
);

NAND2xp5_ASAP7_75t_L g12570 ( 
.A(n_11338),
.B(n_550),
.Y(n_12570)
);

AOI21xp5_ASAP7_75t_L g12571 ( 
.A1(n_11293),
.A2(n_5052),
.B(n_5051),
.Y(n_12571)
);

INVx3_ASAP7_75t_L g12572 ( 
.A(n_11316),
.Y(n_12572)
);

NAND2xp5_ASAP7_75t_L g12573 ( 
.A(n_11338),
.B(n_551),
.Y(n_12573)
);

INVx2_ASAP7_75t_L g12574 ( 
.A(n_11311),
.Y(n_12574)
);

NAND2xp5_ASAP7_75t_L g12575 ( 
.A(n_11338),
.B(n_552),
.Y(n_12575)
);

O2A1O1Ixp33_ASAP7_75t_L g12576 ( 
.A1(n_11920),
.A2(n_555),
.B(n_553),
.C(n_554),
.Y(n_12576)
);

INVx2_ASAP7_75t_L g12577 ( 
.A(n_11311),
.Y(n_12577)
);

INVx1_ASAP7_75t_L g12578 ( 
.A(n_11355),
.Y(n_12578)
);

OAI321xp33_ASAP7_75t_L g12579 ( 
.A1(n_11293),
.A2(n_555),
.A3(n_557),
.B1(n_553),
.B2(n_554),
.C(n_556),
.Y(n_12579)
);

AOI21xp5_ASAP7_75t_L g12580 ( 
.A1(n_11293),
.A2(n_5054),
.B(n_5053),
.Y(n_12580)
);

OAI21xp5_ASAP7_75t_L g12581 ( 
.A1(n_11293),
.A2(n_556),
.B(n_557),
.Y(n_12581)
);

NOR2xp33_ASAP7_75t_L g12582 ( 
.A(n_11293),
.B(n_5055),
.Y(n_12582)
);

AOI21xp5_ASAP7_75t_L g12583 ( 
.A1(n_11293),
.A2(n_5058),
.B(n_5056),
.Y(n_12583)
);

AOI22xp5_ASAP7_75t_L g12584 ( 
.A1(n_11293),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_12584)
);

AOI21xp5_ASAP7_75t_L g12585 ( 
.A1(n_11293),
.A2(n_5060),
.B(n_5059),
.Y(n_12585)
);

AOI21xp5_ASAP7_75t_L g12586 ( 
.A1(n_11293),
.A2(n_5062),
.B(n_5061),
.Y(n_12586)
);

AOI21xp33_ASAP7_75t_L g12587 ( 
.A1(n_11293),
.A2(n_558),
.B(n_559),
.Y(n_12587)
);

NAND2xp5_ASAP7_75t_L g12588 ( 
.A(n_11338),
.B(n_561),
.Y(n_12588)
);

BUFx6f_ASAP7_75t_L g12589 ( 
.A(n_11541),
.Y(n_12589)
);

AOI22xp33_ASAP7_75t_L g12590 ( 
.A1(n_11920),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_12590)
);

AOI21xp5_ASAP7_75t_L g12591 ( 
.A1(n_11293),
.A2(n_5064),
.B(n_5063),
.Y(n_12591)
);

OAI22xp5_ASAP7_75t_L g12592 ( 
.A1(n_11293),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_12592)
);

NAND2xp5_ASAP7_75t_L g12593 ( 
.A(n_11338),
.B(n_564),
.Y(n_12593)
);

A2O1A1Ixp33_ASAP7_75t_L g12594 ( 
.A1(n_11293),
.A2(n_567),
.B(n_565),
.C(n_566),
.Y(n_12594)
);

INVx2_ASAP7_75t_SL g12595 ( 
.A(n_11614),
.Y(n_12595)
);

AND2x4_ASAP7_75t_L g12596 ( 
.A(n_11407),
.B(n_5065),
.Y(n_12596)
);

CKINVDCx10_ASAP7_75t_R g12597 ( 
.A(n_11822),
.Y(n_12597)
);

NAND2xp5_ASAP7_75t_SL g12598 ( 
.A(n_11293),
.B(n_5066),
.Y(n_12598)
);

NAND2xp5_ASAP7_75t_L g12599 ( 
.A(n_11338),
.B(n_566),
.Y(n_12599)
);

INVx3_ASAP7_75t_SL g12600 ( 
.A(n_11765),
.Y(n_12600)
);

OAI21xp5_ASAP7_75t_L g12601 ( 
.A1(n_11293),
.A2(n_567),
.B(n_568),
.Y(n_12601)
);

AOI21xp5_ASAP7_75t_L g12602 ( 
.A1(n_11293),
.A2(n_5068),
.B(n_5067),
.Y(n_12602)
);

NAND2xp5_ASAP7_75t_L g12603 ( 
.A(n_11338),
.B(n_568),
.Y(n_12603)
);

NAND2xp5_ASAP7_75t_L g12604 ( 
.A(n_11338),
.B(n_569),
.Y(n_12604)
);

A2O1A1Ixp33_ASAP7_75t_L g12605 ( 
.A1(n_11293),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_12605)
);

OAI22xp5_ASAP7_75t_L g12606 ( 
.A1(n_11293),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_12606)
);

NAND2xp5_ASAP7_75t_L g12607 ( 
.A(n_11338),
.B(n_573),
.Y(n_12607)
);

AND2x2_ASAP7_75t_L g12608 ( 
.A(n_11598),
.B(n_5069),
.Y(n_12608)
);

NAND2xp5_ASAP7_75t_L g12609 ( 
.A(n_11338),
.B(n_573),
.Y(n_12609)
);

NOR2xp33_ASAP7_75t_L g12610 ( 
.A(n_11293),
.B(n_5070),
.Y(n_12610)
);

AOI22xp33_ASAP7_75t_L g12611 ( 
.A1(n_11920),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_12611)
);

O2A1O1Ixp33_ASAP7_75t_L g12612 ( 
.A1(n_11920),
.A2(n_577),
.B(n_574),
.C(n_576),
.Y(n_12612)
);

AND2x4_ASAP7_75t_L g12613 ( 
.A(n_11407),
.B(n_5071),
.Y(n_12613)
);

INVx2_ASAP7_75t_L g12614 ( 
.A(n_11311),
.Y(n_12614)
);

AOI21xp5_ASAP7_75t_L g12615 ( 
.A1(n_11293),
.A2(n_5074),
.B(n_5073),
.Y(n_12615)
);

CKINVDCx8_ASAP7_75t_R g12616 ( 
.A(n_11559),
.Y(n_12616)
);

NAND2xp5_ASAP7_75t_L g12617 ( 
.A(n_11338),
.B(n_577),
.Y(n_12617)
);

NAND2xp5_ASAP7_75t_L g12618 ( 
.A(n_11338),
.B(n_578),
.Y(n_12618)
);

AND2x2_ASAP7_75t_L g12619 ( 
.A(n_11598),
.B(n_5076),
.Y(n_12619)
);

INVx1_ASAP7_75t_L g12620 ( 
.A(n_11355),
.Y(n_12620)
);

BUFx6f_ASAP7_75t_L g12621 ( 
.A(n_11541),
.Y(n_12621)
);

CKINVDCx5p33_ASAP7_75t_R g12622 ( 
.A(n_11342),
.Y(n_12622)
);

OAI22xp5_ASAP7_75t_L g12623 ( 
.A1(n_11293),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_12623)
);

OAI21xp33_ASAP7_75t_L g12624 ( 
.A1(n_11293),
.A2(n_579),
.B(n_580),
.Y(n_12624)
);

NAND2xp5_ASAP7_75t_L g12625 ( 
.A(n_11338),
.B(n_581),
.Y(n_12625)
);

NOR2x1_ASAP7_75t_L g12626 ( 
.A(n_11870),
.B(n_581),
.Y(n_12626)
);

INVx2_ASAP7_75t_L g12627 ( 
.A(n_11311),
.Y(n_12627)
);

AOI21xp5_ASAP7_75t_L g12628 ( 
.A1(n_11293),
.A2(n_5078),
.B(n_5077),
.Y(n_12628)
);

NAND2xp5_ASAP7_75t_L g12629 ( 
.A(n_11338),
.B(n_582),
.Y(n_12629)
);

OAI21xp5_ASAP7_75t_L g12630 ( 
.A1(n_11293),
.A2(n_582),
.B(n_583),
.Y(n_12630)
);

INVx3_ASAP7_75t_L g12631 ( 
.A(n_11316),
.Y(n_12631)
);

BUFx4f_ASAP7_75t_SL g12632 ( 
.A(n_11908),
.Y(n_12632)
);

NAND2xp5_ASAP7_75t_L g12633 ( 
.A(n_11338),
.B(n_583),
.Y(n_12633)
);

OAI21x1_ASAP7_75t_L g12634 ( 
.A1(n_11549),
.A2(n_5080),
.B(n_5079),
.Y(n_12634)
);

AND2x2_ASAP7_75t_L g12635 ( 
.A(n_11598),
.B(n_5081),
.Y(n_12635)
);

NOR2x1p5_ASAP7_75t_SL g12636 ( 
.A(n_11549),
.B(n_5082),
.Y(n_12636)
);

NAND2xp5_ASAP7_75t_L g12637 ( 
.A(n_11338),
.B(n_584),
.Y(n_12637)
);

BUFx2_ASAP7_75t_L g12638 ( 
.A(n_11838),
.Y(n_12638)
);

AOI21xp5_ASAP7_75t_L g12639 ( 
.A1(n_11293),
.A2(n_5084),
.B(n_5083),
.Y(n_12639)
);

AND2x2_ASAP7_75t_L g12640 ( 
.A(n_11598),
.B(n_5085),
.Y(n_12640)
);

AOI22xp33_ASAP7_75t_L g12641 ( 
.A1(n_11920),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.Y(n_12641)
);

AND2x2_ASAP7_75t_L g12642 ( 
.A(n_11598),
.B(n_5088),
.Y(n_12642)
);

NAND2xp5_ASAP7_75t_L g12643 ( 
.A(n_11338),
.B(n_585),
.Y(n_12643)
);

INVx3_ASAP7_75t_L g12644 ( 
.A(n_11316),
.Y(n_12644)
);

O2A1O1Ixp33_ASAP7_75t_L g12645 ( 
.A1(n_11920),
.A2(n_589),
.B(n_587),
.C(n_588),
.Y(n_12645)
);

O2A1O1Ixp33_ASAP7_75t_L g12646 ( 
.A1(n_11920),
.A2(n_590),
.B(n_587),
.C(n_588),
.Y(n_12646)
);

INVx2_ASAP7_75t_L g12647 ( 
.A(n_11311),
.Y(n_12647)
);

OR2x6_ASAP7_75t_SL g12648 ( 
.A(n_11374),
.B(n_590),
.Y(n_12648)
);

BUFx6f_ASAP7_75t_L g12649 ( 
.A(n_11541),
.Y(n_12649)
);

A2O1A1Ixp33_ASAP7_75t_L g12650 ( 
.A1(n_11293),
.A2(n_594),
.B(n_591),
.C(n_592),
.Y(n_12650)
);

NAND2xp5_ASAP7_75t_L g12651 ( 
.A(n_11338),
.B(n_592),
.Y(n_12651)
);

AND2x2_ASAP7_75t_L g12652 ( 
.A(n_11598),
.B(n_5089),
.Y(n_12652)
);

AOI21xp5_ASAP7_75t_L g12653 ( 
.A1(n_11293),
.A2(n_5092),
.B(n_5090),
.Y(n_12653)
);

O2A1O1Ixp33_ASAP7_75t_L g12654 ( 
.A1(n_11920),
.A2(n_596),
.B(n_594),
.C(n_595),
.Y(n_12654)
);

INVx1_ASAP7_75t_L g12655 ( 
.A(n_11355),
.Y(n_12655)
);

AND2x4_ASAP7_75t_L g12656 ( 
.A(n_11407),
.B(n_5093),
.Y(n_12656)
);

INVx2_ASAP7_75t_L g12657 ( 
.A(n_11311),
.Y(n_12657)
);

AOI21xp5_ASAP7_75t_L g12658 ( 
.A1(n_11293),
.A2(n_5095),
.B(n_5094),
.Y(n_12658)
);

AOI21xp5_ASAP7_75t_L g12659 ( 
.A1(n_11293),
.A2(n_5097),
.B(n_5096),
.Y(n_12659)
);

AOI21x1_ASAP7_75t_L g12660 ( 
.A1(n_11339),
.A2(n_5099),
.B(n_5098),
.Y(n_12660)
);

NAND2xp5_ASAP7_75t_L g12661 ( 
.A(n_11338),
.B(n_597),
.Y(n_12661)
);

AOI21xp5_ASAP7_75t_L g12662 ( 
.A1(n_11293),
.A2(n_5101),
.B(n_5100),
.Y(n_12662)
);

INVxp67_ASAP7_75t_L g12663 ( 
.A(n_11838),
.Y(n_12663)
);

AOI22xp5_ASAP7_75t_L g12664 ( 
.A1(n_11293),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_12664)
);

NAND2xp5_ASAP7_75t_SL g12665 ( 
.A(n_11293),
.B(n_5102),
.Y(n_12665)
);

NAND2xp5_ASAP7_75t_L g12666 ( 
.A(n_11338),
.B(n_598),
.Y(n_12666)
);

INVx1_ASAP7_75t_L g12667 ( 
.A(n_11355),
.Y(n_12667)
);

AOI21xp5_ASAP7_75t_L g12668 ( 
.A1(n_11293),
.A2(n_5105),
.B(n_5104),
.Y(n_12668)
);

AOI21xp5_ASAP7_75t_L g12669 ( 
.A1(n_11293),
.A2(n_5108),
.B(n_5107),
.Y(n_12669)
);

AOI21xp5_ASAP7_75t_L g12670 ( 
.A1(n_11293),
.A2(n_5110),
.B(n_5109),
.Y(n_12670)
);

NAND2xp5_ASAP7_75t_L g12671 ( 
.A(n_11338),
.B(n_599),
.Y(n_12671)
);

NAND2xp5_ASAP7_75t_SL g12672 ( 
.A(n_11293),
.B(n_5111),
.Y(n_12672)
);

NAND2xp5_ASAP7_75t_SL g12673 ( 
.A(n_11293),
.B(n_5112),
.Y(n_12673)
);

AOI22xp5_ASAP7_75t_L g12674 ( 
.A1(n_11293),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_12674)
);

NAND2xp5_ASAP7_75t_L g12675 ( 
.A(n_11338),
.B(n_600),
.Y(n_12675)
);

NAND2xp5_ASAP7_75t_SL g12676 ( 
.A(n_11293),
.B(n_5113),
.Y(n_12676)
);

AOI21xp5_ASAP7_75t_L g12677 ( 
.A1(n_11293),
.A2(n_5115),
.B(n_5114),
.Y(n_12677)
);

NAND2x1_ASAP7_75t_L g12678 ( 
.A(n_11752),
.B(n_5116),
.Y(n_12678)
);

AO21x1_ASAP7_75t_L g12679 ( 
.A1(n_11920),
.A2(n_601),
.B(n_602),
.Y(n_12679)
);

BUFx6f_ASAP7_75t_L g12680 ( 
.A(n_11541),
.Y(n_12680)
);

INVx3_ASAP7_75t_L g12681 ( 
.A(n_11316),
.Y(n_12681)
);

NAND2xp5_ASAP7_75t_L g12682 ( 
.A(n_11338),
.B(n_603),
.Y(n_12682)
);

AOI21xp5_ASAP7_75t_L g12683 ( 
.A1(n_11293),
.A2(n_5118),
.B(n_5117),
.Y(n_12683)
);

A2O1A1Ixp33_ASAP7_75t_L g12684 ( 
.A1(n_11293),
.A2(n_605),
.B(n_603),
.C(n_604),
.Y(n_12684)
);

AOI21xp5_ASAP7_75t_L g12685 ( 
.A1(n_11293),
.A2(n_5120),
.B(n_5119),
.Y(n_12685)
);

INVx2_ASAP7_75t_L g12686 ( 
.A(n_11311),
.Y(n_12686)
);

INVx1_ASAP7_75t_L g12687 ( 
.A(n_11355),
.Y(n_12687)
);

AOI21x1_ASAP7_75t_L g12688 ( 
.A1(n_11339),
.A2(n_5123),
.B(n_5122),
.Y(n_12688)
);

OAI22xp5_ASAP7_75t_L g12689 ( 
.A1(n_11293),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_12689)
);

AOI22xp5_ASAP7_75t_L g12690 ( 
.A1(n_11293),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.Y(n_12690)
);

AOI22xp5_ASAP7_75t_L g12691 ( 
.A1(n_11293),
.A2(n_610),
.B1(n_607),
.B2(n_609),
.Y(n_12691)
);

NOR2xp33_ASAP7_75t_L g12692 ( 
.A(n_11293),
.B(n_5125),
.Y(n_12692)
);

AOI21x1_ASAP7_75t_L g12693 ( 
.A1(n_11339),
.A2(n_5128),
.B(n_5126),
.Y(n_12693)
);

AOI22xp5_ASAP7_75t_L g12694 ( 
.A1(n_11293),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_12694)
);

NOR2xp33_ASAP7_75t_L g12695 ( 
.A(n_11293),
.B(n_5129),
.Y(n_12695)
);

OAI22xp5_ASAP7_75t_SL g12696 ( 
.A1(n_11293),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_12696)
);

NOR3xp33_ASAP7_75t_L g12697 ( 
.A(n_11416),
.B(n_612),
.C(n_613),
.Y(n_12697)
);

NAND2xp5_ASAP7_75t_SL g12698 ( 
.A(n_11293),
.B(n_5130),
.Y(n_12698)
);

NOR2xp33_ASAP7_75t_L g12699 ( 
.A(n_11293),
.B(n_5131),
.Y(n_12699)
);

OAI22xp5_ASAP7_75t_L g12700 ( 
.A1(n_11293),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_12700)
);

NAND2xp5_ASAP7_75t_L g12701 ( 
.A(n_11338),
.B(n_616),
.Y(n_12701)
);

AOI21xp5_ASAP7_75t_L g12702 ( 
.A1(n_11293),
.A2(n_5134),
.B(n_5132),
.Y(n_12702)
);

NAND2xp5_ASAP7_75t_L g12703 ( 
.A(n_11338),
.B(n_617),
.Y(n_12703)
);

O2A1O1Ixp33_ASAP7_75t_L g12704 ( 
.A1(n_11920),
.A2(n_620),
.B(n_618),
.C(n_619),
.Y(n_12704)
);

AND2x2_ASAP7_75t_L g12705 ( 
.A(n_11598),
.B(n_5135),
.Y(n_12705)
);

AOI21xp5_ASAP7_75t_L g12706 ( 
.A1(n_11293),
.A2(n_5137),
.B(n_5136),
.Y(n_12706)
);

AOI21xp5_ASAP7_75t_L g12707 ( 
.A1(n_11293),
.A2(n_5139),
.B(n_5138),
.Y(n_12707)
);

NAND2xp5_ASAP7_75t_L g12708 ( 
.A(n_11338),
.B(n_618),
.Y(n_12708)
);

OAI22xp5_ASAP7_75t_L g12709 ( 
.A1(n_11293),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_12709)
);

OAI21xp5_ASAP7_75t_L g12710 ( 
.A1(n_11293),
.A2(n_621),
.B(n_622),
.Y(n_12710)
);

AOI21xp5_ASAP7_75t_L g12711 ( 
.A1(n_11293),
.A2(n_5143),
.B(n_5140),
.Y(n_12711)
);

NAND2xp5_ASAP7_75t_SL g12712 ( 
.A(n_11293),
.B(n_5145),
.Y(n_12712)
);

INVx2_ASAP7_75t_L g12713 ( 
.A(n_11311),
.Y(n_12713)
);

AOI21xp5_ASAP7_75t_L g12714 ( 
.A1(n_11293),
.A2(n_5147),
.B(n_5146),
.Y(n_12714)
);

NOR2x1_ASAP7_75t_L g12715 ( 
.A(n_11870),
.B(n_622),
.Y(n_12715)
);

AOI21xp5_ASAP7_75t_L g12716 ( 
.A1(n_11293),
.A2(n_5149),
.B(n_5148),
.Y(n_12716)
);

INVx3_ASAP7_75t_L g12717 ( 
.A(n_11316),
.Y(n_12717)
);

A2O1A1Ixp33_ASAP7_75t_L g12718 ( 
.A1(n_11293),
.A2(n_625),
.B(n_623),
.C(n_624),
.Y(n_12718)
);

AOI21xp5_ASAP7_75t_L g12719 ( 
.A1(n_11293),
.A2(n_5152),
.B(n_5150),
.Y(n_12719)
);

NOR2xp33_ASAP7_75t_SL g12720 ( 
.A(n_11361),
.B(n_5153),
.Y(n_12720)
);

AOI21x1_ASAP7_75t_L g12721 ( 
.A1(n_11339),
.A2(n_5155),
.B(n_5154),
.Y(n_12721)
);

AOI33xp33_ASAP7_75t_L g12722 ( 
.A1(n_11293),
.A2(n_625),
.A3(n_628),
.B1(n_623),
.B2(n_624),
.B3(n_626),
.Y(n_12722)
);

NAND2xp5_ASAP7_75t_L g12723 ( 
.A(n_11338),
.B(n_626),
.Y(n_12723)
);

AOI21xp5_ASAP7_75t_L g12724 ( 
.A1(n_11293),
.A2(n_5157),
.B(n_5156),
.Y(n_12724)
);

AOI21xp5_ASAP7_75t_L g12725 ( 
.A1(n_11293),
.A2(n_5159),
.B(n_5158),
.Y(n_12725)
);

INVx3_ASAP7_75t_L g12726 ( 
.A(n_11316),
.Y(n_12726)
);

NAND2xp5_ASAP7_75t_SL g12727 ( 
.A(n_11293),
.B(n_5160),
.Y(n_12727)
);

INVx2_ASAP7_75t_SL g12728 ( 
.A(n_11614),
.Y(n_12728)
);

A2O1A1Ixp33_ASAP7_75t_L g12729 ( 
.A1(n_11293),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_12729)
);

NOR2xp33_ASAP7_75t_L g12730 ( 
.A(n_11293),
.B(n_5161),
.Y(n_12730)
);

AO32x2_ASAP7_75t_L g12731 ( 
.A1(n_11529),
.A2(n_631),
.A3(n_629),
.B1(n_630),
.B2(n_632),
.Y(n_12731)
);

OAI321xp33_ASAP7_75t_L g12732 ( 
.A1(n_11293),
.A2(n_634),
.A3(n_636),
.B1(n_631),
.B2(n_633),
.C(n_635),
.Y(n_12732)
);

OR2x4_ASAP7_75t_L g12733 ( 
.A(n_11373),
.B(n_633),
.Y(n_12733)
);

INVx1_ASAP7_75t_L g12734 ( 
.A(n_11355),
.Y(n_12734)
);

NAND2xp5_ASAP7_75t_L g12735 ( 
.A(n_11338),
.B(n_634),
.Y(n_12735)
);

INVx1_ASAP7_75t_L g12736 ( 
.A(n_11355),
.Y(n_12736)
);

AND2x2_ASAP7_75t_L g12737 ( 
.A(n_11598),
.B(n_5162),
.Y(n_12737)
);

OAI21xp5_ASAP7_75t_L g12738 ( 
.A1(n_11293),
.A2(n_635),
.B(n_637),
.Y(n_12738)
);

BUFx6f_ASAP7_75t_L g12739 ( 
.A(n_11541),
.Y(n_12739)
);

AOI22xp5_ASAP7_75t_L g12740 ( 
.A1(n_11293),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.Y(n_12740)
);

AOI21xp5_ASAP7_75t_L g12741 ( 
.A1(n_11293),
.A2(n_5164),
.B(n_5163),
.Y(n_12741)
);

NAND2xp5_ASAP7_75t_SL g12742 ( 
.A(n_11293),
.B(n_5165),
.Y(n_12742)
);

NAND2xp5_ASAP7_75t_L g12743 ( 
.A(n_11338),
.B(n_638),
.Y(n_12743)
);

O2A1O1Ixp33_ASAP7_75t_L g12744 ( 
.A1(n_11920),
.A2(n_641),
.B(n_639),
.C(n_640),
.Y(n_12744)
);

INVx1_ASAP7_75t_L g12745 ( 
.A(n_11355),
.Y(n_12745)
);

NAND2xp5_ASAP7_75t_L g12746 ( 
.A(n_11338),
.B(n_640),
.Y(n_12746)
);

AOI21xp5_ASAP7_75t_L g12747 ( 
.A1(n_11293),
.A2(n_5168),
.B(n_5166),
.Y(n_12747)
);

INVx2_ASAP7_75t_L g12748 ( 
.A(n_11311),
.Y(n_12748)
);

NAND2xp33_ASAP7_75t_L g12749 ( 
.A(n_11293),
.B(n_642),
.Y(n_12749)
);

AOI21xp5_ASAP7_75t_L g12750 ( 
.A1(n_11293),
.A2(n_5170),
.B(n_5169),
.Y(n_12750)
);

NAND2xp5_ASAP7_75t_L g12751 ( 
.A(n_11338),
.B(n_642),
.Y(n_12751)
);

O2A1O1Ixp5_ASAP7_75t_L g12752 ( 
.A1(n_11529),
.A2(n_645),
.B(n_643),
.C(n_644),
.Y(n_12752)
);

NAND2xp5_ASAP7_75t_L g12753 ( 
.A(n_11338),
.B(n_643),
.Y(n_12753)
);

AOI22xp33_ASAP7_75t_L g12754 ( 
.A1(n_11920),
.A2(n_647),
.B1(n_645),
.B2(n_646),
.Y(n_12754)
);

NAND2xp5_ASAP7_75t_L g12755 ( 
.A(n_11338),
.B(n_646),
.Y(n_12755)
);

NAND2xp5_ASAP7_75t_L g12756 ( 
.A(n_11338),
.B(n_647),
.Y(n_12756)
);

AND2x2_ASAP7_75t_L g12757 ( 
.A(n_11598),
.B(n_5171),
.Y(n_12757)
);

NAND2xp5_ASAP7_75t_SL g12758 ( 
.A(n_11293),
.B(n_5172),
.Y(n_12758)
);

O2A1O1Ixp5_ASAP7_75t_L g12759 ( 
.A1(n_11529),
.A2(n_650),
.B(n_648),
.C(n_649),
.Y(n_12759)
);

INVx2_ASAP7_75t_L g12760 ( 
.A(n_11311),
.Y(n_12760)
);

HB1xp67_ASAP7_75t_L g12761 ( 
.A(n_11838),
.Y(n_12761)
);

NAND2xp5_ASAP7_75t_L g12762 ( 
.A(n_11338),
.B(n_648),
.Y(n_12762)
);

NAND2xp5_ASAP7_75t_L g12763 ( 
.A(n_11338),
.B(n_649),
.Y(n_12763)
);

NAND2xp5_ASAP7_75t_L g12764 ( 
.A(n_11338),
.B(n_650),
.Y(n_12764)
);

AND2x2_ASAP7_75t_L g12765 ( 
.A(n_11598),
.B(n_5173),
.Y(n_12765)
);

AOI22xp5_ASAP7_75t_L g12766 ( 
.A1(n_11293),
.A2(n_653),
.B1(n_651),
.B2(n_652),
.Y(n_12766)
);

NAND2xp5_ASAP7_75t_L g12767 ( 
.A(n_11338),
.B(n_651),
.Y(n_12767)
);

AOI21xp5_ASAP7_75t_L g12768 ( 
.A1(n_11293),
.A2(n_5175),
.B(n_5174),
.Y(n_12768)
);

HB1xp67_ASAP7_75t_L g12769 ( 
.A(n_11838),
.Y(n_12769)
);

AOI21xp5_ASAP7_75t_L g12770 ( 
.A1(n_11293),
.A2(n_5177),
.B(n_5176),
.Y(n_12770)
);

INVx2_ASAP7_75t_L g12771 ( 
.A(n_11311),
.Y(n_12771)
);

INVx3_ASAP7_75t_L g12772 ( 
.A(n_11316),
.Y(n_12772)
);

OAI22xp5_ASAP7_75t_L g12773 ( 
.A1(n_11293),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_12773)
);

NAND2xp5_ASAP7_75t_L g12774 ( 
.A(n_11338),
.B(n_654),
.Y(n_12774)
);

NOR2xp67_ASAP7_75t_L g12775 ( 
.A(n_11288),
.B(n_5178),
.Y(n_12775)
);

AOI21xp5_ASAP7_75t_L g12776 ( 
.A1(n_11293),
.A2(n_5180),
.B(n_5179),
.Y(n_12776)
);

OAI21xp5_ASAP7_75t_L g12777 ( 
.A1(n_11293),
.A2(n_655),
.B(n_656),
.Y(n_12777)
);

BUFx3_ASAP7_75t_L g12778 ( 
.A(n_11523),
.Y(n_12778)
);

AOI21xp5_ASAP7_75t_L g12779 ( 
.A1(n_11293),
.A2(n_5184),
.B(n_5181),
.Y(n_12779)
);

NOR2xp33_ASAP7_75t_L g12780 ( 
.A(n_11293),
.B(n_5185),
.Y(n_12780)
);

OAI21xp5_ASAP7_75t_L g12781 ( 
.A1(n_11293),
.A2(n_655),
.B(n_656),
.Y(n_12781)
);

NOR2xp33_ASAP7_75t_L g12782 ( 
.A(n_11293),
.B(n_5186),
.Y(n_12782)
);

AOI21xp5_ASAP7_75t_L g12783 ( 
.A1(n_11293),
.A2(n_5188),
.B(n_5187),
.Y(n_12783)
);

INVx1_ASAP7_75t_SL g12784 ( 
.A(n_11907),
.Y(n_12784)
);

AOI22xp5_ASAP7_75t_L g12785 ( 
.A1(n_11293),
.A2(n_660),
.B1(n_657),
.B2(n_659),
.Y(n_12785)
);

NOR2x1_ASAP7_75t_L g12786 ( 
.A(n_11870),
.B(n_657),
.Y(n_12786)
);

BUFx3_ASAP7_75t_L g12787 ( 
.A(n_11523),
.Y(n_12787)
);

AOI21xp5_ASAP7_75t_L g12788 ( 
.A1(n_11293),
.A2(n_5190),
.B(n_5189),
.Y(n_12788)
);

AND2x2_ASAP7_75t_L g12789 ( 
.A(n_11598),
.B(n_5191),
.Y(n_12789)
);

NOR2xp33_ASAP7_75t_SL g12790 ( 
.A(n_11361),
.B(n_5193),
.Y(n_12790)
);

AOI22xp5_ASAP7_75t_L g12791 ( 
.A1(n_11293),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.Y(n_12791)
);

NAND3xp33_ASAP7_75t_L g12792 ( 
.A(n_12749),
.B(n_662),
.C(n_663),
.Y(n_12792)
);

INVx5_ASAP7_75t_L g12793 ( 
.A(n_11970),
.Y(n_12793)
);

OAI22xp5_ASAP7_75t_L g12794 ( 
.A1(n_12155),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.Y(n_12794)
);

AOI21xp5_ASAP7_75t_L g12795 ( 
.A1(n_11937),
.A2(n_12326),
.B(n_11934),
.Y(n_12795)
);

AOI21xp5_ASAP7_75t_L g12796 ( 
.A1(n_12304),
.A2(n_5196),
.B(n_5195),
.Y(n_12796)
);

BUFx6f_ASAP7_75t_L g12797 ( 
.A(n_11999),
.Y(n_12797)
);

AOI21xp5_ASAP7_75t_L g12798 ( 
.A1(n_12315),
.A2(n_5198),
.B(n_5197),
.Y(n_12798)
);

OAI22xp5_ASAP7_75t_L g12799 ( 
.A1(n_12568),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_12799)
);

NOR2xp33_ASAP7_75t_L g12800 ( 
.A(n_12098),
.B(n_666),
.Y(n_12800)
);

AOI21xp5_ASAP7_75t_L g12801 ( 
.A1(n_11993),
.A2(n_5200),
.B(n_5199),
.Y(n_12801)
);

AOI21xp5_ASAP7_75t_L g12802 ( 
.A1(n_12010),
.A2(n_5202),
.B(n_5201),
.Y(n_12802)
);

O2A1O1Ixp33_ASAP7_75t_L g12803 ( 
.A1(n_11955),
.A2(n_669),
.B(n_667),
.C(n_668),
.Y(n_12803)
);

AND2x4_ASAP7_75t_L g12804 ( 
.A(n_12638),
.B(n_5203),
.Y(n_12804)
);

NOR2x1_ASAP7_75t_L g12805 ( 
.A(n_12049),
.B(n_668),
.Y(n_12805)
);

A2O1A1Ixp33_ASAP7_75t_L g12806 ( 
.A1(n_11952),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_12806)
);

INVx1_ASAP7_75t_L g12807 ( 
.A(n_12185),
.Y(n_12807)
);

INVx1_ASAP7_75t_L g12808 ( 
.A(n_12246),
.Y(n_12808)
);

AOI22xp33_ASAP7_75t_L g12809 ( 
.A1(n_12561),
.A2(n_672),
.B1(n_670),
.B2(n_671),
.Y(n_12809)
);

NAND2xp5_ASAP7_75t_L g12810 ( 
.A(n_12761),
.B(n_672),
.Y(n_12810)
);

CKINVDCx5p33_ASAP7_75t_R g12811 ( 
.A(n_11958),
.Y(n_12811)
);

BUFx12f_ASAP7_75t_L g12812 ( 
.A(n_12396),
.Y(n_12812)
);

NOR2xp33_ASAP7_75t_L g12813 ( 
.A(n_12632),
.B(n_12548),
.Y(n_12813)
);

AOI21xp5_ASAP7_75t_L g12814 ( 
.A1(n_12017),
.A2(n_5206),
.B(n_5204),
.Y(n_12814)
);

NAND2xp5_ASAP7_75t_L g12815 ( 
.A(n_12769),
.B(n_673),
.Y(n_12815)
);

AOI21xp5_ASAP7_75t_L g12816 ( 
.A1(n_12042),
.A2(n_5208),
.B(n_5207),
.Y(n_12816)
);

AOI21xp5_ASAP7_75t_L g12817 ( 
.A1(n_11935),
.A2(n_5212),
.B(n_5211),
.Y(n_12817)
);

NAND2xp5_ASAP7_75t_L g12818 ( 
.A(n_11938),
.B(n_673),
.Y(n_12818)
);

AND2x2_ASAP7_75t_L g12819 ( 
.A(n_12302),
.B(n_674),
.Y(n_12819)
);

O2A1O1Ixp33_ASAP7_75t_L g12820 ( 
.A1(n_11930),
.A2(n_676),
.B(n_674),
.C(n_675),
.Y(n_12820)
);

AOI22xp5_ASAP7_75t_L g12821 ( 
.A1(n_12697),
.A2(n_678),
.B1(n_676),
.B2(n_677),
.Y(n_12821)
);

INVx3_ASAP7_75t_L g12822 ( 
.A(n_12097),
.Y(n_12822)
);

BUFx12f_ASAP7_75t_L g12823 ( 
.A(n_12303),
.Y(n_12823)
);

NAND2xp5_ASAP7_75t_SL g12824 ( 
.A(n_11949),
.B(n_5213),
.Y(n_12824)
);

NOR2xp33_ASAP7_75t_L g12825 ( 
.A(n_12784),
.B(n_677),
.Y(n_12825)
);

NOR2xp33_ASAP7_75t_L g12826 ( 
.A(n_12007),
.B(n_11940),
.Y(n_12826)
);

NAND3xp33_ASAP7_75t_L g12827 ( 
.A(n_12002),
.B(n_678),
.C(n_679),
.Y(n_12827)
);

OAI21xp33_ASAP7_75t_SL g12828 ( 
.A1(n_12327),
.A2(n_679),
.B(n_680),
.Y(n_12828)
);

A2O1A1Ixp33_ASAP7_75t_L g12829 ( 
.A1(n_12088),
.A2(n_682),
.B(n_680),
.C(n_681),
.Y(n_12829)
);

AOI21xp5_ASAP7_75t_L g12830 ( 
.A1(n_12207),
.A2(n_5217),
.B(n_5214),
.Y(n_12830)
);

NAND2xp5_ASAP7_75t_L g12831 ( 
.A(n_12423),
.B(n_682),
.Y(n_12831)
);

AOI21xp5_ASAP7_75t_L g12832 ( 
.A1(n_12044),
.A2(n_5220),
.B(n_5219),
.Y(n_12832)
);

O2A1O1Ixp33_ASAP7_75t_L g12833 ( 
.A1(n_12501),
.A2(n_685),
.B(n_683),
.C(n_684),
.Y(n_12833)
);

INVx2_ASAP7_75t_L g12834 ( 
.A(n_12400),
.Y(n_12834)
);

NAND2xp5_ASAP7_75t_L g12835 ( 
.A(n_12551),
.B(n_683),
.Y(n_12835)
);

AOI22x1_ASAP7_75t_L g12836 ( 
.A1(n_11946),
.A2(n_687),
.B1(n_684),
.B2(n_686),
.Y(n_12836)
);

OAI21xp33_ASAP7_75t_SL g12837 ( 
.A1(n_12722),
.A2(n_686),
.B(n_687),
.Y(n_12837)
);

AOI21xp5_ASAP7_75t_L g12838 ( 
.A1(n_12546),
.A2(n_12598),
.B(n_12554),
.Y(n_12838)
);

AOI21x1_ASAP7_75t_L g12839 ( 
.A1(n_12660),
.A2(n_688),
.B(n_689),
.Y(n_12839)
);

O2A1O1Ixp5_ASAP7_75t_L g12840 ( 
.A1(n_12524),
.A2(n_690),
.B(n_688),
.C(n_689),
.Y(n_12840)
);

NAND2xp5_ASAP7_75t_SL g12841 ( 
.A(n_12012),
.B(n_5223),
.Y(n_12841)
);

INVx2_ASAP7_75t_L g12842 ( 
.A(n_12375),
.Y(n_12842)
);

O2A1O1Ixp5_ASAP7_75t_L g12843 ( 
.A1(n_12527),
.A2(n_692),
.B(n_690),
.C(n_691),
.Y(n_12843)
);

AOI21xp5_ASAP7_75t_L g12844 ( 
.A1(n_12665),
.A2(n_5225),
.B(n_5224),
.Y(n_12844)
);

AOI221xp5_ASAP7_75t_L g12845 ( 
.A1(n_12587),
.A2(n_693),
.B1(n_691),
.B2(n_692),
.C(n_694),
.Y(n_12845)
);

NAND2xp5_ASAP7_75t_L g12846 ( 
.A(n_12541),
.B(n_693),
.Y(n_12846)
);

NAND2xp5_ASAP7_75t_SL g12847 ( 
.A(n_11995),
.B(n_12432),
.Y(n_12847)
);

NAND2xp5_ASAP7_75t_L g12848 ( 
.A(n_12663),
.B(n_695),
.Y(n_12848)
);

NOR2x1_ASAP7_75t_L g12849 ( 
.A(n_12153),
.B(n_696),
.Y(n_12849)
);

OAI22xp5_ASAP7_75t_L g12850 ( 
.A1(n_12563),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.Y(n_12850)
);

OAI22x1_ASAP7_75t_L g12851 ( 
.A1(n_12120),
.A2(n_700),
.B1(n_697),
.B2(n_699),
.Y(n_12851)
);

BUFx2_ASAP7_75t_L g12852 ( 
.A(n_12121),
.Y(n_12852)
);

NAND2xp5_ASAP7_75t_L g12853 ( 
.A(n_12051),
.B(n_700),
.Y(n_12853)
);

INVx1_ASAP7_75t_L g12854 ( 
.A(n_12260),
.Y(n_12854)
);

NAND2xp5_ASAP7_75t_L g12855 ( 
.A(n_12075),
.B(n_701),
.Y(n_12855)
);

AOI21xp5_ASAP7_75t_L g12856 ( 
.A1(n_12672),
.A2(n_5227),
.B(n_5226),
.Y(n_12856)
);

AOI21xp5_ASAP7_75t_L g12857 ( 
.A1(n_12673),
.A2(n_5230),
.B(n_5229),
.Y(n_12857)
);

NAND2xp5_ASAP7_75t_L g12858 ( 
.A(n_11985),
.B(n_701),
.Y(n_12858)
);

INVx2_ASAP7_75t_SL g12859 ( 
.A(n_12167),
.Y(n_12859)
);

OAI22xp5_ASAP7_75t_L g12860 ( 
.A1(n_12590),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_12860)
);

NAND2xp5_ASAP7_75t_L g12861 ( 
.A(n_12113),
.B(n_703),
.Y(n_12861)
);

INVx2_ASAP7_75t_SL g12862 ( 
.A(n_12097),
.Y(n_12862)
);

INVx2_ASAP7_75t_L g12863 ( 
.A(n_11931),
.Y(n_12863)
);

AND2x2_ASAP7_75t_L g12864 ( 
.A(n_12388),
.B(n_704),
.Y(n_12864)
);

OR2x6_ASAP7_75t_L g12865 ( 
.A(n_12159),
.B(n_5231),
.Y(n_12865)
);

AOI21xp5_ASAP7_75t_L g12866 ( 
.A1(n_12676),
.A2(n_5234),
.B(n_5233),
.Y(n_12866)
);

CKINVDCx6p67_ASAP7_75t_R g12867 ( 
.A(n_12597),
.Y(n_12867)
);

AOI21xp5_ASAP7_75t_L g12868 ( 
.A1(n_12698),
.A2(n_5237),
.B(n_5235),
.Y(n_12868)
);

OR2x6_ASAP7_75t_L g12869 ( 
.A(n_11950),
.B(n_5239),
.Y(n_12869)
);

AOI21xp5_ASAP7_75t_L g12870 ( 
.A1(n_12712),
.A2(n_5242),
.B(n_5240),
.Y(n_12870)
);

AOI21xp5_ASAP7_75t_L g12871 ( 
.A1(n_12727),
.A2(n_5244),
.B(n_5243),
.Y(n_12871)
);

AO21x2_ASAP7_75t_L g12872 ( 
.A1(n_11959),
.A2(n_705),
.B(n_706),
.Y(n_12872)
);

AOI22xp33_ASAP7_75t_SL g12873 ( 
.A1(n_12537),
.A2(n_708),
.B1(n_705),
.B2(n_707),
.Y(n_12873)
);

OAI21xp5_ASAP7_75t_L g12874 ( 
.A1(n_12552),
.A2(n_5247),
.B(n_5245),
.Y(n_12874)
);

AOI21xp5_ASAP7_75t_L g12875 ( 
.A1(n_12742),
.A2(n_5250),
.B(n_5248),
.Y(n_12875)
);

INVx1_ASAP7_75t_L g12876 ( 
.A(n_12351),
.Y(n_12876)
);

NAND2xp5_ASAP7_75t_L g12877 ( 
.A(n_12030),
.B(n_707),
.Y(n_12877)
);

AOI21xp5_ASAP7_75t_L g12878 ( 
.A1(n_12758),
.A2(n_5252),
.B(n_5251),
.Y(n_12878)
);

AOI21xp5_ASAP7_75t_L g12879 ( 
.A1(n_12499),
.A2(n_5254),
.B(n_5253),
.Y(n_12879)
);

NAND2xp5_ASAP7_75t_L g12880 ( 
.A(n_11953),
.B(n_708),
.Y(n_12880)
);

INVx2_ASAP7_75t_L g12881 ( 
.A(n_11933),
.Y(n_12881)
);

AOI22xp5_ASAP7_75t_L g12882 ( 
.A1(n_12016),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.Y(n_12882)
);

NAND2xp5_ASAP7_75t_L g12883 ( 
.A(n_11967),
.B(n_709),
.Y(n_12883)
);

NOR2xp33_ASAP7_75t_L g12884 ( 
.A(n_12622),
.B(n_12337),
.Y(n_12884)
);

NAND2xp5_ASAP7_75t_L g12885 ( 
.A(n_12412),
.B(n_710),
.Y(n_12885)
);

AOI21xp5_ASAP7_75t_L g12886 ( 
.A1(n_12506),
.A2(n_5257),
.B(n_5255),
.Y(n_12886)
);

AOI21xp5_ASAP7_75t_L g12887 ( 
.A1(n_12517),
.A2(n_5260),
.B(n_5258),
.Y(n_12887)
);

NOR2xp33_ASAP7_75t_L g12888 ( 
.A(n_12353),
.B(n_712),
.Y(n_12888)
);

BUFx6f_ASAP7_75t_L g12889 ( 
.A(n_11968),
.Y(n_12889)
);

NOR3xp33_ASAP7_75t_L g12890 ( 
.A(n_12581),
.B(n_712),
.C(n_713),
.Y(n_12890)
);

AOI22xp5_ASAP7_75t_L g12891 ( 
.A1(n_12582),
.A2(n_715),
.B1(n_713),
.B2(n_714),
.Y(n_12891)
);

INVx2_ASAP7_75t_L g12892 ( 
.A(n_11991),
.Y(n_12892)
);

INVx2_ASAP7_75t_L g12893 ( 
.A(n_12015),
.Y(n_12893)
);

AND2x2_ASAP7_75t_L g12894 ( 
.A(n_12472),
.B(n_714),
.Y(n_12894)
);

BUFx2_ASAP7_75t_L g12895 ( 
.A(n_12068),
.Y(n_12895)
);

AOI21x1_ASAP7_75t_L g12896 ( 
.A1(n_12688),
.A2(n_715),
.B(n_716),
.Y(n_12896)
);

OAI22xp5_ASAP7_75t_L g12897 ( 
.A1(n_12611),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_12897)
);

INVx1_ASAP7_75t_L g12898 ( 
.A(n_12032),
.Y(n_12898)
);

AOI22xp5_ASAP7_75t_L g12899 ( 
.A1(n_12610),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_12899)
);

NAND2xp5_ASAP7_75t_L g12900 ( 
.A(n_12445),
.B(n_719),
.Y(n_12900)
);

OR2x6_ASAP7_75t_SL g12901 ( 
.A(n_12471),
.B(n_720),
.Y(n_12901)
);

AOI21x1_ASAP7_75t_L g12902 ( 
.A1(n_12693),
.A2(n_720),
.B(n_721),
.Y(n_12902)
);

NAND2xp5_ASAP7_75t_SL g12903 ( 
.A(n_12601),
.B(n_5262),
.Y(n_12903)
);

AOI21xp5_ASAP7_75t_L g12904 ( 
.A1(n_12530),
.A2(n_12553),
.B(n_12549),
.Y(n_12904)
);

O2A1O1Ixp33_ASAP7_75t_L g12905 ( 
.A1(n_12523),
.A2(n_723),
.B(n_721),
.C(n_722),
.Y(n_12905)
);

AOI21xp5_ASAP7_75t_L g12906 ( 
.A1(n_12556),
.A2(n_5264),
.B(n_5263),
.Y(n_12906)
);

AOI21xp5_ASAP7_75t_L g12907 ( 
.A1(n_12576),
.A2(n_12645),
.B(n_12612),
.Y(n_12907)
);

O2A1O1Ixp5_ASAP7_75t_L g12908 ( 
.A1(n_12544),
.A2(n_724),
.B(n_722),
.C(n_723),
.Y(n_12908)
);

INVx1_ASAP7_75t_L g12909 ( 
.A(n_12080),
.Y(n_12909)
);

INVx1_ASAP7_75t_L g12910 ( 
.A(n_12118),
.Y(n_12910)
);

AND2x4_ASAP7_75t_L g12911 ( 
.A(n_11986),
.B(n_5265),
.Y(n_12911)
);

NAND2xp5_ASAP7_75t_L g12912 ( 
.A(n_12424),
.B(n_724),
.Y(n_12912)
);

INVx3_ASAP7_75t_L g12913 ( 
.A(n_12097),
.Y(n_12913)
);

INVx1_ASAP7_75t_L g12914 ( 
.A(n_12126),
.Y(n_12914)
);

NAND3xp33_ASAP7_75t_SL g12915 ( 
.A(n_12630),
.B(n_725),
.C(n_726),
.Y(n_12915)
);

CKINVDCx20_ASAP7_75t_R g12916 ( 
.A(n_12079),
.Y(n_12916)
);

AND2x4_ASAP7_75t_L g12917 ( 
.A(n_12198),
.B(n_5267),
.Y(n_12917)
);

NOR2xp67_ASAP7_75t_SL g12918 ( 
.A(n_12122),
.B(n_5268),
.Y(n_12918)
);

AOI22xp5_ASAP7_75t_L g12919 ( 
.A1(n_12692),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.Y(n_12919)
);

INVx2_ASAP7_75t_L g12920 ( 
.A(n_12197),
.Y(n_12920)
);

AO22x1_ASAP7_75t_L g12921 ( 
.A1(n_12265),
.A2(n_731),
.B1(n_728),
.B2(n_730),
.Y(n_12921)
);

NAND2xp5_ASAP7_75t_SL g12922 ( 
.A(n_12710),
.B(n_5269),
.Y(n_12922)
);

NAND2xp5_ASAP7_75t_SL g12923 ( 
.A(n_12738),
.B(n_5270),
.Y(n_12923)
);

AND2x2_ASAP7_75t_L g12924 ( 
.A(n_12431),
.B(n_12255),
.Y(n_12924)
);

AOI22xp33_ASAP7_75t_L g12925 ( 
.A1(n_12040),
.A2(n_732),
.B1(n_728),
.B2(n_731),
.Y(n_12925)
);

BUFx6f_ASAP7_75t_L g12926 ( 
.A(n_11968),
.Y(n_12926)
);

OAI22xp5_ASAP7_75t_L g12927 ( 
.A1(n_12641),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_12285),
.Y(n_12928)
);

AOI21x1_ASAP7_75t_L g12929 ( 
.A1(n_12721),
.A2(n_733),
.B(n_735),
.Y(n_12929)
);

NAND2xp5_ASAP7_75t_L g12930 ( 
.A(n_12340),
.B(n_735),
.Y(n_12930)
);

AO22x1_ASAP7_75t_L g12931 ( 
.A1(n_12777),
.A2(n_738),
.B1(n_736),
.B2(n_737),
.Y(n_12931)
);

OA22x2_ASAP7_75t_L g12932 ( 
.A1(n_12454),
.A2(n_738),
.B1(n_736),
.B2(n_737),
.Y(n_12932)
);

NAND2xp5_ASAP7_75t_L g12933 ( 
.A(n_12323),
.B(n_739),
.Y(n_12933)
);

INVx1_ASAP7_75t_L g12934 ( 
.A(n_12288),
.Y(n_12934)
);

INVx2_ASAP7_75t_L g12935 ( 
.A(n_12325),
.Y(n_12935)
);

INVx3_ASAP7_75t_L g12936 ( 
.A(n_12101),
.Y(n_12936)
);

AOI21xp5_ASAP7_75t_L g12937 ( 
.A1(n_12646),
.A2(n_12704),
.B(n_12654),
.Y(n_12937)
);

AOI21xp5_ASAP7_75t_L g12938 ( 
.A1(n_12744),
.A2(n_5273),
.B(n_5271),
.Y(n_12938)
);

OAI21x1_ASAP7_75t_L g12939 ( 
.A1(n_12213),
.A2(n_5275),
.B(n_5274),
.Y(n_12939)
);

NAND2xp5_ASAP7_75t_L g12940 ( 
.A(n_12377),
.B(n_740),
.Y(n_12940)
);

AOI21x1_ASAP7_75t_L g12941 ( 
.A1(n_12435),
.A2(n_740),
.B(n_741),
.Y(n_12941)
);

NOR2xp33_ASAP7_75t_L g12942 ( 
.A(n_12368),
.B(n_741),
.Y(n_12942)
);

NAND2xp5_ASAP7_75t_SL g12943 ( 
.A(n_12781),
.B(n_5276),
.Y(n_12943)
);

AOI21xp5_ASAP7_75t_L g12944 ( 
.A1(n_12189),
.A2(n_11944),
.B(n_12500),
.Y(n_12944)
);

AOI21xp5_ASAP7_75t_L g12945 ( 
.A1(n_12504),
.A2(n_5282),
.B(n_5279),
.Y(n_12945)
);

AOI21xp5_ASAP7_75t_L g12946 ( 
.A1(n_12510),
.A2(n_5284),
.B(n_5283),
.Y(n_12946)
);

NAND2xp5_ASAP7_75t_SL g12947 ( 
.A(n_12679),
.B(n_5285),
.Y(n_12947)
);

AOI21xp5_ASAP7_75t_L g12948 ( 
.A1(n_12514),
.A2(n_5287),
.B(n_5286),
.Y(n_12948)
);

AOI21xp5_ASAP7_75t_L g12949 ( 
.A1(n_12518),
.A2(n_5290),
.B(n_5288),
.Y(n_12949)
);

NAND2xp5_ASAP7_75t_L g12950 ( 
.A(n_11964),
.B(n_742),
.Y(n_12950)
);

NAND2xp5_ASAP7_75t_SL g12951 ( 
.A(n_11975),
.B(n_5291),
.Y(n_12951)
);

AND2x2_ASAP7_75t_L g12952 ( 
.A(n_12369),
.B(n_742),
.Y(n_12952)
);

AOI21x1_ASAP7_75t_L g12953 ( 
.A1(n_12493),
.A2(n_743),
.B(n_744),
.Y(n_12953)
);

AND2x2_ASAP7_75t_L g12954 ( 
.A(n_12374),
.B(n_743),
.Y(n_12954)
);

INVx1_ASAP7_75t_SL g12955 ( 
.A(n_12050),
.Y(n_12955)
);

AOI21xp5_ASAP7_75t_L g12956 ( 
.A1(n_12522),
.A2(n_5294),
.B(n_5292),
.Y(n_12956)
);

O2A1O1Ixp5_ASAP7_75t_L g12957 ( 
.A1(n_12244),
.A2(n_746),
.B(n_744),
.C(n_745),
.Y(n_12957)
);

OR2x2_ASAP7_75t_L g12958 ( 
.A(n_12301),
.B(n_745),
.Y(n_12958)
);

NAND2xp5_ASAP7_75t_SL g12959 ( 
.A(n_12626),
.B(n_5295),
.Y(n_12959)
);

NOR2xp33_ASAP7_75t_L g12960 ( 
.A(n_12383),
.B(n_746),
.Y(n_12960)
);

NOR2xp33_ASAP7_75t_L g12961 ( 
.A(n_12045),
.B(n_747),
.Y(n_12961)
);

AND2x2_ASAP7_75t_L g12962 ( 
.A(n_12508),
.B(n_747),
.Y(n_12962)
);

NAND2xp5_ASAP7_75t_SL g12963 ( 
.A(n_12715),
.B(n_5296),
.Y(n_12963)
);

AND2x2_ASAP7_75t_L g12964 ( 
.A(n_12512),
.B(n_748),
.Y(n_12964)
);

NAND2xp5_ASAP7_75t_SL g12965 ( 
.A(n_12786),
.B(n_5297),
.Y(n_12965)
);

A2O1A1Ixp33_ASAP7_75t_L g12966 ( 
.A1(n_12144),
.A2(n_12211),
.B(n_12624),
.C(n_12528),
.Y(n_12966)
);

NAND2xp5_ASAP7_75t_L g12967 ( 
.A(n_11969),
.B(n_748),
.Y(n_12967)
);

AND2x4_ASAP7_75t_L g12968 ( 
.A(n_12226),
.B(n_5298),
.Y(n_12968)
);

BUFx6f_ASAP7_75t_L g12969 ( 
.A(n_11968),
.Y(n_12969)
);

AOI21xp5_ASAP7_75t_L g12970 ( 
.A1(n_12538),
.A2(n_12559),
.B(n_12540),
.Y(n_12970)
);

NAND2xp5_ASAP7_75t_L g12971 ( 
.A(n_12003),
.B(n_12037),
.Y(n_12971)
);

O2A1O1Ixp5_ASAP7_75t_L g12972 ( 
.A1(n_12257),
.A2(n_752),
.B(n_750),
.C(n_751),
.Y(n_12972)
);

INVx1_ASAP7_75t_L g12973 ( 
.A(n_12529),
.Y(n_12973)
);

AOI21xp5_ASAP7_75t_L g12974 ( 
.A1(n_12565),
.A2(n_5300),
.B(n_5299),
.Y(n_12974)
);

NOR2xp67_ASAP7_75t_SL g12975 ( 
.A(n_12156),
.B(n_5301),
.Y(n_12975)
);

NAND2xp5_ASAP7_75t_L g12976 ( 
.A(n_12063),
.B(n_750),
.Y(n_12976)
);

AND2x2_ASAP7_75t_L g12977 ( 
.A(n_12578),
.B(n_751),
.Y(n_12977)
);

AOI21xp5_ASAP7_75t_L g12978 ( 
.A1(n_12571),
.A2(n_5303),
.B(n_5302),
.Y(n_12978)
);

AOI21xp5_ASAP7_75t_L g12979 ( 
.A1(n_12580),
.A2(n_5306),
.B(n_5304),
.Y(n_12979)
);

O2A1O1Ixp33_ASAP7_75t_L g12980 ( 
.A1(n_12532),
.A2(n_12547),
.B(n_12594),
.C(n_12555),
.Y(n_12980)
);

BUFx4f_ASAP7_75t_SL g12981 ( 
.A(n_12558),
.Y(n_12981)
);

INVx2_ASAP7_75t_L g12982 ( 
.A(n_12620),
.Y(n_12982)
);

INVx1_ASAP7_75t_L g12983 ( 
.A(n_12655),
.Y(n_12983)
);

AOI21xp5_ASAP7_75t_L g12984 ( 
.A1(n_12583),
.A2(n_5309),
.B(n_5308),
.Y(n_12984)
);

AND2x2_ASAP7_75t_L g12985 ( 
.A(n_12667),
.B(n_12687),
.Y(n_12985)
);

NAND2xp5_ASAP7_75t_L g12986 ( 
.A(n_12066),
.B(n_752),
.Y(n_12986)
);

INVx1_ASAP7_75t_L g12987 ( 
.A(n_12734),
.Y(n_12987)
);

AOI21xp5_ASAP7_75t_L g12988 ( 
.A1(n_12585),
.A2(n_5313),
.B(n_5312),
.Y(n_12988)
);

INVx1_ASAP7_75t_L g12989 ( 
.A(n_12736),
.Y(n_12989)
);

NAND2xp5_ASAP7_75t_L g12990 ( 
.A(n_12073),
.B(n_753),
.Y(n_12990)
);

INVx3_ASAP7_75t_L g12991 ( 
.A(n_12101),
.Y(n_12991)
);

OAI21x1_ASAP7_75t_L g12992 ( 
.A1(n_12363),
.A2(n_5315),
.B(n_5314),
.Y(n_12992)
);

INVx8_ASAP7_75t_L g12993 ( 
.A(n_12380),
.Y(n_12993)
);

NOR2xp67_ASAP7_75t_L g12994 ( 
.A(n_12191),
.B(n_753),
.Y(n_12994)
);

BUFx4f_ASAP7_75t_L g12995 ( 
.A(n_12142),
.Y(n_12995)
);

OAI21xp33_ASAP7_75t_L g12996 ( 
.A1(n_11956),
.A2(n_12754),
.B(n_12224),
.Y(n_12996)
);

NOR2xp33_ASAP7_75t_L g12997 ( 
.A(n_12733),
.B(n_754),
.Y(n_12997)
);

OAI22xp5_ASAP7_75t_L g12998 ( 
.A1(n_12410),
.A2(n_756),
.B1(n_754),
.B2(n_755),
.Y(n_12998)
);

NAND2xp5_ASAP7_75t_L g12999 ( 
.A(n_12082),
.B(n_755),
.Y(n_12999)
);

OR2x2_ASAP7_75t_L g13000 ( 
.A(n_12745),
.B(n_756),
.Y(n_13000)
);

NAND3xp33_ASAP7_75t_L g13001 ( 
.A(n_12235),
.B(n_757),
.C(n_758),
.Y(n_13001)
);

AOI21xp5_ASAP7_75t_L g13002 ( 
.A1(n_12586),
.A2(n_5317),
.B(n_5316),
.Y(n_13002)
);

OAI22xp5_ASAP7_75t_L g13003 ( 
.A1(n_11942),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_13003)
);

AOI21xp5_ASAP7_75t_L g13004 ( 
.A1(n_12591),
.A2(n_5319),
.B(n_5318),
.Y(n_13004)
);

AND2x2_ASAP7_75t_L g13005 ( 
.A(n_12023),
.B(n_12389),
.Y(n_13005)
);

OAI21xp5_ASAP7_75t_L g13006 ( 
.A1(n_12695),
.A2(n_5321),
.B(n_5320),
.Y(n_13006)
);

NAND2xp5_ASAP7_75t_L g13007 ( 
.A(n_12139),
.B(n_759),
.Y(n_13007)
);

INVx1_ASAP7_75t_L g13008 ( 
.A(n_12398),
.Y(n_13008)
);

AOI21x1_ASAP7_75t_L g13009 ( 
.A1(n_11983),
.A2(n_12166),
.B(n_12498),
.Y(n_13009)
);

BUFx8_ASAP7_75t_L g13010 ( 
.A(n_12199),
.Y(n_13010)
);

AOI21xp5_ASAP7_75t_L g13011 ( 
.A1(n_12602),
.A2(n_5323),
.B(n_5322),
.Y(n_13011)
);

BUFx6f_ASAP7_75t_L g13012 ( 
.A(n_11943),
.Y(n_13012)
);

INVx1_ASAP7_75t_L g13013 ( 
.A(n_12373),
.Y(n_13013)
);

NOR2xp33_ASAP7_75t_L g13014 ( 
.A(n_12616),
.B(n_760),
.Y(n_13014)
);

OAI21xp5_ASAP7_75t_L g13015 ( 
.A1(n_12699),
.A2(n_5326),
.B(n_5325),
.Y(n_13015)
);

NAND2xp5_ASAP7_75t_L g13016 ( 
.A(n_12152),
.B(n_760),
.Y(n_13016)
);

NAND2xp5_ASAP7_75t_L g13017 ( 
.A(n_12168),
.B(n_761),
.Y(n_13017)
);

INVx1_ASAP7_75t_L g13018 ( 
.A(n_12385),
.Y(n_13018)
);

INVx3_ASAP7_75t_L g13019 ( 
.A(n_12101),
.Y(n_13019)
);

AOI21xp5_ASAP7_75t_L g13020 ( 
.A1(n_12615),
.A2(n_5329),
.B(n_5328),
.Y(n_13020)
);

NAND2xp5_ASAP7_75t_SL g13021 ( 
.A(n_12173),
.B(n_5330),
.Y(n_13021)
);

NAND2xp5_ASAP7_75t_SL g13022 ( 
.A(n_12730),
.B(n_5331),
.Y(n_13022)
);

NOR2xp67_ASAP7_75t_L g13023 ( 
.A(n_12089),
.B(n_761),
.Y(n_13023)
);

NAND2xp5_ASAP7_75t_L g13024 ( 
.A(n_12188),
.B(n_762),
.Y(n_13024)
);

NAND2xp5_ASAP7_75t_SL g13025 ( 
.A(n_12780),
.B(n_5332),
.Y(n_13025)
);

NAND2xp5_ASAP7_75t_L g13026 ( 
.A(n_12502),
.B(n_762),
.Y(n_13026)
);

AOI21xp5_ASAP7_75t_L g13027 ( 
.A1(n_12628),
.A2(n_5334),
.B(n_5333),
.Y(n_13027)
);

AOI21xp5_ASAP7_75t_L g13028 ( 
.A1(n_12639),
.A2(n_5337),
.B(n_5336),
.Y(n_13028)
);

AOI22xp5_ASAP7_75t_L g13029 ( 
.A1(n_12782),
.A2(n_765),
.B1(n_763),
.B2(n_764),
.Y(n_13029)
);

NAND2xp5_ASAP7_75t_L g13030 ( 
.A(n_12503),
.B(n_763),
.Y(n_13030)
);

AOI221xp5_ASAP7_75t_L g13031 ( 
.A1(n_12411),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.C(n_767),
.Y(n_13031)
);

NAND2xp5_ASAP7_75t_L g13032 ( 
.A(n_12516),
.B(n_766),
.Y(n_13032)
);

OAI21xp33_ASAP7_75t_L g13033 ( 
.A1(n_11990),
.A2(n_767),
.B(n_768),
.Y(n_13033)
);

OR2x6_ASAP7_75t_L g13034 ( 
.A(n_12305),
.B(n_5338),
.Y(n_13034)
);

AOI21xp5_ASAP7_75t_L g13035 ( 
.A1(n_12653),
.A2(n_12659),
.B(n_12658),
.Y(n_13035)
);

NAND2xp5_ASAP7_75t_SL g13036 ( 
.A(n_12309),
.B(n_5339),
.Y(n_13036)
);

NAND2xp5_ASAP7_75t_SL g13037 ( 
.A(n_12252),
.B(n_5340),
.Y(n_13037)
);

NOR2x1_ASAP7_75t_L g13038 ( 
.A(n_12494),
.B(n_768),
.Y(n_13038)
);

AOI21xp5_ASAP7_75t_L g13039 ( 
.A1(n_12662),
.A2(n_5342),
.B(n_5341),
.Y(n_13039)
);

BUFx3_ASAP7_75t_L g13040 ( 
.A(n_12178),
.Y(n_13040)
);

BUFx2_ASAP7_75t_L g13041 ( 
.A(n_12481),
.Y(n_13041)
);

NAND2xp5_ASAP7_75t_L g13042 ( 
.A(n_12520),
.B(n_12526),
.Y(n_13042)
);

AOI21xp5_ASAP7_75t_L g13043 ( 
.A1(n_12668),
.A2(n_5344),
.B(n_5343),
.Y(n_13043)
);

NAND2xp5_ASAP7_75t_L g13044 ( 
.A(n_12531),
.B(n_770),
.Y(n_13044)
);

BUFx2_ASAP7_75t_L g13045 ( 
.A(n_12438),
.Y(n_13045)
);

INVx4_ASAP7_75t_L g13046 ( 
.A(n_12507),
.Y(n_13046)
);

AOI21xp5_ASAP7_75t_L g13047 ( 
.A1(n_12669),
.A2(n_5346),
.B(n_5345),
.Y(n_13047)
);

INVx2_ASAP7_75t_L g13048 ( 
.A(n_12536),
.Y(n_13048)
);

NOR2xp33_ASAP7_75t_L g13049 ( 
.A(n_12187),
.B(n_770),
.Y(n_13049)
);

NAND2xp5_ASAP7_75t_L g13050 ( 
.A(n_12543),
.B(n_771),
.Y(n_13050)
);

O2A1O1Ixp33_ASAP7_75t_L g13051 ( 
.A1(n_12605),
.A2(n_774),
.B(n_772),
.C(n_773),
.Y(n_13051)
);

INVx1_ASAP7_75t_L g13052 ( 
.A(n_12261),
.Y(n_13052)
);

AO21x1_ASAP7_75t_L g13053 ( 
.A1(n_12345),
.A2(n_772),
.B(n_773),
.Y(n_13053)
);

INVx11_ASAP7_75t_L g13054 ( 
.A(n_12014),
.Y(n_13054)
);

AND2x4_ASAP7_75t_L g13055 ( 
.A(n_12451),
.B(n_5347),
.Y(n_13055)
);

OAI22xp5_ASAP7_75t_L g13056 ( 
.A1(n_12312),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_13056)
);

NAND2xp5_ASAP7_75t_SL g13057 ( 
.A(n_12505),
.B(n_5348),
.Y(n_13057)
);

NAND2xp5_ASAP7_75t_L g13058 ( 
.A(n_12550),
.B(n_775),
.Y(n_13058)
);

OAI21x1_ASAP7_75t_L g13059 ( 
.A1(n_12348),
.A2(n_5350),
.B(n_5349),
.Y(n_13059)
);

OAI21xp33_ASAP7_75t_L g13060 ( 
.A1(n_12194),
.A2(n_776),
.B(n_777),
.Y(n_13060)
);

NOR2xp33_ASAP7_75t_L g13061 ( 
.A(n_12026),
.B(n_778),
.Y(n_13061)
);

INVx2_ASAP7_75t_L g13062 ( 
.A(n_12569),
.Y(n_13062)
);

NAND2xp5_ASAP7_75t_L g13063 ( 
.A(n_12574),
.B(n_778),
.Y(n_13063)
);

OAI22xp5_ASAP7_75t_L g13064 ( 
.A1(n_12074),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_13064)
);

AOI21xp5_ASAP7_75t_L g13065 ( 
.A1(n_12670),
.A2(n_12683),
.B(n_12677),
.Y(n_13065)
);

INVx1_ASAP7_75t_L g13066 ( 
.A(n_12277),
.Y(n_13066)
);

NAND2xp5_ASAP7_75t_L g13067 ( 
.A(n_12577),
.B(n_781),
.Y(n_13067)
);

INVx2_ASAP7_75t_L g13068 ( 
.A(n_12771),
.Y(n_13068)
);

AOI21x1_ASAP7_75t_L g13069 ( 
.A1(n_12034),
.A2(n_782),
.B(n_783),
.Y(n_13069)
);

NOR2xp33_ASAP7_75t_L g13070 ( 
.A(n_12482),
.B(n_782),
.Y(n_13070)
);

NAND2xp5_ASAP7_75t_L g13071 ( 
.A(n_12614),
.B(n_783),
.Y(n_13071)
);

OAI22xp5_ASAP7_75t_L g13072 ( 
.A1(n_12231),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.Y(n_13072)
);

NOR2xp33_ASAP7_75t_L g13073 ( 
.A(n_11939),
.B(n_12521),
.Y(n_13073)
);

OAI21xp33_ASAP7_75t_L g13074 ( 
.A1(n_12210),
.A2(n_784),
.B(n_785),
.Y(n_13074)
);

AOI21xp5_ASAP7_75t_L g13075 ( 
.A1(n_12685),
.A2(n_5353),
.B(n_5352),
.Y(n_13075)
);

AOI21xp5_ASAP7_75t_L g13076 ( 
.A1(n_12702),
.A2(n_5355),
.B(n_5354),
.Y(n_13076)
);

CKINVDCx5p33_ASAP7_75t_R g13077 ( 
.A(n_12072),
.Y(n_13077)
);

INVx1_ASAP7_75t_L g13078 ( 
.A(n_12316),
.Y(n_13078)
);

AOI21xp5_ASAP7_75t_L g13079 ( 
.A1(n_12706),
.A2(n_5358),
.B(n_5356),
.Y(n_13079)
);

NOR2xp33_ASAP7_75t_R g13080 ( 
.A(n_12250),
.B(n_5359),
.Y(n_13080)
);

AND2x2_ASAP7_75t_L g13081 ( 
.A(n_12475),
.B(n_786),
.Y(n_13081)
);

A2O1A1Ixp33_ASAP7_75t_L g13082 ( 
.A1(n_12234),
.A2(n_789),
.B(n_787),
.C(n_788),
.Y(n_13082)
);

INVx3_ASAP7_75t_L g13083 ( 
.A(n_11943),
.Y(n_13083)
);

INVx2_ASAP7_75t_L g13084 ( 
.A(n_12627),
.Y(n_13084)
);

AOI21xp5_ASAP7_75t_L g13085 ( 
.A1(n_12707),
.A2(n_5362),
.B(n_5360),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12397),
.Y(n_13086)
);

CKINVDCx5p33_ASAP7_75t_R g13087 ( 
.A(n_12449),
.Y(n_13087)
);

AOI22xp5_ASAP7_75t_L g13088 ( 
.A1(n_12392),
.A2(n_790),
.B1(n_788),
.B2(n_789),
.Y(n_13088)
);

INVx1_ASAP7_75t_L g13089 ( 
.A(n_12225),
.Y(n_13089)
);

AND2x2_ASAP7_75t_SL g13090 ( 
.A(n_12495),
.B(n_790),
.Y(n_13090)
);

INVxp67_ASAP7_75t_SL g13091 ( 
.A(n_12242),
.Y(n_13091)
);

INVx2_ASAP7_75t_L g13092 ( 
.A(n_12647),
.Y(n_13092)
);

NAND2xp5_ASAP7_75t_SL g13093 ( 
.A(n_12775),
.B(n_5366),
.Y(n_13093)
);

AOI21xp5_ASAP7_75t_L g13094 ( 
.A1(n_12711),
.A2(n_5368),
.B(n_5367),
.Y(n_13094)
);

O2A1O1Ixp33_ASAP7_75t_L g13095 ( 
.A1(n_12650),
.A2(n_793),
.B(n_791),
.C(n_792),
.Y(n_13095)
);

AOI21xp5_ASAP7_75t_L g13096 ( 
.A1(n_12714),
.A2(n_5370),
.B(n_5369),
.Y(n_13096)
);

NAND2xp5_ASAP7_75t_L g13097 ( 
.A(n_12657),
.B(n_791),
.Y(n_13097)
);

A2O1A1Ixp33_ASAP7_75t_L g13098 ( 
.A1(n_12179),
.A2(n_795),
.B(n_792),
.C(n_794),
.Y(n_13098)
);

NAND2xp5_ASAP7_75t_L g13099 ( 
.A(n_12686),
.B(n_794),
.Y(n_13099)
);

AOI22xp5_ASAP7_75t_L g13100 ( 
.A1(n_12696),
.A2(n_797),
.B1(n_795),
.B2(n_796),
.Y(n_13100)
);

NOR2xp33_ASAP7_75t_L g13101 ( 
.A(n_12572),
.B(n_796),
.Y(n_13101)
);

AOI22xp5_ASAP7_75t_L g13102 ( 
.A1(n_12275),
.A2(n_799),
.B1(n_797),
.B2(n_798),
.Y(n_13102)
);

AO32x2_ASAP7_75t_L g13103 ( 
.A1(n_12491),
.A2(n_800),
.A3(n_798),
.B1(n_799),
.B2(n_801),
.Y(n_13103)
);

AND2x2_ASAP7_75t_SL g13104 ( 
.A(n_12467),
.B(n_800),
.Y(n_13104)
);

AOI22xp5_ASAP7_75t_L g13105 ( 
.A1(n_12005),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_13105)
);

AOI21xp5_ASAP7_75t_L g13106 ( 
.A1(n_12716),
.A2(n_5372),
.B(n_5371),
.Y(n_13106)
);

NAND2xp5_ASAP7_75t_SL g13107 ( 
.A(n_12237),
.B(n_5373),
.Y(n_13107)
);

NAND2xp5_ASAP7_75t_L g13108 ( 
.A(n_12713),
.B(n_802),
.Y(n_13108)
);

AOI21xp5_ASAP7_75t_L g13109 ( 
.A1(n_12719),
.A2(n_5376),
.B(n_5375),
.Y(n_13109)
);

INVxp67_ASAP7_75t_L g13110 ( 
.A(n_12631),
.Y(n_13110)
);

INVx1_ASAP7_75t_L g13111 ( 
.A(n_12748),
.Y(n_13111)
);

AOI21xp5_ASAP7_75t_L g13112 ( 
.A1(n_12724),
.A2(n_5378),
.B(n_5377),
.Y(n_13112)
);

NAND2xp5_ASAP7_75t_SL g13113 ( 
.A(n_12426),
.B(n_5380),
.Y(n_13113)
);

BUFx2_ASAP7_75t_L g13114 ( 
.A(n_11943),
.Y(n_13114)
);

NOR3xp33_ASAP7_75t_L g13115 ( 
.A(n_12355),
.B(n_803),
.C(n_805),
.Y(n_13115)
);

NOR2xp33_ASAP7_75t_L g13116 ( 
.A(n_12644),
.B(n_805),
.Y(n_13116)
);

NAND2xp5_ASAP7_75t_SL g13117 ( 
.A(n_12429),
.B(n_5381),
.Y(n_13117)
);

OR2x2_ASAP7_75t_L g13118 ( 
.A(n_12170),
.B(n_806),
.Y(n_13118)
);

OR2x6_ASAP7_75t_SL g13119 ( 
.A(n_12407),
.B(n_806),
.Y(n_13119)
);

NAND2xp5_ASAP7_75t_SL g13120 ( 
.A(n_12104),
.B(n_5384),
.Y(n_13120)
);

NOR2x1_ASAP7_75t_L g13121 ( 
.A(n_12043),
.B(n_807),
.Y(n_13121)
);

INVx2_ASAP7_75t_L g13122 ( 
.A(n_12760),
.Y(n_13122)
);

AND2x2_ASAP7_75t_L g13123 ( 
.A(n_11988),
.B(n_807),
.Y(n_13123)
);

AOI21xp5_ASAP7_75t_L g13124 ( 
.A1(n_12725),
.A2(n_5386),
.B(n_5385),
.Y(n_13124)
);

INVx2_ASAP7_75t_L g13125 ( 
.A(n_12209),
.Y(n_13125)
);

INVx4_ASAP7_75t_L g13126 ( 
.A(n_12600),
.Y(n_13126)
);

OAI21xp5_ASAP7_75t_L g13127 ( 
.A1(n_12741),
.A2(n_12750),
.B(n_12747),
.Y(n_13127)
);

AOI21xp5_ASAP7_75t_L g13128 ( 
.A1(n_12768),
.A2(n_5389),
.B(n_5387),
.Y(n_13128)
);

NAND2xp5_ASAP7_75t_L g13129 ( 
.A(n_12221),
.B(n_808),
.Y(n_13129)
);

AND2x2_ASAP7_75t_SL g13130 ( 
.A(n_12047),
.B(n_808),
.Y(n_13130)
);

NAND2xp5_ASAP7_75t_L g13131 ( 
.A(n_12232),
.B(n_809),
.Y(n_13131)
);

INVx1_ASAP7_75t_L g13132 ( 
.A(n_12281),
.Y(n_13132)
);

AND2x2_ASAP7_75t_L g13133 ( 
.A(n_12525),
.B(n_809),
.Y(n_13133)
);

AOI22xp5_ASAP7_75t_L g13134 ( 
.A1(n_12008),
.A2(n_812),
.B1(n_810),
.B2(n_811),
.Y(n_13134)
);

NAND2xp5_ASAP7_75t_L g13135 ( 
.A(n_12331),
.B(n_810),
.Y(n_13135)
);

INVx3_ASAP7_75t_L g13136 ( 
.A(n_11966),
.Y(n_13136)
);

INVx2_ASAP7_75t_SL g13137 ( 
.A(n_11966),
.Y(n_13137)
);

OAI22xp5_ASAP7_75t_L g13138 ( 
.A1(n_12249),
.A2(n_813),
.B1(n_811),
.B2(n_812),
.Y(n_13138)
);

AOI21xp5_ASAP7_75t_L g13139 ( 
.A1(n_12770),
.A2(n_5391),
.B(n_5390),
.Y(n_13139)
);

BUFx3_ASAP7_75t_L g13140 ( 
.A(n_12142),
.Y(n_13140)
);

OAI22xp5_ASAP7_75t_L g13141 ( 
.A1(n_12263),
.A2(n_12095),
.B1(n_12164),
.B2(n_12162),
.Y(n_13141)
);

NAND2xp5_ASAP7_75t_L g13142 ( 
.A(n_12356),
.B(n_813),
.Y(n_13142)
);

NAND2xp5_ASAP7_75t_L g13143 ( 
.A(n_12404),
.B(n_814),
.Y(n_13143)
);

INVx3_ASAP7_75t_SL g13144 ( 
.A(n_12142),
.Y(n_13144)
);

INVx1_ASAP7_75t_L g13145 ( 
.A(n_12358),
.Y(n_13145)
);

AND2x6_ASAP7_75t_SL g13146 ( 
.A(n_12480),
.B(n_814),
.Y(n_13146)
);

AOI21xp5_ASAP7_75t_L g13147 ( 
.A1(n_12776),
.A2(n_12783),
.B(n_12779),
.Y(n_13147)
);

AND2x2_ASAP7_75t_SL g13148 ( 
.A(n_12273),
.B(n_815),
.Y(n_13148)
);

NAND2xp5_ASAP7_75t_SL g13149 ( 
.A(n_12200),
.B(n_12282),
.Y(n_13149)
);

AND2x2_ASAP7_75t_SL g13150 ( 
.A(n_12479),
.B(n_816),
.Y(n_13150)
);

AOI221xp5_ASAP7_75t_L g13151 ( 
.A1(n_12293),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.C(n_819),
.Y(n_13151)
);

HB1xp67_ASAP7_75t_L g13152 ( 
.A(n_12497),
.Y(n_13152)
);

NAND2xp5_ASAP7_75t_SL g13153 ( 
.A(n_12350),
.B(n_12013),
.Y(n_13153)
);

AOI21xp5_ASAP7_75t_L g13154 ( 
.A1(n_12788),
.A2(n_5393),
.B(n_5392),
.Y(n_13154)
);

INVx1_ASAP7_75t_SL g13155 ( 
.A(n_12289),
.Y(n_13155)
);

OAI22xp5_ASAP7_75t_L g13156 ( 
.A1(n_12317),
.A2(n_820),
.B1(n_817),
.B2(n_819),
.Y(n_13156)
);

INVx3_ASAP7_75t_L g13157 ( 
.A(n_11966),
.Y(n_13157)
);

INVx2_ASAP7_75t_L g13158 ( 
.A(n_12341),
.Y(n_13158)
);

AO32x1_ASAP7_75t_L g13159 ( 
.A1(n_12485),
.A2(n_822),
.A3(n_820),
.B1(n_821),
.B2(n_823),
.Y(n_13159)
);

INVx2_ASAP7_75t_L g13160 ( 
.A(n_12357),
.Y(n_13160)
);

OAI22xp5_ASAP7_75t_L g13161 ( 
.A1(n_12584),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.Y(n_13161)
);

AND2x2_ASAP7_75t_SL g13162 ( 
.A(n_12455),
.B(n_824),
.Y(n_13162)
);

A2O1A1Ixp33_ASAP7_75t_SL g13163 ( 
.A1(n_12048),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_13163)
);

OA22x2_ASAP7_75t_L g13164 ( 
.A1(n_12413),
.A2(n_827),
.B1(n_825),
.B2(n_826),
.Y(n_13164)
);

NAND2xp5_ASAP7_75t_L g13165 ( 
.A(n_12390),
.B(n_827),
.Y(n_13165)
);

NOR2xp33_ASAP7_75t_SL g13166 ( 
.A(n_12128),
.B(n_5394),
.Y(n_13166)
);

AND2x2_ASAP7_75t_L g13167 ( 
.A(n_12608),
.B(n_828),
.Y(n_13167)
);

AO22x1_ASAP7_75t_L g13168 ( 
.A1(n_12394),
.A2(n_830),
.B1(n_828),
.B2(n_829),
.Y(n_13168)
);

A2O1A1Ixp33_ASAP7_75t_L g13169 ( 
.A1(n_12105),
.A2(n_832),
.B(n_829),
.C(n_831),
.Y(n_13169)
);

NAND2xp5_ASAP7_75t_L g13170 ( 
.A(n_12298),
.B(n_831),
.Y(n_13170)
);

INVx4_ASAP7_75t_L g13171 ( 
.A(n_12380),
.Y(n_13171)
);

AOI21xp5_ASAP7_75t_L g13172 ( 
.A1(n_11948),
.A2(n_5396),
.B(n_5395),
.Y(n_13172)
);

NAND2xp5_ASAP7_75t_L g13173 ( 
.A(n_12509),
.B(n_833),
.Y(n_13173)
);

AOI21xp5_ASAP7_75t_L g13174 ( 
.A1(n_12223),
.A2(n_5398),
.B(n_5397),
.Y(n_13174)
);

INVx2_ASAP7_75t_L g13175 ( 
.A(n_12214),
.Y(n_13175)
);

NAND2xp5_ASAP7_75t_SL g13176 ( 
.A(n_12116),
.B(n_5400),
.Y(n_13176)
);

AO21x1_ASAP7_75t_L g13177 ( 
.A1(n_12443),
.A2(n_833),
.B(n_834),
.Y(n_13177)
);

AOI21xp5_ASAP7_75t_L g13178 ( 
.A1(n_12229),
.A2(n_5402),
.B(n_5401),
.Y(n_13178)
);

AND2x4_ASAP7_75t_L g13179 ( 
.A(n_12402),
.B(n_5403),
.Y(n_13179)
);

OAI22xp5_ASAP7_75t_L g13180 ( 
.A1(n_12664),
.A2(n_836),
.B1(n_834),
.B2(n_835),
.Y(n_13180)
);

O2A1O1Ixp5_ASAP7_75t_L g13181 ( 
.A1(n_12177),
.A2(n_837),
.B(n_835),
.C(n_836),
.Y(n_13181)
);

INVx1_ASAP7_75t_L g13182 ( 
.A(n_12358),
.Y(n_13182)
);

O2A1O1Ixp5_ASAP7_75t_L g13183 ( 
.A1(n_12060),
.A2(n_839),
.B(n_837),
.C(n_838),
.Y(n_13183)
);

BUFx6f_ASAP7_75t_L g13184 ( 
.A(n_12589),
.Y(n_13184)
);

AOI21xp5_ASAP7_75t_L g13185 ( 
.A1(n_12215),
.A2(n_5406),
.B(n_5405),
.Y(n_13185)
);

BUFx2_ASAP7_75t_L g13186 ( 
.A(n_12589),
.Y(n_13186)
);

NAND2xp5_ASAP7_75t_SL g13187 ( 
.A(n_12129),
.B(n_5407),
.Y(n_13187)
);

AOI21xp5_ASAP7_75t_L g13188 ( 
.A1(n_12280),
.A2(n_5409),
.B(n_5408),
.Y(n_13188)
);

AND2x2_ASAP7_75t_L g13189 ( 
.A(n_12619),
.B(n_838),
.Y(n_13189)
);

A2O1A1Ixp33_ASAP7_75t_L g13190 ( 
.A1(n_12102),
.A2(n_12035),
.B(n_12070),
.C(n_12011),
.Y(n_13190)
);

OAI22xp5_ASAP7_75t_L g13191 ( 
.A1(n_12674),
.A2(n_12690),
.B1(n_12694),
.B2(n_12691),
.Y(n_13191)
);

BUFx12f_ASAP7_75t_L g13192 ( 
.A(n_12205),
.Y(n_13192)
);

AO21x1_ASAP7_75t_L g13193 ( 
.A1(n_12488),
.A2(n_839),
.B(n_840),
.Y(n_13193)
);

NAND2xp5_ASAP7_75t_L g13194 ( 
.A(n_12511),
.B(n_840),
.Y(n_13194)
);

NOR2xp33_ASAP7_75t_SL g13195 ( 
.A(n_12534),
.B(n_12419),
.Y(n_13195)
);

AOI22xp33_ASAP7_75t_L g13196 ( 
.A1(n_12364),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_13196)
);

AOI22xp33_ASAP7_75t_L g13197 ( 
.A1(n_12236),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_13197)
);

AOI21xp5_ASAP7_75t_L g13198 ( 
.A1(n_12280),
.A2(n_5412),
.B(n_5410),
.Y(n_13198)
);

AOI21xp5_ASAP7_75t_L g13199 ( 
.A1(n_12174),
.A2(n_5414),
.B(n_5413),
.Y(n_13199)
);

OAI22xp5_ASAP7_75t_L g13200 ( 
.A1(n_12740),
.A2(n_846),
.B1(n_844),
.B2(n_845),
.Y(n_13200)
);

NAND2xp5_ASAP7_75t_SL g13201 ( 
.A(n_12401),
.B(n_5415),
.Y(n_13201)
);

OAI22xp5_ASAP7_75t_L g13202 ( 
.A1(n_12766),
.A2(n_847),
.B1(n_844),
.B2(n_845),
.Y(n_13202)
);

INVxp67_ASAP7_75t_L g13203 ( 
.A(n_12681),
.Y(n_13203)
);

OAI21xp5_ASAP7_75t_L g13204 ( 
.A1(n_11996),
.A2(n_5418),
.B(n_5417),
.Y(n_13204)
);

AND2x4_ASAP7_75t_L g13205 ( 
.A(n_12428),
.B(n_5419),
.Y(n_13205)
);

AOI21xp5_ASAP7_75t_L g13206 ( 
.A1(n_12176),
.A2(n_5421),
.B(n_5420),
.Y(n_13206)
);

A2O1A1Ixp33_ASAP7_75t_L g13207 ( 
.A1(n_12308),
.A2(n_851),
.B(n_848),
.C(n_849),
.Y(n_13207)
);

INVx1_ASAP7_75t_L g13208 ( 
.A(n_12372),
.Y(n_13208)
);

INVx3_ASAP7_75t_L g13209 ( 
.A(n_12589),
.Y(n_13209)
);

OAI22xp5_ASAP7_75t_SL g13210 ( 
.A1(n_12262),
.A2(n_851),
.B1(n_848),
.B2(n_849),
.Y(n_13210)
);

NOR2xp33_ASAP7_75t_L g13211 ( 
.A(n_12717),
.B(n_852),
.Y(n_13211)
);

AOI21xp5_ASAP7_75t_L g13212 ( 
.A1(n_12329),
.A2(n_5423),
.B(n_5422),
.Y(n_13212)
);

AOI22xp5_ASAP7_75t_L g13213 ( 
.A1(n_12785),
.A2(n_12791),
.B1(n_12131),
.B2(n_12186),
.Y(n_13213)
);

AND2x4_ASAP7_75t_L g13214 ( 
.A(n_12436),
.B(n_5424),
.Y(n_13214)
);

AOI21x1_ASAP7_75t_L g13215 ( 
.A1(n_12492),
.A2(n_852),
.B(n_853),
.Y(n_13215)
);

NAND2xp5_ASAP7_75t_L g13216 ( 
.A(n_12515),
.B(n_853),
.Y(n_13216)
);

NOR2xp33_ASAP7_75t_L g13217 ( 
.A(n_12726),
.B(n_854),
.Y(n_13217)
);

OAI22xp5_ASAP7_75t_L g13218 ( 
.A1(n_12362),
.A2(n_857),
.B1(n_855),
.B2(n_856),
.Y(n_13218)
);

AOI21x1_ASAP7_75t_L g13219 ( 
.A1(n_12109),
.A2(n_855),
.B(n_856),
.Y(n_13219)
);

HB1xp67_ASAP7_75t_L g13220 ( 
.A(n_12193),
.Y(n_13220)
);

NAND2xp5_ASAP7_75t_SL g13221 ( 
.A(n_12401),
.B(n_5426),
.Y(n_13221)
);

NAND2xp5_ASAP7_75t_SL g13222 ( 
.A(n_12401),
.B(n_5428),
.Y(n_13222)
);

NAND2xp5_ASAP7_75t_L g13223 ( 
.A(n_12545),
.B(n_857),
.Y(n_13223)
);

AND2x2_ASAP7_75t_L g13224 ( 
.A(n_12635),
.B(n_858),
.Y(n_13224)
);

BUFx8_ASAP7_75t_L g13225 ( 
.A(n_12344),
.Y(n_13225)
);

AOI21xp5_ASAP7_75t_L g13226 ( 
.A1(n_12513),
.A2(n_5430),
.B(n_5429),
.Y(n_13226)
);

NOR2xp33_ASAP7_75t_SL g13227 ( 
.A(n_11976),
.B(n_5431),
.Y(n_13227)
);

OR2x6_ASAP7_75t_SL g13228 ( 
.A(n_12446),
.B(n_858),
.Y(n_13228)
);

AOI21xp5_ASAP7_75t_L g13229 ( 
.A1(n_12535),
.A2(n_5433),
.B(n_5432),
.Y(n_13229)
);

NAND2xp5_ASAP7_75t_L g13230 ( 
.A(n_12557),
.B(n_12560),
.Y(n_13230)
);

AOI22xp5_ASAP7_75t_L g13231 ( 
.A1(n_12592),
.A2(n_861),
.B1(n_859),
.B2(n_860),
.Y(n_13231)
);

O2A1O1Ixp33_ASAP7_75t_L g13232 ( 
.A1(n_12684),
.A2(n_863),
.B(n_861),
.C(n_862),
.Y(n_13232)
);

INVx1_ASAP7_75t_L g13233 ( 
.A(n_12378),
.Y(n_13233)
);

NOR2xp33_ASAP7_75t_R g13234 ( 
.A(n_12283),
.B(n_5434),
.Y(n_13234)
);

NAND2xp5_ASAP7_75t_L g13235 ( 
.A(n_12562),
.B(n_862),
.Y(n_13235)
);

NAND2xp5_ASAP7_75t_L g13236 ( 
.A(n_12564),
.B(n_863),
.Y(n_13236)
);

INVxp67_ASAP7_75t_L g13237 ( 
.A(n_12772),
.Y(n_13237)
);

AOI21xp5_ASAP7_75t_L g13238 ( 
.A1(n_12452),
.A2(n_5436),
.B(n_5435),
.Y(n_13238)
);

AOI21xp5_ASAP7_75t_L g13239 ( 
.A1(n_12365),
.A2(n_5438),
.B(n_5437),
.Y(n_13239)
);

NAND2xp5_ASAP7_75t_L g13240 ( 
.A(n_12566),
.B(n_864),
.Y(n_13240)
);

NAND2xp5_ASAP7_75t_SL g13241 ( 
.A(n_12473),
.B(n_5443),
.Y(n_13241)
);

AOI21xp5_ASAP7_75t_L g13242 ( 
.A1(n_11936),
.A2(n_5447),
.B(n_5446),
.Y(n_13242)
);

AOI21xp5_ASAP7_75t_L g13243 ( 
.A1(n_12286),
.A2(n_5449),
.B(n_5448),
.Y(n_13243)
);

AOI21xp5_ASAP7_75t_L g13244 ( 
.A1(n_11945),
.A2(n_5451),
.B(n_5450),
.Y(n_13244)
);

AOI21xp5_ASAP7_75t_L g13245 ( 
.A1(n_12382),
.A2(n_5453),
.B(n_5452),
.Y(n_13245)
);

NAND3xp33_ASAP7_75t_L g13246 ( 
.A(n_12239),
.B(n_864),
.C(n_865),
.Y(n_13246)
);

INVx1_ASAP7_75t_L g13247 ( 
.A(n_12379),
.Y(n_13247)
);

INVx2_ASAP7_75t_L g13248 ( 
.A(n_12222),
.Y(n_13248)
);

AOI21xp5_ASAP7_75t_L g13249 ( 
.A1(n_11947),
.A2(n_12284),
.B(n_12321),
.Y(n_13249)
);

BUFx6f_ASAP7_75t_L g13250 ( 
.A(n_12621),
.Y(n_13250)
);

AO32x2_ASAP7_75t_L g13251 ( 
.A1(n_12461),
.A2(n_867),
.A3(n_865),
.B1(n_866),
.B2(n_868),
.Y(n_13251)
);

NOR2xp33_ASAP7_75t_L g13252 ( 
.A(n_12020),
.B(n_866),
.Y(n_13252)
);

NOR2xp33_ASAP7_75t_L g13253 ( 
.A(n_11932),
.B(n_867),
.Y(n_13253)
);

NAND2xp5_ASAP7_75t_L g13254 ( 
.A(n_12567),
.B(n_868),
.Y(n_13254)
);

OAI22xp5_ASAP7_75t_L g13255 ( 
.A1(n_12430),
.A2(n_872),
.B1(n_869),
.B2(n_871),
.Y(n_13255)
);

NAND2xp5_ASAP7_75t_SL g13256 ( 
.A(n_12399),
.B(n_12409),
.Y(n_13256)
);

A2O1A1Ixp33_ASAP7_75t_L g13257 ( 
.A1(n_12314),
.A2(n_12395),
.B(n_12729),
.C(n_12718),
.Y(n_13257)
);

NAND2xp5_ASAP7_75t_SL g13258 ( 
.A(n_12444),
.B(n_5454),
.Y(n_13258)
);

AOI21x1_ASAP7_75t_L g13259 ( 
.A1(n_12243),
.A2(n_871),
.B(n_872),
.Y(n_13259)
);

AOI21xp5_ASAP7_75t_L g13260 ( 
.A1(n_11962),
.A2(n_5456),
.B(n_5455),
.Y(n_13260)
);

AOI22xp5_ASAP7_75t_L g13261 ( 
.A1(n_12606),
.A2(n_875),
.B1(n_873),
.B2(n_874),
.Y(n_13261)
);

AOI21xp5_ASAP7_75t_L g13262 ( 
.A1(n_11963),
.A2(n_5458),
.B(n_5457),
.Y(n_13262)
);

AOI21xp5_ASAP7_75t_L g13263 ( 
.A1(n_11965),
.A2(n_5461),
.B(n_5459),
.Y(n_13263)
);

CKINVDCx5p33_ASAP7_75t_R g13264 ( 
.A(n_12240),
.Y(n_13264)
);

OAI21xp5_ASAP7_75t_L g13265 ( 
.A1(n_12533),
.A2(n_12752),
.B(n_12542),
.Y(n_13265)
);

O2A1O1Ixp33_ASAP7_75t_L g13266 ( 
.A1(n_12266),
.A2(n_875),
.B(n_873),
.C(n_874),
.Y(n_13266)
);

NAND2xp5_ASAP7_75t_L g13267 ( 
.A(n_12570),
.B(n_12573),
.Y(n_13267)
);

AOI21xp5_ASAP7_75t_L g13268 ( 
.A1(n_11971),
.A2(n_5463),
.B(n_5462),
.Y(n_13268)
);

INVx2_ASAP7_75t_L g13269 ( 
.A(n_12238),
.Y(n_13269)
);

INVx5_ASAP7_75t_L g13270 ( 
.A(n_11970),
.Y(n_13270)
);

INVx3_ASAP7_75t_L g13271 ( 
.A(n_12621),
.Y(n_13271)
);

HB1xp67_ASAP7_75t_L g13272 ( 
.A(n_12203),
.Y(n_13272)
);

AOI21xp5_ASAP7_75t_L g13273 ( 
.A1(n_11974),
.A2(n_5465),
.B(n_5464),
.Y(n_13273)
);

AOI221xp5_ASAP7_75t_L g13274 ( 
.A1(n_12440),
.A2(n_878),
.B1(n_876),
.B2(n_877),
.C(n_879),
.Y(n_13274)
);

AND2x2_ASAP7_75t_L g13275 ( 
.A(n_12640),
.B(n_878),
.Y(n_13275)
);

NAND2xp5_ASAP7_75t_L g13276 ( 
.A(n_12575),
.B(n_880),
.Y(n_13276)
);

NAND2xp5_ASAP7_75t_SL g13277 ( 
.A(n_12248),
.B(n_5467),
.Y(n_13277)
);

INVx2_ASAP7_75t_L g13278 ( 
.A(n_12245),
.Y(n_13278)
);

AND2x2_ASAP7_75t_SL g13279 ( 
.A(n_12464),
.B(n_880),
.Y(n_13279)
);

NOR2xp33_ASAP7_75t_L g13280 ( 
.A(n_11984),
.B(n_881),
.Y(n_13280)
);

OAI22xp5_ASAP7_75t_L g13281 ( 
.A1(n_12268),
.A2(n_12384),
.B1(n_12487),
.B2(n_12069),
.Y(n_13281)
);

NAND2xp5_ASAP7_75t_L g13282 ( 
.A(n_12588),
.B(n_882),
.Y(n_13282)
);

NAND2xp5_ASAP7_75t_SL g13283 ( 
.A(n_12124),
.B(n_5469),
.Y(n_13283)
);

NAND3xp33_ASAP7_75t_L g13284 ( 
.A(n_12114),
.B(n_882),
.C(n_883),
.Y(n_13284)
);

INVx3_ASAP7_75t_L g13285 ( 
.A(n_12621),
.Y(n_13285)
);

A2O1A1Ixp33_ASAP7_75t_L g13286 ( 
.A1(n_12366),
.A2(n_885),
.B(n_883),
.C(n_884),
.Y(n_13286)
);

NAND2xp5_ASAP7_75t_L g13287 ( 
.A(n_12593),
.B(n_884),
.Y(n_13287)
);

NOR2xp33_ASAP7_75t_L g13288 ( 
.A(n_12001),
.B(n_885),
.Y(n_13288)
);

NAND2xp5_ASAP7_75t_L g13289 ( 
.A(n_12599),
.B(n_886),
.Y(n_13289)
);

BUFx12f_ASAP7_75t_L g13290 ( 
.A(n_12094),
.Y(n_13290)
);

NOR2xp33_ASAP7_75t_L g13291 ( 
.A(n_12427),
.B(n_887),
.Y(n_13291)
);

NOR2xp33_ASAP7_75t_SL g13292 ( 
.A(n_12720),
.B(n_5470),
.Y(n_13292)
);

AOI21xp5_ASAP7_75t_L g13293 ( 
.A1(n_11979),
.A2(n_5474),
.B(n_5472),
.Y(n_13293)
);

BUFx3_ASAP7_75t_L g13294 ( 
.A(n_12649),
.Y(n_13294)
);

HB1xp67_ASAP7_75t_L g13295 ( 
.A(n_12204),
.Y(n_13295)
);

NAND2xp5_ASAP7_75t_L g13296 ( 
.A(n_12603),
.B(n_888),
.Y(n_13296)
);

AND2x2_ASAP7_75t_L g13297 ( 
.A(n_12642),
.B(n_888),
.Y(n_13297)
);

BUFx2_ASAP7_75t_L g13298 ( 
.A(n_12649),
.Y(n_13298)
);

NOR2xp33_ASAP7_75t_R g13299 ( 
.A(n_12324),
.B(n_5475),
.Y(n_13299)
);

AOI21xp5_ASAP7_75t_L g13300 ( 
.A1(n_11980),
.A2(n_5477),
.B(n_5476),
.Y(n_13300)
);

INVx1_ASAP7_75t_L g13301 ( 
.A(n_12381),
.Y(n_13301)
);

NAND2x1p5_ASAP7_75t_L g13302 ( 
.A(n_12004),
.B(n_5478),
.Y(n_13302)
);

INVxp67_ASAP7_75t_SL g13303 ( 
.A(n_12318),
.Y(n_13303)
);

INVxp67_ASAP7_75t_L g13304 ( 
.A(n_12649),
.Y(n_13304)
);

NAND2xp5_ASAP7_75t_SL g13305 ( 
.A(n_12403),
.B(n_5479),
.Y(n_13305)
);

AOI22xp5_ASAP7_75t_L g13306 ( 
.A1(n_12623),
.A2(n_891),
.B1(n_889),
.B2(n_890),
.Y(n_13306)
);

HB1xp67_ASAP7_75t_L g13307 ( 
.A(n_12320),
.Y(n_13307)
);

INVx1_ASAP7_75t_SL g13308 ( 
.A(n_12680),
.Y(n_13308)
);

AO22x1_ASAP7_75t_L g13309 ( 
.A1(n_12041),
.A2(n_891),
.B1(n_889),
.B2(n_890),
.Y(n_13309)
);

INVx1_ASAP7_75t_L g13310 ( 
.A(n_12386),
.Y(n_13310)
);

AOI21xp5_ASAP7_75t_L g13311 ( 
.A1(n_11982),
.A2(n_5481),
.B(n_5480),
.Y(n_13311)
);

OAI22xp5_ASAP7_75t_L g13312 ( 
.A1(n_12466),
.A2(n_894),
.B1(n_892),
.B2(n_893),
.Y(n_13312)
);

BUFx3_ASAP7_75t_L g13313 ( 
.A(n_12680),
.Y(n_13313)
);

NOR2xp33_ASAP7_75t_L g13314 ( 
.A(n_12427),
.B(n_12463),
.Y(n_13314)
);

AOI21xp5_ASAP7_75t_L g13315 ( 
.A1(n_11997),
.A2(n_12006),
.B(n_12000),
.Y(n_13315)
);

NOR2xp33_ASAP7_75t_L g13316 ( 
.A(n_12427),
.B(n_892),
.Y(n_13316)
);

NAND2xp5_ASAP7_75t_SL g13317 ( 
.A(n_11973),
.B(n_5482),
.Y(n_13317)
);

AND2x6_ASAP7_75t_L g13318 ( 
.A(n_12434),
.B(n_5483),
.Y(n_13318)
);

AOI21xp5_ASAP7_75t_L g13319 ( 
.A1(n_12009),
.A2(n_5487),
.B(n_5485),
.Y(n_13319)
);

AOI22xp33_ASAP7_75t_L g13320 ( 
.A1(n_12247),
.A2(n_896),
.B1(n_893),
.B2(n_895),
.Y(n_13320)
);

INVx2_ASAP7_75t_L g13321 ( 
.A(n_12256),
.Y(n_13321)
);

NAND2xp5_ASAP7_75t_L g13322 ( 
.A(n_12604),
.B(n_895),
.Y(n_13322)
);

AOI21xp5_ASAP7_75t_L g13323 ( 
.A1(n_12019),
.A2(n_5490),
.B(n_5488),
.Y(n_13323)
);

INVx1_ASAP7_75t_L g13324 ( 
.A(n_12258),
.Y(n_13324)
);

NAND2xp5_ASAP7_75t_L g13325 ( 
.A(n_12607),
.B(n_897),
.Y(n_13325)
);

INVx1_ASAP7_75t_L g13326 ( 
.A(n_12267),
.Y(n_13326)
);

AOI21xp5_ASAP7_75t_L g13327 ( 
.A1(n_12021),
.A2(n_5492),
.B(n_5491),
.Y(n_13327)
);

OAI22xp5_ASAP7_75t_L g13328 ( 
.A1(n_12137),
.A2(n_899),
.B1(n_897),
.B2(n_898),
.Y(n_13328)
);

AOI21xp5_ASAP7_75t_L g13329 ( 
.A1(n_12029),
.A2(n_5494),
.B(n_5493),
.Y(n_13329)
);

AOI21xp5_ASAP7_75t_L g13330 ( 
.A1(n_12033),
.A2(n_5497),
.B(n_5496),
.Y(n_13330)
);

BUFx6f_ASAP7_75t_L g13331 ( 
.A(n_12680),
.Y(n_13331)
);

NAND2xp5_ASAP7_75t_L g13332 ( 
.A(n_12609),
.B(n_898),
.Y(n_13332)
);

INVx1_ASAP7_75t_L g13333 ( 
.A(n_12269),
.Y(n_13333)
);

NOR2xp33_ASAP7_75t_L g13334 ( 
.A(n_12025),
.B(n_899),
.Y(n_13334)
);

INVx2_ASAP7_75t_L g13335 ( 
.A(n_12270),
.Y(n_13335)
);

A2O1A1Ixp33_ASAP7_75t_L g13336 ( 
.A1(n_11981),
.A2(n_902),
.B(n_900),
.C(n_901),
.Y(n_13336)
);

AOI21xp5_ASAP7_75t_L g13337 ( 
.A1(n_12038),
.A2(n_5500),
.B(n_5498),
.Y(n_13337)
);

INVx3_ASAP7_75t_L g13338 ( 
.A(n_12739),
.Y(n_13338)
);

INVx1_ASAP7_75t_L g13339 ( 
.A(n_12271),
.Y(n_13339)
);

AOI21xp5_ASAP7_75t_L g13340 ( 
.A1(n_12053),
.A2(n_5502),
.B(n_5501),
.Y(n_13340)
);

NOR2xp33_ASAP7_75t_L g13341 ( 
.A(n_12346),
.B(n_900),
.Y(n_13341)
);

A2O1A1Ixp33_ASAP7_75t_L g13342 ( 
.A1(n_12046),
.A2(n_905),
.B(n_902),
.C(n_904),
.Y(n_13342)
);

AOI21xp5_ASAP7_75t_L g13343 ( 
.A1(n_12055),
.A2(n_12062),
.B(n_12058),
.Y(n_13343)
);

AOI21xp5_ASAP7_75t_L g13344 ( 
.A1(n_12083),
.A2(n_5504),
.B(n_5503),
.Y(n_13344)
);

INVx2_ASAP7_75t_L g13345 ( 
.A(n_12272),
.Y(n_13345)
);

AOI21xp5_ASAP7_75t_L g13346 ( 
.A1(n_12084),
.A2(n_5506),
.B(n_5505),
.Y(n_13346)
);

AOI21xp5_ASAP7_75t_L g13347 ( 
.A1(n_12085),
.A2(n_5508),
.B(n_5507),
.Y(n_13347)
);

O2A1O1Ixp33_ASAP7_75t_L g13348 ( 
.A1(n_12057),
.A2(n_906),
.B(n_904),
.C(n_905),
.Y(n_13348)
);

AOI21xp5_ASAP7_75t_L g13349 ( 
.A1(n_12086),
.A2(n_5510),
.B(n_5509),
.Y(n_13349)
);

A2O1A1Ixp33_ASAP7_75t_L g13350 ( 
.A1(n_12759),
.A2(n_908),
.B(n_906),
.C(n_907),
.Y(n_13350)
);

AOI21xp5_ASAP7_75t_L g13351 ( 
.A1(n_12087),
.A2(n_5513),
.B(n_5512),
.Y(n_13351)
);

NAND2xp5_ASAP7_75t_L g13352 ( 
.A(n_12617),
.B(n_907),
.Y(n_13352)
);

NOR3xp33_ASAP7_75t_L g13353 ( 
.A(n_12297),
.B(n_908),
.C(n_909),
.Y(n_13353)
);

INVx2_ASAP7_75t_L g13354 ( 
.A(n_12274),
.Y(n_13354)
);

NOR2xp33_ASAP7_75t_L g13355 ( 
.A(n_12115),
.B(n_910),
.Y(n_13355)
);

INVxp67_ASAP7_75t_L g13356 ( 
.A(n_12739),
.Y(n_13356)
);

AOI22xp5_ASAP7_75t_L g13357 ( 
.A1(n_12689),
.A2(n_12700),
.B1(n_12773),
.B2(n_12709),
.Y(n_13357)
);

AO21x2_ASAP7_75t_L g13358 ( 
.A1(n_12253),
.A2(n_910),
.B(n_911),
.Y(n_13358)
);

AND2x2_ASAP7_75t_L g13359 ( 
.A(n_12652),
.B(n_911),
.Y(n_13359)
);

NAND3xp33_ASAP7_75t_L g13360 ( 
.A(n_12175),
.B(n_912),
.C(n_913),
.Y(n_13360)
);

O2A1O1Ixp33_ASAP7_75t_L g13361 ( 
.A1(n_12059),
.A2(n_914),
.B(n_912),
.C(n_913),
.Y(n_13361)
);

AOI21xp5_ASAP7_75t_L g13362 ( 
.A1(n_12090),
.A2(n_5516),
.B(n_5515),
.Y(n_13362)
);

NAND2xp5_ASAP7_75t_SL g13363 ( 
.A(n_12184),
.B(n_5517),
.Y(n_13363)
);

INVx1_ASAP7_75t_L g13364 ( 
.A(n_12292),
.Y(n_13364)
);

BUFx8_ASAP7_75t_SL g13365 ( 
.A(n_12519),
.Y(n_13365)
);

NAND2xp5_ASAP7_75t_L g13366 ( 
.A(n_12618),
.B(n_915),
.Y(n_13366)
);

NAND2xp5_ASAP7_75t_L g13367 ( 
.A(n_12625),
.B(n_915),
.Y(n_13367)
);

NAND2xp5_ASAP7_75t_SL g13368 ( 
.A(n_12208),
.B(n_5518),
.Y(n_13368)
);

INVx2_ASAP7_75t_L g13369 ( 
.A(n_12295),
.Y(n_13369)
);

BUFx12f_ASAP7_75t_L g13370 ( 
.A(n_12192),
.Y(n_13370)
);

NOR2xp33_ASAP7_75t_L g13371 ( 
.A(n_12259),
.B(n_916),
.Y(n_13371)
);

NOR2xp33_ASAP7_75t_L g13372 ( 
.A(n_12278),
.B(n_917),
.Y(n_13372)
);

OAI21xp5_ASAP7_75t_L g13373 ( 
.A1(n_12146),
.A2(n_5521),
.B(n_5520),
.Y(n_13373)
);

OAI22xp5_ASAP7_75t_L g13374 ( 
.A1(n_12064),
.A2(n_11957),
.B1(n_12433),
.B2(n_12148),
.Y(n_13374)
);

OAI22xp5_ASAP7_75t_L g13375 ( 
.A1(n_12134),
.A2(n_919),
.B1(n_917),
.B2(n_918),
.Y(n_13375)
);

CKINVDCx5p33_ASAP7_75t_R g13376 ( 
.A(n_12778),
.Y(n_13376)
);

BUFx2_ASAP7_75t_L g13377 ( 
.A(n_12739),
.Y(n_13377)
);

NAND2x1p5_ASAP7_75t_L g13378 ( 
.A(n_12422),
.B(n_5523),
.Y(n_13378)
);

AOI21xp5_ASAP7_75t_L g13379 ( 
.A1(n_12092),
.A2(n_5525),
.B(n_5524),
.Y(n_13379)
);

AOI21xp5_ASAP7_75t_L g13380 ( 
.A1(n_12052),
.A2(n_5527),
.B(n_5526),
.Y(n_13380)
);

OAI21xp5_ASAP7_75t_L g13381 ( 
.A1(n_12230),
.A2(n_5529),
.B(n_5528),
.Y(n_13381)
);

NAND2xp5_ASAP7_75t_L g13382 ( 
.A(n_12629),
.B(n_918),
.Y(n_13382)
);

OAI22xp5_ASAP7_75t_L g13383 ( 
.A1(n_12149),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.Y(n_13383)
);

NAND3xp33_ASAP7_75t_L g13384 ( 
.A(n_12172),
.B(n_920),
.C(n_921),
.Y(n_13384)
);

AOI22xp5_ASAP7_75t_L g13385 ( 
.A1(n_12107),
.A2(n_926),
.B1(n_923),
.B2(n_925),
.Y(n_13385)
);

CKINVDCx8_ASAP7_75t_R g13386 ( 
.A(n_12335),
.Y(n_13386)
);

NAND2xp5_ASAP7_75t_L g13387 ( 
.A(n_12633),
.B(n_923),
.Y(n_13387)
);

BUFx12f_ASAP7_75t_L g13388 ( 
.A(n_12313),
.Y(n_13388)
);

NAND2xp5_ASAP7_75t_L g13389 ( 
.A(n_12637),
.B(n_925),
.Y(n_13389)
);

AOI22xp33_ASAP7_75t_SL g13390 ( 
.A1(n_12483),
.A2(n_928),
.B1(n_926),
.B2(n_927),
.Y(n_13390)
);

INVx1_ASAP7_75t_L g13391 ( 
.A(n_12296),
.Y(n_13391)
);

INVx2_ASAP7_75t_SL g13392 ( 
.A(n_12299),
.Y(n_13392)
);

INVx1_ASAP7_75t_L g13393 ( 
.A(n_12310),
.Y(n_13393)
);

AOI21xp5_ASAP7_75t_L g13394 ( 
.A1(n_12071),
.A2(n_5533),
.B(n_5530),
.Y(n_13394)
);

INVx5_ASAP7_75t_L g13395 ( 
.A(n_12299),
.Y(n_13395)
);

A2O1A1Ixp33_ASAP7_75t_L g13396 ( 
.A1(n_12328),
.A2(n_929),
.B(n_927),
.C(n_928),
.Y(n_13396)
);

AOI21xp5_ASAP7_75t_L g13397 ( 
.A1(n_12096),
.A2(n_5535),
.B(n_5534),
.Y(n_13397)
);

AO21x1_ASAP7_75t_L g13398 ( 
.A1(n_12334),
.A2(n_929),
.B(n_930),
.Y(n_13398)
);

AOI21xp5_ASAP7_75t_L g13399 ( 
.A1(n_12147),
.A2(n_12154),
.B(n_11987),
.Y(n_13399)
);

NAND2xp5_ASAP7_75t_L g13400 ( 
.A(n_12643),
.B(n_930),
.Y(n_13400)
);

CKINVDCx11_ASAP7_75t_R g13401 ( 
.A(n_12648),
.Y(n_13401)
);

NAND2xp5_ASAP7_75t_L g13402 ( 
.A(n_12651),
.B(n_931),
.Y(n_13402)
);

NAND2xp5_ASAP7_75t_L g13403 ( 
.A(n_12661),
.B(n_932),
.Y(n_13403)
);

AOI21xp5_ASAP7_75t_L g13404 ( 
.A1(n_11977),
.A2(n_5537),
.B(n_5536),
.Y(n_13404)
);

OAI21xp5_ASAP7_75t_L g13405 ( 
.A1(n_12183),
.A2(n_5541),
.B(n_5539),
.Y(n_13405)
);

OAI21x1_ASAP7_75t_L g13406 ( 
.A1(n_12319),
.A2(n_5545),
.B(n_5544),
.Y(n_13406)
);

NAND2xp5_ASAP7_75t_L g13407 ( 
.A(n_12666),
.B(n_932),
.Y(n_13407)
);

BUFx6f_ASAP7_75t_L g13408 ( 
.A(n_12299),
.Y(n_13408)
);

A2O1A1Ixp33_ASAP7_75t_L g13409 ( 
.A1(n_12342),
.A2(n_935),
.B(n_933),
.C(n_934),
.Y(n_13409)
);

INVx5_ASAP7_75t_L g13410 ( 
.A(n_12450),
.Y(n_13410)
);

AOI22xp5_ASAP7_75t_L g13411 ( 
.A1(n_12279),
.A2(n_935),
.B1(n_933),
.B2(n_934),
.Y(n_13411)
);

NOR2xp33_ASAP7_75t_L g13412 ( 
.A(n_12171),
.B(n_936),
.Y(n_13412)
);

AOI22xp5_ASAP7_75t_L g13413 ( 
.A1(n_12307),
.A2(n_938),
.B1(n_936),
.B2(n_937),
.Y(n_13413)
);

OAI22xp5_ASAP7_75t_L g13414 ( 
.A1(n_12206),
.A2(n_939),
.B1(n_937),
.B2(n_938),
.Y(n_13414)
);

NAND2xp5_ASAP7_75t_L g13415 ( 
.A(n_12671),
.B(n_939),
.Y(n_13415)
);

OAI22xp5_ASAP7_75t_L g13416 ( 
.A1(n_12219),
.A2(n_942),
.B1(n_940),
.B2(n_941),
.Y(n_13416)
);

AOI21xp5_ASAP7_75t_L g13417 ( 
.A1(n_11992),
.A2(n_5548),
.B(n_5547),
.Y(n_13417)
);

O2A1O1Ixp33_ASAP7_75t_L g13418 ( 
.A1(n_12036),
.A2(n_944),
.B(n_940),
.C(n_943),
.Y(n_13418)
);

OAI22xp5_ASAP7_75t_L g13419 ( 
.A1(n_12414),
.A2(n_945),
.B1(n_943),
.B2(n_944),
.Y(n_13419)
);

OAI22xp5_ASAP7_75t_L g13420 ( 
.A1(n_12294),
.A2(n_947),
.B1(n_945),
.B2(n_946),
.Y(n_13420)
);

NOR2xp33_ASAP7_75t_L g13421 ( 
.A(n_12202),
.B(n_946),
.Y(n_13421)
);

INVx1_ASAP7_75t_L g13422 ( 
.A(n_12201),
.Y(n_13422)
);

AND2x4_ASAP7_75t_L g13423 ( 
.A(n_12447),
.B(n_5549),
.Y(n_13423)
);

AND2x4_ASAP7_75t_L g13424 ( 
.A(n_11960),
.B(n_5550),
.Y(n_13424)
);

AOI21x1_ASAP7_75t_L g13425 ( 
.A1(n_12264),
.A2(n_948),
.B(n_949),
.Y(n_13425)
);

AO22x1_ASAP7_75t_L g13426 ( 
.A1(n_12441),
.A2(n_950),
.B1(n_948),
.B2(n_949),
.Y(n_13426)
);

INVx1_ASAP7_75t_L g13427 ( 
.A(n_12453),
.Y(n_13427)
);

NAND2xp5_ASAP7_75t_SL g13428 ( 
.A(n_12218),
.B(n_5551),
.Y(n_13428)
);

O2A1O1Ixp33_ASAP7_75t_L g13429 ( 
.A1(n_12018),
.A2(n_952),
.B(n_950),
.C(n_951),
.Y(n_13429)
);

INVx3_ASAP7_75t_L g13430 ( 
.A(n_12787),
.Y(n_13430)
);

BUFx6f_ASAP7_75t_L g13431 ( 
.A(n_12595),
.Y(n_13431)
);

BUFx6f_ASAP7_75t_L g13432 ( 
.A(n_12728),
.Y(n_13432)
);

NAND2xp5_ASAP7_75t_L g13433 ( 
.A(n_12675),
.B(n_952),
.Y(n_13433)
);

INVx3_ASAP7_75t_L g13434 ( 
.A(n_12596),
.Y(n_13434)
);

AOI21xp5_ASAP7_75t_L g13435 ( 
.A1(n_12241),
.A2(n_5553),
.B(n_5552),
.Y(n_13435)
);

AOI21xp5_ASAP7_75t_L g13436 ( 
.A1(n_12251),
.A2(n_5556),
.B(n_5554),
.Y(n_13436)
);

NOR2xp67_ASAP7_75t_SL g13437 ( 
.A(n_12539),
.B(n_5557),
.Y(n_13437)
);

INVx1_ASAP7_75t_L g13438 ( 
.A(n_12453),
.Y(n_13438)
);

INVxp33_ASAP7_75t_SL g13439 ( 
.A(n_12332),
.Y(n_13439)
);

AND2x4_ASAP7_75t_L g13440 ( 
.A(n_12613),
.B(n_5558),
.Y(n_13440)
);

NOR2xp33_ASAP7_75t_L g13441 ( 
.A(n_12705),
.B(n_953),
.Y(n_13441)
);

AOI21xp5_ASAP7_75t_L g13442 ( 
.A1(n_12287),
.A2(n_5560),
.B(n_5559),
.Y(n_13442)
);

NOR2xp33_ASAP7_75t_L g13443 ( 
.A(n_12737),
.B(n_953),
.Y(n_13443)
);

OA22x2_ASAP7_75t_L g13444 ( 
.A1(n_12456),
.A2(n_956),
.B1(n_954),
.B2(n_955),
.Y(n_13444)
);

INVx2_ASAP7_75t_L g13445 ( 
.A(n_12336),
.Y(n_13445)
);

NAND2xp5_ASAP7_75t_L g13446 ( 
.A(n_12682),
.B(n_955),
.Y(n_13446)
);

NAND2xp5_ASAP7_75t_SL g13447 ( 
.A(n_12322),
.B(n_5561),
.Y(n_13447)
);

A2O1A1Ixp33_ASAP7_75t_L g13448 ( 
.A1(n_12470),
.A2(n_959),
.B(n_957),
.C(n_958),
.Y(n_13448)
);

NAND2xp5_ASAP7_75t_L g13449 ( 
.A(n_12701),
.B(n_957),
.Y(n_13449)
);

OR2x6_ASAP7_75t_SL g13450 ( 
.A(n_12457),
.B(n_12462),
.Y(n_13450)
);

NAND2xp5_ASAP7_75t_L g13451 ( 
.A(n_12703),
.B(n_958),
.Y(n_13451)
);

OAI21xp5_ASAP7_75t_L g13452 ( 
.A1(n_12338),
.A2(n_12133),
.B(n_12132),
.Y(n_13452)
);

NOR2xp33_ASAP7_75t_L g13453 ( 
.A(n_12757),
.B(n_959),
.Y(n_13453)
);

BUFx2_ASAP7_75t_L g13454 ( 
.A(n_12254),
.Y(n_13454)
);

INVx2_ASAP7_75t_L g13455 ( 
.A(n_12421),
.Y(n_13455)
);

HB1xp67_ASAP7_75t_L g13456 ( 
.A(n_12465),
.Y(n_13456)
);

OAI22xp5_ASAP7_75t_L g13457 ( 
.A1(n_12165),
.A2(n_962),
.B1(n_960),
.B2(n_961),
.Y(n_13457)
);

INVx2_ASAP7_75t_L g13458 ( 
.A(n_12108),
.Y(n_13458)
);

AOI22xp33_ASAP7_75t_L g13459 ( 
.A1(n_12054),
.A2(n_962),
.B1(n_960),
.B2(n_961),
.Y(n_13459)
);

NAND2xp5_ASAP7_75t_SL g13460 ( 
.A(n_12347),
.B(n_5562),
.Y(n_13460)
);

NAND2xp5_ASAP7_75t_SL g13461 ( 
.A(n_12349),
.B(n_5563),
.Y(n_13461)
);

A2O1A1Ixp33_ASAP7_75t_L g13462 ( 
.A1(n_12276),
.A2(n_965),
.B(n_963),
.C(n_964),
.Y(n_13462)
);

OAI22xp5_ASAP7_75t_L g13463 ( 
.A1(n_12708),
.A2(n_966),
.B1(n_963),
.B2(n_965),
.Y(n_13463)
);

OAI22xp5_ASAP7_75t_L g13464 ( 
.A1(n_12723),
.A2(n_968),
.B1(n_966),
.B2(n_967),
.Y(n_13464)
);

OAI22xp5_ASAP7_75t_L g13465 ( 
.A1(n_12735),
.A2(n_969),
.B1(n_967),
.B2(n_968),
.Y(n_13465)
);

NAND2xp5_ASAP7_75t_L g13466 ( 
.A(n_12743),
.B(n_969),
.Y(n_13466)
);

AOI21xp5_ASAP7_75t_L g13467 ( 
.A1(n_12291),
.A2(n_5566),
.B(n_5565),
.Y(n_13467)
);

AOI33xp33_ASAP7_75t_L g13468 ( 
.A1(n_12490),
.A2(n_972),
.A3(n_974),
.B1(n_970),
.B2(n_971),
.B3(n_973),
.Y(n_13468)
);

AOI21xp5_ASAP7_75t_L g13469 ( 
.A1(n_12300),
.A2(n_5568),
.B(n_5567),
.Y(n_13469)
);

INVx3_ASAP7_75t_L g13470 ( 
.A(n_12656),
.Y(n_13470)
);

NAND2xp5_ASAP7_75t_SL g13471 ( 
.A(n_12484),
.B(n_5569),
.Y(n_13471)
);

AOI21xp5_ASAP7_75t_L g13472 ( 
.A1(n_12306),
.A2(n_5576),
.B(n_5574),
.Y(n_13472)
);

AND2x2_ASAP7_75t_L g13473 ( 
.A(n_12765),
.B(n_972),
.Y(n_13473)
);

NAND2xp5_ASAP7_75t_L g13474 ( 
.A(n_12746),
.B(n_12751),
.Y(n_13474)
);

AOI21xp5_ASAP7_75t_L g13475 ( 
.A1(n_12135),
.A2(n_5578),
.B(n_5577),
.Y(n_13475)
);

NOR2xp33_ASAP7_75t_L g13476 ( 
.A(n_12789),
.B(n_973),
.Y(n_13476)
);

BUFx6f_ASAP7_75t_L g13477 ( 
.A(n_12361),
.Y(n_13477)
);

INVx3_ASAP7_75t_L g13478 ( 
.A(n_12160),
.Y(n_13478)
);

AND2x2_ASAP7_75t_L g13479 ( 
.A(n_12091),
.B(n_974),
.Y(n_13479)
);

NAND2xp5_ASAP7_75t_L g13480 ( 
.A(n_12753),
.B(n_12755),
.Y(n_13480)
);

NAND2xp5_ASAP7_75t_SL g13481 ( 
.A(n_12486),
.B(n_5579),
.Y(n_13481)
);

AOI21xp5_ASAP7_75t_L g13482 ( 
.A1(n_12136),
.A2(n_12143),
.B(n_12141),
.Y(n_13482)
);

NAND3xp33_ASAP7_75t_L g13483 ( 
.A(n_12489),
.B(n_975),
.C(n_976),
.Y(n_13483)
);

AOI21xp5_ASAP7_75t_L g13484 ( 
.A1(n_12161),
.A2(n_5581),
.B(n_5580),
.Y(n_13484)
);

AOI21xp5_ASAP7_75t_L g13485 ( 
.A1(n_12330),
.A2(n_5583),
.B(n_5582),
.Y(n_13485)
);

AOI21xp5_ASAP7_75t_L g13486 ( 
.A1(n_12406),
.A2(n_5585),
.B(n_5584),
.Y(n_13486)
);

OR2x2_ASAP7_75t_L g13487 ( 
.A(n_12415),
.B(n_975),
.Y(n_13487)
);

INVx1_ASAP7_75t_L g13488 ( 
.A(n_12453),
.Y(n_13488)
);

NAND2xp5_ASAP7_75t_L g13489 ( 
.A(n_12756),
.B(n_976),
.Y(n_13489)
);

BUFx2_ASAP7_75t_L g13490 ( 
.A(n_12376),
.Y(n_13490)
);

NOR2xp33_ASAP7_75t_L g13491 ( 
.A(n_12408),
.B(n_977),
.Y(n_13491)
);

NAND2xp5_ASAP7_75t_SL g13492 ( 
.A(n_12425),
.B(n_5586),
.Y(n_13492)
);

AOI21xp5_ASAP7_75t_L g13493 ( 
.A1(n_12416),
.A2(n_5588),
.B(n_5587),
.Y(n_13493)
);

BUFx6f_ASAP7_75t_L g13494 ( 
.A(n_12343),
.Y(n_13494)
);

A2O1A1Ixp33_ASAP7_75t_L g13495 ( 
.A1(n_12579),
.A2(n_979),
.B(n_977),
.C(n_978),
.Y(n_13495)
);

NAND2xp5_ASAP7_75t_L g13496 ( 
.A(n_12762),
.B(n_978),
.Y(n_13496)
);

NAND2xp5_ASAP7_75t_L g13497 ( 
.A(n_12763),
.B(n_979),
.Y(n_13497)
);

NAND2xp5_ASAP7_75t_L g13498 ( 
.A(n_12764),
.B(n_980),
.Y(n_13498)
);

INVx1_ASAP7_75t_L g13499 ( 
.A(n_11998),
.Y(n_13499)
);

NAND2x1p5_ASAP7_75t_L g13500 ( 
.A(n_11972),
.B(n_5589),
.Y(n_13500)
);

NAND2xp5_ASAP7_75t_L g13501 ( 
.A(n_12767),
.B(n_980),
.Y(n_13501)
);

OAI22xp5_ASAP7_75t_L g13502 ( 
.A1(n_12774),
.A2(n_983),
.B1(n_981),
.B2(n_982),
.Y(n_13502)
);

NAND2xp5_ASAP7_75t_SL g13503 ( 
.A(n_12496),
.B(n_5590),
.Y(n_13503)
);

AOI21xp5_ASAP7_75t_L g13504 ( 
.A1(n_12417),
.A2(n_5592),
.B(n_5591),
.Y(n_13504)
);

INVx3_ASAP7_75t_SL g13505 ( 
.A(n_12056),
.Y(n_13505)
);

NAND2xp5_ASAP7_75t_SL g13506 ( 
.A(n_12468),
.B(n_5594),
.Y(n_13506)
);

AOI21xp5_ASAP7_75t_L g13507 ( 
.A1(n_12420),
.A2(n_5597),
.B(n_5595),
.Y(n_13507)
);

NAND2xp5_ASAP7_75t_L g13508 ( 
.A(n_12022),
.B(n_981),
.Y(n_13508)
);

AOI21xp5_ASAP7_75t_L g13509 ( 
.A1(n_12439),
.A2(n_5599),
.B(n_5598),
.Y(n_13509)
);

NAND2xp5_ASAP7_75t_L g13510 ( 
.A(n_12027),
.B(n_12031),
.Y(n_13510)
);

A2O1A1Ixp33_ASAP7_75t_L g13511 ( 
.A1(n_12732),
.A2(n_984),
.B(n_982),
.C(n_983),
.Y(n_13511)
);

AOI21xp5_ASAP7_75t_L g13512 ( 
.A1(n_12130),
.A2(n_5601),
.B(n_5600),
.Y(n_13512)
);

NOR2xp33_ASAP7_75t_L g13513 ( 
.A(n_12100),
.B(n_984),
.Y(n_13513)
);

NAND2xp5_ASAP7_75t_L g13514 ( 
.A(n_12061),
.B(n_985),
.Y(n_13514)
);

AOI21xp5_ASAP7_75t_L g13515 ( 
.A1(n_12311),
.A2(n_5603),
.B(n_5602),
.Y(n_13515)
);

O2A1O1Ixp33_ASAP7_75t_L g13516 ( 
.A1(n_12028),
.A2(n_987),
.B(n_985),
.C(n_986),
.Y(n_13516)
);

OR2x6_ASAP7_75t_L g13517 ( 
.A(n_12476),
.B(n_5604),
.Y(n_13517)
);

AOI22xp33_ASAP7_75t_L g13518 ( 
.A1(n_12110),
.A2(n_988),
.B1(n_986),
.B2(n_987),
.Y(n_13518)
);

OAI22xp5_ASAP7_75t_L g13519 ( 
.A1(n_12039),
.A2(n_990),
.B1(n_988),
.B2(n_989),
.Y(n_13519)
);

NOR2xp67_ASAP7_75t_L g13520 ( 
.A(n_11951),
.B(n_11954),
.Y(n_13520)
);

OAI22xp5_ASAP7_75t_L g13521 ( 
.A1(n_12469),
.A2(n_993),
.B1(n_989),
.B2(n_992),
.Y(n_13521)
);

AO21x1_ASAP7_75t_L g13522 ( 
.A1(n_12157),
.A2(n_993),
.B(n_994),
.Y(n_13522)
);

AOI21xp5_ASAP7_75t_L g13523 ( 
.A1(n_12371),
.A2(n_5607),
.B(n_5606),
.Y(n_13523)
);

NAND2xp5_ASAP7_75t_SL g13524 ( 
.A(n_11994),
.B(n_5609),
.Y(n_13524)
);

INVx2_ASAP7_75t_SL g13525 ( 
.A(n_12103),
.Y(n_13525)
);

AOI21xp5_ASAP7_75t_L g13526 ( 
.A1(n_12459),
.A2(n_5614),
.B(n_5612),
.Y(n_13526)
);

AND2x2_ASAP7_75t_L g13527 ( 
.A(n_12217),
.B(n_994),
.Y(n_13527)
);

NAND2xp5_ASAP7_75t_L g13528 ( 
.A(n_12065),
.B(n_995),
.Y(n_13528)
);

NAND2x1p5_ASAP7_75t_L g13529 ( 
.A(n_12678),
.B(n_5616),
.Y(n_13529)
);

INVx2_ASAP7_75t_L g13530 ( 
.A(n_12163),
.Y(n_13530)
);

OAI22xp5_ASAP7_75t_L g13531 ( 
.A1(n_12478),
.A2(n_998),
.B1(n_995),
.B2(n_996),
.Y(n_13531)
);

AOI21xp5_ASAP7_75t_L g13532 ( 
.A1(n_12354),
.A2(n_5619),
.B(n_5618),
.Y(n_13532)
);

AOI22xp5_ASAP7_75t_L g13533 ( 
.A1(n_12458),
.A2(n_1000),
.B1(n_996),
.B2(n_999),
.Y(n_13533)
);

AOI21xp5_ASAP7_75t_L g13534 ( 
.A1(n_12360),
.A2(n_5622),
.B(n_5621),
.Y(n_13534)
);

OAI22xp5_ASAP7_75t_L g13535 ( 
.A1(n_12067),
.A2(n_1002),
.B1(n_999),
.B2(n_1001),
.Y(n_13535)
);

NAND2xp5_ASAP7_75t_L g13536 ( 
.A(n_12076),
.B(n_1001),
.Y(n_13536)
);

NOR2xp67_ASAP7_75t_L g13537 ( 
.A(n_11961),
.B(n_1002),
.Y(n_13537)
);

INVx2_ASAP7_75t_L g13538 ( 
.A(n_12077),
.Y(n_13538)
);

INVxp67_ASAP7_75t_L g13539 ( 
.A(n_11978),
.Y(n_13539)
);

OAI22xp5_ASAP7_75t_L g13540 ( 
.A1(n_12078),
.A2(n_1005),
.B1(n_1003),
.B2(n_1004),
.Y(n_13540)
);

NOR2xp33_ASAP7_75t_L g13541 ( 
.A(n_12233),
.B(n_1003),
.Y(n_13541)
);

NAND2xp5_ASAP7_75t_L g13542 ( 
.A(n_12081),
.B(n_1004),
.Y(n_13542)
);

INVx2_ASAP7_75t_L g13543 ( 
.A(n_12093),
.Y(n_13543)
);

NOR2xp33_ASAP7_75t_L g13544 ( 
.A(n_12290),
.B(n_1005),
.Y(n_13544)
);

AOI22xp5_ASAP7_75t_L g13545 ( 
.A1(n_12437),
.A2(n_1008),
.B1(n_1006),
.B2(n_1007),
.Y(n_13545)
);

NAND2xp5_ASAP7_75t_L g13546 ( 
.A(n_12112),
.B(n_1006),
.Y(n_13546)
);

INVx2_ASAP7_75t_L g13547 ( 
.A(n_12391),
.Y(n_13547)
);

O2A1O1Ixp33_ASAP7_75t_SL g13548 ( 
.A1(n_12111),
.A2(n_1010),
.B(n_1007),
.C(n_1009),
.Y(n_13548)
);

NAND2xp5_ASAP7_75t_L g13549 ( 
.A(n_12123),
.B(n_1009),
.Y(n_13549)
);

AOI22xp5_ASAP7_75t_L g13550 ( 
.A1(n_12442),
.A2(n_1013),
.B1(n_1011),
.B2(n_1012),
.Y(n_13550)
);

A2O1A1Ixp33_ASAP7_75t_L g13551 ( 
.A1(n_12158),
.A2(n_1014),
.B(n_1011),
.C(n_1013),
.Y(n_13551)
);

BUFx6f_ASAP7_75t_L g13552 ( 
.A(n_12150),
.Y(n_13552)
);

NAND2xp5_ASAP7_75t_SL g13553 ( 
.A(n_12333),
.B(n_5623),
.Y(n_13553)
);

AOI21xp5_ASAP7_75t_L g13554 ( 
.A1(n_12370),
.A2(n_5626),
.B(n_5625),
.Y(n_13554)
);

INVx1_ASAP7_75t_L g13555 ( 
.A(n_12125),
.Y(n_13555)
);

INVx2_ASAP7_75t_L g13556 ( 
.A(n_12127),
.Y(n_13556)
);

INVx2_ASAP7_75t_L g13557 ( 
.A(n_12138),
.Y(n_13557)
);

OAI21xp5_ASAP7_75t_L g13558 ( 
.A1(n_12387),
.A2(n_5628),
.B(n_5627),
.Y(n_13558)
);

NAND2xp5_ASAP7_75t_L g13559 ( 
.A(n_12140),
.B(n_1014),
.Y(n_13559)
);

NAND2xp5_ASAP7_75t_L g13560 ( 
.A(n_12145),
.B(n_1015),
.Y(n_13560)
);

NAND2xp5_ASAP7_75t_SL g13561 ( 
.A(n_12181),
.B(n_5629),
.Y(n_13561)
);

NOR2xp33_ASAP7_75t_L g13562 ( 
.A(n_12359),
.B(n_1015),
.Y(n_13562)
);

OR2x6_ASAP7_75t_SL g13563 ( 
.A(n_11989),
.B(n_1016),
.Y(n_13563)
);

INVx1_ASAP7_75t_SL g13564 ( 
.A(n_12393),
.Y(n_13564)
);

INVx1_ASAP7_75t_L g13565 ( 
.A(n_12151),
.Y(n_13565)
);

NAND2xp5_ASAP7_75t_L g13566 ( 
.A(n_12339),
.B(n_1016),
.Y(n_13566)
);

BUFx4f_ASAP7_75t_L g13567 ( 
.A(n_12367),
.Y(n_13567)
);

AOI21xp5_ASAP7_75t_L g13568 ( 
.A1(n_12212),
.A2(n_5633),
.B(n_5631),
.Y(n_13568)
);

AO21x1_ASAP7_75t_L g13569 ( 
.A1(n_12106),
.A2(n_1017),
.B(n_1018),
.Y(n_13569)
);

INVx2_ASAP7_75t_SL g13570 ( 
.A(n_12228),
.Y(n_13570)
);

HB1xp67_ASAP7_75t_L g13571 ( 
.A(n_12405),
.Y(n_13571)
);

OR2x2_ASAP7_75t_L g13572 ( 
.A(n_12352),
.B(n_1017),
.Y(n_13572)
);

OAI22xp5_ASAP7_75t_L g13573 ( 
.A1(n_12474),
.A2(n_1020),
.B1(n_1018),
.B2(n_1019),
.Y(n_13573)
);

O2A1O1Ixp33_ASAP7_75t_L g13574 ( 
.A1(n_12180),
.A2(n_1021),
.B(n_1019),
.C(n_1020),
.Y(n_13574)
);

AOI21xp5_ASAP7_75t_L g13575 ( 
.A1(n_12216),
.A2(n_5635),
.B(n_5634),
.Y(n_13575)
);

OAI22xp5_ASAP7_75t_L g13576 ( 
.A1(n_12460),
.A2(n_1024),
.B1(n_1022),
.B2(n_1023),
.Y(n_13576)
);

INVx1_ASAP7_75t_L g13577 ( 
.A(n_11941),
.Y(n_13577)
);

AND2x2_ASAP7_75t_L g13578 ( 
.A(n_12418),
.B(n_1022),
.Y(n_13578)
);

OAI22xp5_ASAP7_75t_L g13579 ( 
.A1(n_12477),
.A2(n_12117),
.B1(n_12182),
.B2(n_12220),
.Y(n_13579)
);

NAND2xp5_ASAP7_75t_SL g13580 ( 
.A(n_12448),
.B(n_5636),
.Y(n_13580)
);

AOI21xp5_ASAP7_75t_L g13581 ( 
.A1(n_12190),
.A2(n_5638),
.B(n_5637),
.Y(n_13581)
);

NOR2xp67_ASAP7_75t_L g13582 ( 
.A(n_12195),
.B(n_1024),
.Y(n_13582)
);

OAI22xp5_ASAP7_75t_L g13583 ( 
.A1(n_12196),
.A2(n_1027),
.B1(n_1025),
.B2(n_1026),
.Y(n_13583)
);

AOI21xp5_ASAP7_75t_L g13584 ( 
.A1(n_12790),
.A2(n_5640),
.B(n_5639),
.Y(n_13584)
);

AOI21xp5_ASAP7_75t_L g13585 ( 
.A1(n_12099),
.A2(n_5642),
.B(n_5641),
.Y(n_13585)
);

CKINVDCx11_ASAP7_75t_R g13586 ( 
.A(n_12227),
.Y(n_13586)
);

NOR2xp33_ASAP7_75t_L g13587 ( 
.A(n_12169),
.B(n_1026),
.Y(n_13587)
);

AOI21xp5_ASAP7_75t_L g13588 ( 
.A1(n_12634),
.A2(n_5644),
.B(n_5643),
.Y(n_13588)
);

AOI21xp5_ASAP7_75t_L g13589 ( 
.A1(n_11941),
.A2(n_12731),
.B(n_12636),
.Y(n_13589)
);

AOI22xp5_ASAP7_75t_L g13590 ( 
.A1(n_11941),
.A2(n_1029),
.B1(n_1027),
.B2(n_1028),
.Y(n_13590)
);

AO21x2_ASAP7_75t_L g13591 ( 
.A1(n_12024),
.A2(n_1029),
.B(n_1030),
.Y(n_13591)
);

OAI22xp5_ASAP7_75t_L g13592 ( 
.A1(n_12731),
.A2(n_12119),
.B1(n_1032),
.B2(n_1030),
.Y(n_13592)
);

INVx2_ASAP7_75t_L g13593 ( 
.A(n_12731),
.Y(n_13593)
);

AOI22xp33_ASAP7_75t_L g13594 ( 
.A1(n_12749),
.A2(n_1034),
.B1(n_1031),
.B2(n_1033),
.Y(n_13594)
);

HB1xp67_ASAP7_75t_L g13595 ( 
.A(n_12761),
.Y(n_13595)
);

O2A1O1Ixp5_ASAP7_75t_L g13596 ( 
.A1(n_11937),
.A2(n_1034),
.B(n_1031),
.C(n_1033),
.Y(n_13596)
);

INVxp67_ASAP7_75t_SL g13597 ( 
.A(n_12761),
.Y(n_13597)
);

AOI21xp5_ASAP7_75t_L g13598 ( 
.A1(n_11937),
.A2(n_5649),
.B(n_5646),
.Y(n_13598)
);

OR2x6_ASAP7_75t_L g13599 ( 
.A(n_12432),
.B(n_5651),
.Y(n_13599)
);

INVx2_ASAP7_75t_L g13600 ( 
.A(n_12400),
.Y(n_13600)
);

AOI22xp33_ASAP7_75t_L g13601 ( 
.A1(n_12749),
.A2(n_1037),
.B1(n_1035),
.B2(n_1036),
.Y(n_13601)
);

AOI22x1_ASAP7_75t_L g13602 ( 
.A1(n_11937),
.A2(n_1038),
.B1(n_1035),
.B2(n_1036),
.Y(n_13602)
);

OAI22xp5_ASAP7_75t_L g13603 ( 
.A1(n_12155),
.A2(n_1040),
.B1(n_1038),
.B2(n_1039),
.Y(n_13603)
);

NOR2xp33_ASAP7_75t_L g13604 ( 
.A(n_12098),
.B(n_1039),
.Y(n_13604)
);

O2A1O1Ixp33_ASAP7_75t_L g13605 ( 
.A1(n_12749),
.A2(n_1042),
.B(n_1040),
.C(n_1041),
.Y(n_13605)
);

AOI22xp5_ASAP7_75t_L g13606 ( 
.A1(n_12749),
.A2(n_1044),
.B1(n_1041),
.B2(n_1043),
.Y(n_13606)
);

INVx3_ASAP7_75t_L g13607 ( 
.A(n_12097),
.Y(n_13607)
);

AOI22x1_ASAP7_75t_L g13608 ( 
.A1(n_11937),
.A2(n_1045),
.B1(n_1043),
.B2(n_1044),
.Y(n_13608)
);

BUFx2_ASAP7_75t_L g13609 ( 
.A(n_12638),
.Y(n_13609)
);

OAI21xp5_ASAP7_75t_L g13610 ( 
.A1(n_11937),
.A2(n_5653),
.B(n_5652),
.Y(n_13610)
);

OR2x6_ASAP7_75t_SL g13611 ( 
.A(n_12396),
.B(n_1045),
.Y(n_13611)
);

OAI21xp5_ASAP7_75t_L g13612 ( 
.A1(n_11937),
.A2(n_5655),
.B(n_5654),
.Y(n_13612)
);

AOI21xp5_ASAP7_75t_L g13613 ( 
.A1(n_11937),
.A2(n_5657),
.B(n_5656),
.Y(n_13613)
);

AOI21xp5_ASAP7_75t_L g13614 ( 
.A1(n_11937),
.A2(n_5660),
.B(n_5658),
.Y(n_13614)
);

AOI22xp5_ASAP7_75t_L g13615 ( 
.A1(n_12749),
.A2(n_1048),
.B1(n_1046),
.B2(n_1047),
.Y(n_13615)
);

O2A1O1Ixp33_ASAP7_75t_L g13616 ( 
.A1(n_12749),
.A2(n_1049),
.B(n_1047),
.C(n_1048),
.Y(n_13616)
);

INVxp67_ASAP7_75t_L g13617 ( 
.A(n_12761),
.Y(n_13617)
);

INVx2_ASAP7_75t_L g13618 ( 
.A(n_12400),
.Y(n_13618)
);

OAI21x1_ASAP7_75t_L g13619 ( 
.A1(n_12207),
.A2(n_5663),
.B(n_5662),
.Y(n_13619)
);

AOI21xp5_ASAP7_75t_L g13620 ( 
.A1(n_11937),
.A2(n_5665),
.B(n_5664),
.Y(n_13620)
);

OAI22xp5_ASAP7_75t_SL g13621 ( 
.A1(n_12696),
.A2(n_1051),
.B1(n_1049),
.B2(n_1050),
.Y(n_13621)
);

NAND2xp5_ASAP7_75t_L g13622 ( 
.A(n_12761),
.B(n_1051),
.Y(n_13622)
);

OR2x6_ASAP7_75t_SL g13623 ( 
.A(n_12396),
.B(n_1054),
.Y(n_13623)
);

NAND2xp5_ASAP7_75t_L g13624 ( 
.A(n_12761),
.B(n_1054),
.Y(n_13624)
);

INVx2_ASAP7_75t_SL g13625 ( 
.A(n_12167),
.Y(n_13625)
);

NAND2xp5_ASAP7_75t_L g13626 ( 
.A(n_12761),
.B(n_1055),
.Y(n_13626)
);

AOI21xp5_ASAP7_75t_L g13627 ( 
.A1(n_11937),
.A2(n_5667),
.B(n_5666),
.Y(n_13627)
);

AOI21xp5_ASAP7_75t_L g13628 ( 
.A1(n_11937),
.A2(n_5669),
.B(n_5668),
.Y(n_13628)
);

NAND2xp5_ASAP7_75t_L g13629 ( 
.A(n_12761),
.B(n_1055),
.Y(n_13629)
);

NAND2x1_ASAP7_75t_L g13630 ( 
.A(n_12189),
.B(n_5671),
.Y(n_13630)
);

BUFx6f_ASAP7_75t_L g13631 ( 
.A(n_11999),
.Y(n_13631)
);

NAND2xp5_ASAP7_75t_L g13632 ( 
.A(n_12761),
.B(n_1056),
.Y(n_13632)
);

O2A1O1Ixp5_ASAP7_75t_SL g13633 ( 
.A1(n_12440),
.A2(n_1059),
.B(n_1057),
.C(n_1058),
.Y(n_13633)
);

NAND2xp5_ASAP7_75t_L g13634 ( 
.A(n_12761),
.B(n_1057),
.Y(n_13634)
);

CKINVDCx11_ASAP7_75t_R g13635 ( 
.A(n_12072),
.Y(n_13635)
);

O2A1O1Ixp5_ASAP7_75t_L g13636 ( 
.A1(n_11937),
.A2(n_1060),
.B(n_1058),
.C(n_1059),
.Y(n_13636)
);

NAND2xp5_ASAP7_75t_L g13637 ( 
.A(n_12761),
.B(n_1061),
.Y(n_13637)
);

O2A1O1Ixp33_ASAP7_75t_L g13638 ( 
.A1(n_12749),
.A2(n_1063),
.B(n_1061),
.C(n_1062),
.Y(n_13638)
);

INVx3_ASAP7_75t_L g13639 ( 
.A(n_12097),
.Y(n_13639)
);

NAND2xp5_ASAP7_75t_L g13640 ( 
.A(n_12761),
.B(n_1062),
.Y(n_13640)
);

OAI22xp5_ASAP7_75t_L g13641 ( 
.A1(n_12155),
.A2(n_1065),
.B1(n_1063),
.B2(n_1064),
.Y(n_13641)
);

AOI21xp5_ASAP7_75t_L g13642 ( 
.A1(n_11937),
.A2(n_5675),
.B(n_5674),
.Y(n_13642)
);

O2A1O1Ixp33_ASAP7_75t_L g13643 ( 
.A1(n_12749),
.A2(n_1066),
.B(n_1064),
.C(n_1065),
.Y(n_13643)
);

INVx1_ASAP7_75t_L g13644 ( 
.A(n_12185),
.Y(n_13644)
);

OAI22xp5_ASAP7_75t_L g13645 ( 
.A1(n_12155),
.A2(n_1068),
.B1(n_1066),
.B2(n_1067),
.Y(n_13645)
);

AND2x2_ASAP7_75t_L g13646 ( 
.A(n_12302),
.B(n_1067),
.Y(n_13646)
);

AOI21xp5_ASAP7_75t_L g13647 ( 
.A1(n_11937),
.A2(n_5677),
.B(n_5676),
.Y(n_13647)
);

AOI21xp5_ASAP7_75t_L g13648 ( 
.A1(n_11937),
.A2(n_5683),
.B(n_5681),
.Y(n_13648)
);

AOI21xp5_ASAP7_75t_L g13649 ( 
.A1(n_11937),
.A2(n_5687),
.B(n_5685),
.Y(n_13649)
);

INVx1_ASAP7_75t_L g13650 ( 
.A(n_12185),
.Y(n_13650)
);

NOR2xp67_ASAP7_75t_L g13651 ( 
.A(n_12153),
.B(n_1068),
.Y(n_13651)
);

OAI22x1_ASAP7_75t_L g13652 ( 
.A1(n_12012),
.A2(n_1071),
.B1(n_1069),
.B2(n_1070),
.Y(n_13652)
);

A2O1A1Ixp33_ASAP7_75t_L g13653 ( 
.A1(n_11937),
.A2(n_1071),
.B(n_1069),
.C(n_1070),
.Y(n_13653)
);

NAND2xp5_ASAP7_75t_L g13654 ( 
.A(n_12761),
.B(n_1072),
.Y(n_13654)
);

INVx1_ASAP7_75t_SL g13655 ( 
.A(n_12548),
.Y(n_13655)
);

INVx1_ASAP7_75t_L g13656 ( 
.A(n_12185),
.Y(n_13656)
);

INVx2_ASAP7_75t_L g13657 ( 
.A(n_12400),
.Y(n_13657)
);

AOI21xp5_ASAP7_75t_L g13658 ( 
.A1(n_11937),
.A2(n_5689),
.B(n_5688),
.Y(n_13658)
);

NAND2xp5_ASAP7_75t_L g13659 ( 
.A(n_12761),
.B(n_1072),
.Y(n_13659)
);

NOR2xp33_ASAP7_75t_L g13660 ( 
.A(n_12098),
.B(n_1073),
.Y(n_13660)
);

O2A1O1Ixp33_ASAP7_75t_L g13661 ( 
.A1(n_12749),
.A2(n_1075),
.B(n_1073),
.C(n_1074),
.Y(n_13661)
);

AOI21xp5_ASAP7_75t_L g13662 ( 
.A1(n_11937),
.A2(n_5691),
.B(n_5690),
.Y(n_13662)
);

NAND2xp5_ASAP7_75t_SL g13663 ( 
.A(n_11937),
.B(n_5693),
.Y(n_13663)
);

NAND2xp5_ASAP7_75t_L g13664 ( 
.A(n_12761),
.B(n_1074),
.Y(n_13664)
);

BUFx2_ASAP7_75t_L g13665 ( 
.A(n_12638),
.Y(n_13665)
);

NAND2xp5_ASAP7_75t_SL g13666 ( 
.A(n_11937),
.B(n_5695),
.Y(n_13666)
);

NAND2xp5_ASAP7_75t_L g13667 ( 
.A(n_12761),
.B(n_1075),
.Y(n_13667)
);

NAND2xp5_ASAP7_75t_L g13668 ( 
.A(n_12761),
.B(n_1076),
.Y(n_13668)
);

AOI22xp33_ASAP7_75t_L g13669 ( 
.A1(n_12749),
.A2(n_1078),
.B1(n_1076),
.B2(n_1077),
.Y(n_13669)
);

NOR2xp33_ASAP7_75t_L g13670 ( 
.A(n_12098),
.B(n_1077),
.Y(n_13670)
);

NOR2xp33_ASAP7_75t_L g13671 ( 
.A(n_12098),
.B(n_1078),
.Y(n_13671)
);

AOI21xp5_ASAP7_75t_L g13672 ( 
.A1(n_11937),
.A2(n_5697),
.B(n_5696),
.Y(n_13672)
);

NAND2xp5_ASAP7_75t_L g13673 ( 
.A(n_12761),
.B(n_1079),
.Y(n_13673)
);

BUFx6f_ASAP7_75t_L g13674 ( 
.A(n_11999),
.Y(n_13674)
);

O2A1O1Ixp33_ASAP7_75t_L g13675 ( 
.A1(n_12749),
.A2(n_1081),
.B(n_1079),
.C(n_1080),
.Y(n_13675)
);

INVx1_ASAP7_75t_L g13676 ( 
.A(n_12185),
.Y(n_13676)
);

NAND2xp5_ASAP7_75t_L g13677 ( 
.A(n_12761),
.B(n_1080),
.Y(n_13677)
);

AND2x2_ASAP7_75t_L g13678 ( 
.A(n_12302),
.B(n_1081),
.Y(n_13678)
);

AOI21x1_ASAP7_75t_L g13679 ( 
.A1(n_11952),
.A2(n_1082),
.B(n_1083),
.Y(n_13679)
);

NAND2xp5_ASAP7_75t_L g13680 ( 
.A(n_12761),
.B(n_1082),
.Y(n_13680)
);

AOI21xp5_ASAP7_75t_L g13681 ( 
.A1(n_11937),
.A2(n_5699),
.B(n_5698),
.Y(n_13681)
);

BUFx6f_ASAP7_75t_L g13682 ( 
.A(n_11999),
.Y(n_13682)
);

HB1xp67_ASAP7_75t_L g13683 ( 
.A(n_12761),
.Y(n_13683)
);

AND2x2_ASAP7_75t_L g13684 ( 
.A(n_12302),
.B(n_1083),
.Y(n_13684)
);

AOI21xp5_ASAP7_75t_L g13685 ( 
.A1(n_11937),
.A2(n_5702),
.B(n_5701),
.Y(n_13685)
);

NOR2xp33_ASAP7_75t_L g13686 ( 
.A(n_12098),
.B(n_1084),
.Y(n_13686)
);

HB1xp67_ASAP7_75t_L g13687 ( 
.A(n_12761),
.Y(n_13687)
);

AOI22xp5_ASAP7_75t_L g13688 ( 
.A1(n_12749),
.A2(n_1087),
.B1(n_1085),
.B2(n_1086),
.Y(n_13688)
);

INVx1_ASAP7_75t_L g13689 ( 
.A(n_12185),
.Y(n_13689)
);

OAI22xp5_ASAP7_75t_L g13690 ( 
.A1(n_12155),
.A2(n_1087),
.B1(n_1085),
.B2(n_1086),
.Y(n_13690)
);

INVx2_ASAP7_75t_SL g13691 ( 
.A(n_12167),
.Y(n_13691)
);

NOR2xp33_ASAP7_75t_SL g13692 ( 
.A(n_12072),
.B(n_5703),
.Y(n_13692)
);

AOI22xp5_ASAP7_75t_L g13693 ( 
.A1(n_12749),
.A2(n_1090),
.B1(n_1088),
.B2(n_1089),
.Y(n_13693)
);

NAND2xp5_ASAP7_75t_L g13694 ( 
.A(n_12761),
.B(n_1088),
.Y(n_13694)
);

OAI21xp33_ASAP7_75t_SL g13695 ( 
.A1(n_12327),
.A2(n_1089),
.B(n_1090),
.Y(n_13695)
);

NAND2xp5_ASAP7_75t_L g13696 ( 
.A(n_12761),
.B(n_1091),
.Y(n_13696)
);

INVx1_ASAP7_75t_L g13697 ( 
.A(n_12185),
.Y(n_13697)
);

INVx2_ASAP7_75t_L g13698 ( 
.A(n_12400),
.Y(n_13698)
);

INVxp67_ASAP7_75t_L g13699 ( 
.A(n_12761),
.Y(n_13699)
);

BUFx6f_ASAP7_75t_L g13700 ( 
.A(n_11999),
.Y(n_13700)
);

AOI21xp5_ASAP7_75t_L g13701 ( 
.A1(n_11937),
.A2(n_5707),
.B(n_5706),
.Y(n_13701)
);

NOR2xp33_ASAP7_75t_SL g13702 ( 
.A(n_12072),
.B(n_5709),
.Y(n_13702)
);

AOI22xp33_ASAP7_75t_L g13703 ( 
.A1(n_12749),
.A2(n_1093),
.B1(n_1091),
.B2(n_1092),
.Y(n_13703)
);

A2O1A1Ixp33_ASAP7_75t_L g13704 ( 
.A1(n_11937),
.A2(n_1094),
.B(n_1092),
.C(n_1093),
.Y(n_13704)
);

AOI21xp5_ASAP7_75t_L g13705 ( 
.A1(n_11937),
.A2(n_5712),
.B(n_5711),
.Y(n_13705)
);

BUFx2_ASAP7_75t_L g13706 ( 
.A(n_12638),
.Y(n_13706)
);

NOR2xp33_ASAP7_75t_L g13707 ( 
.A(n_12098),
.B(n_1094),
.Y(n_13707)
);

AOI21xp5_ASAP7_75t_L g13708 ( 
.A1(n_11937),
.A2(n_5714),
.B(n_5713),
.Y(n_13708)
);

NOR2xp33_ASAP7_75t_L g13709 ( 
.A(n_12098),
.B(n_1095),
.Y(n_13709)
);

BUFx4f_ASAP7_75t_L g13710 ( 
.A(n_12303),
.Y(n_13710)
);

OAI22xp5_ASAP7_75t_L g13711 ( 
.A1(n_12155),
.A2(n_1098),
.B1(n_1096),
.B2(n_1097),
.Y(n_13711)
);

AOI221xp5_ASAP7_75t_L g13712 ( 
.A1(n_12561),
.A2(n_1099),
.B1(n_1097),
.B2(n_1098),
.C(n_1100),
.Y(n_13712)
);

AOI22x1_ASAP7_75t_L g13713 ( 
.A1(n_11937),
.A2(n_1101),
.B1(n_1099),
.B2(n_1100),
.Y(n_13713)
);

AOI21xp5_ASAP7_75t_L g13714 ( 
.A1(n_11937),
.A2(n_5716),
.B(n_5715),
.Y(n_13714)
);

INVx1_ASAP7_75t_SL g13715 ( 
.A(n_12548),
.Y(n_13715)
);

INVx3_ASAP7_75t_L g13716 ( 
.A(n_12097),
.Y(n_13716)
);

NAND2xp5_ASAP7_75t_L g13717 ( 
.A(n_12761),
.B(n_1101),
.Y(n_13717)
);

AOI21xp5_ASAP7_75t_L g13718 ( 
.A1(n_11937),
.A2(n_5719),
.B(n_5718),
.Y(n_13718)
);

BUFx2_ASAP7_75t_L g13719 ( 
.A(n_12638),
.Y(n_13719)
);

NAND2x1_ASAP7_75t_L g13720 ( 
.A(n_12189),
.B(n_5720),
.Y(n_13720)
);

BUFx6f_ASAP7_75t_L g13721 ( 
.A(n_11999),
.Y(n_13721)
);

INVx2_ASAP7_75t_SL g13722 ( 
.A(n_12167),
.Y(n_13722)
);

A2O1A1Ixp33_ASAP7_75t_L g13723 ( 
.A1(n_11937),
.A2(n_1104),
.B(n_1102),
.C(n_1103),
.Y(n_13723)
);

NOR2xp33_ASAP7_75t_L g13724 ( 
.A(n_12098),
.B(n_1102),
.Y(n_13724)
);

AOI22xp5_ASAP7_75t_L g13725 ( 
.A1(n_12749),
.A2(n_1105),
.B1(n_1103),
.B2(n_1104),
.Y(n_13725)
);

BUFx6f_ASAP7_75t_L g13726 ( 
.A(n_11999),
.Y(n_13726)
);

AOI21xp5_ASAP7_75t_L g13727 ( 
.A1(n_11937),
.A2(n_5722),
.B(n_5721),
.Y(n_13727)
);

AOI22xp5_ASAP7_75t_L g13728 ( 
.A1(n_12749),
.A2(n_1107),
.B1(n_1105),
.B2(n_1106),
.Y(n_13728)
);

NOR2xp67_ASAP7_75t_L g13729 ( 
.A(n_12153),
.B(n_1107),
.Y(n_13729)
);

INVx3_ASAP7_75t_L g13730 ( 
.A(n_12097),
.Y(n_13730)
);

INVx1_ASAP7_75t_L g13731 ( 
.A(n_12185),
.Y(n_13731)
);

INVx1_ASAP7_75t_L g13732 ( 
.A(n_12185),
.Y(n_13732)
);

INVx1_ASAP7_75t_L g13733 ( 
.A(n_12185),
.Y(n_13733)
);

AOI21xp5_ASAP7_75t_L g13734 ( 
.A1(n_11937),
.A2(n_5724),
.B(n_5723),
.Y(n_13734)
);

INVx1_ASAP7_75t_SL g13735 ( 
.A(n_12548),
.Y(n_13735)
);

NOR2xp33_ASAP7_75t_L g13736 ( 
.A(n_12098),
.B(n_1108),
.Y(n_13736)
);

NAND2xp5_ASAP7_75t_L g13737 ( 
.A(n_12761),
.B(n_1108),
.Y(n_13737)
);

O2A1O1Ixp33_ASAP7_75t_L g13738 ( 
.A1(n_12749),
.A2(n_1111),
.B(n_1109),
.C(n_1110),
.Y(n_13738)
);

NAND2xp5_ASAP7_75t_SL g13739 ( 
.A(n_11937),
.B(n_5725),
.Y(n_13739)
);

AOI21xp5_ASAP7_75t_L g13740 ( 
.A1(n_11937),
.A2(n_5727),
.B(n_5726),
.Y(n_13740)
);

NAND3xp33_ASAP7_75t_L g13741 ( 
.A(n_12749),
.B(n_1110),
.C(n_1111),
.Y(n_13741)
);

AND2x2_ASAP7_75t_L g13742 ( 
.A(n_12302),
.B(n_1112),
.Y(n_13742)
);

INVx1_ASAP7_75t_L g13743 ( 
.A(n_12185),
.Y(n_13743)
);

NAND2xp5_ASAP7_75t_L g13744 ( 
.A(n_12761),
.B(n_1112),
.Y(n_13744)
);

AOI21xp5_ASAP7_75t_L g13745 ( 
.A1(n_11937),
.A2(n_5729),
.B(n_5728),
.Y(n_13745)
);

AOI22xp5_ASAP7_75t_L g13746 ( 
.A1(n_12749),
.A2(n_1116),
.B1(n_1113),
.B2(n_1115),
.Y(n_13746)
);

INVx1_ASAP7_75t_SL g13747 ( 
.A(n_12548),
.Y(n_13747)
);

OAI21xp5_ASAP7_75t_L g13748 ( 
.A1(n_11937),
.A2(n_5731),
.B(n_5730),
.Y(n_13748)
);

OR2x2_ASAP7_75t_L g13749 ( 
.A(n_12761),
.B(n_1113),
.Y(n_13749)
);

BUFx12f_ASAP7_75t_L g13750 ( 
.A(n_12396),
.Y(n_13750)
);

OAI22xp5_ASAP7_75t_L g13751 ( 
.A1(n_12155),
.A2(n_1117),
.B1(n_1115),
.B2(n_1116),
.Y(n_13751)
);

BUFx8_ASAP7_75t_SL g13752 ( 
.A(n_12303),
.Y(n_13752)
);

AND2x2_ASAP7_75t_L g13753 ( 
.A(n_12302),
.B(n_1117),
.Y(n_13753)
);

INVx4_ASAP7_75t_L g13754 ( 
.A(n_12507),
.Y(n_13754)
);

NAND3xp33_ASAP7_75t_L g13755 ( 
.A(n_12749),
.B(n_1118),
.C(n_1119),
.Y(n_13755)
);

AOI21xp5_ASAP7_75t_L g13756 ( 
.A1(n_11937),
.A2(n_5735),
.B(n_5733),
.Y(n_13756)
);

AOI21xp5_ASAP7_75t_L g13757 ( 
.A1(n_11937),
.A2(n_5737),
.B(n_5736),
.Y(n_13757)
);

O2A1O1Ixp33_ASAP7_75t_L g13758 ( 
.A1(n_12749),
.A2(n_1120),
.B(n_1118),
.C(n_1119),
.Y(n_13758)
);

AND2x4_ASAP7_75t_L g13759 ( 
.A(n_12638),
.B(n_5738),
.Y(n_13759)
);

NAND2xp5_ASAP7_75t_L g13760 ( 
.A(n_12761),
.B(n_1120),
.Y(n_13760)
);

NAND2xp5_ASAP7_75t_L g13761 ( 
.A(n_12761),
.B(n_1121),
.Y(n_13761)
);

AOI21xp5_ASAP7_75t_L g13762 ( 
.A1(n_11937),
.A2(n_5741),
.B(n_5739),
.Y(n_13762)
);

INVx1_ASAP7_75t_L g13763 ( 
.A(n_12185),
.Y(n_13763)
);

AOI21xp5_ASAP7_75t_L g13764 ( 
.A1(n_11937),
.A2(n_5744),
.B(n_5742),
.Y(n_13764)
);

BUFx12f_ASAP7_75t_L g13765 ( 
.A(n_12396),
.Y(n_13765)
);

NAND2xp5_ASAP7_75t_L g13766 ( 
.A(n_12761),
.B(n_1121),
.Y(n_13766)
);

INVx2_ASAP7_75t_L g13767 ( 
.A(n_12400),
.Y(n_13767)
);

A2O1A1Ixp33_ASAP7_75t_L g13768 ( 
.A1(n_11937),
.A2(n_1124),
.B(n_1122),
.C(n_1123),
.Y(n_13768)
);

NAND2xp5_ASAP7_75t_SL g13769 ( 
.A(n_11937),
.B(n_5745),
.Y(n_13769)
);

AOI21xp5_ASAP7_75t_L g13770 ( 
.A1(n_11937),
.A2(n_5750),
.B(n_5748),
.Y(n_13770)
);

OAI22xp5_ASAP7_75t_L g13771 ( 
.A1(n_12155),
.A2(n_1124),
.B1(n_1122),
.B2(n_1123),
.Y(n_13771)
);

OAI22xp5_ASAP7_75t_L g13772 ( 
.A1(n_12155),
.A2(n_1127),
.B1(n_1125),
.B2(n_1126),
.Y(n_13772)
);

INVx1_ASAP7_75t_L g13773 ( 
.A(n_12185),
.Y(n_13773)
);

OR2x6_ASAP7_75t_L g13774 ( 
.A(n_12432),
.B(n_5752),
.Y(n_13774)
);

NAND2xp5_ASAP7_75t_SL g13775 ( 
.A(n_11937),
.B(n_5753),
.Y(n_13775)
);

AOI21xp5_ASAP7_75t_L g13776 ( 
.A1(n_11937),
.A2(n_5755),
.B(n_5754),
.Y(n_13776)
);

NAND2xp5_ASAP7_75t_SL g13777 ( 
.A(n_11937),
.B(n_5756),
.Y(n_13777)
);

AOI21xp5_ASAP7_75t_L g13778 ( 
.A1(n_11937),
.A2(n_5758),
.B(n_5757),
.Y(n_13778)
);

NAND2xp5_ASAP7_75t_L g13779 ( 
.A(n_12761),
.B(n_1125),
.Y(n_13779)
);

AOI21xp5_ASAP7_75t_L g13780 ( 
.A1(n_11937),
.A2(n_5761),
.B(n_5760),
.Y(n_13780)
);

AOI21xp5_ASAP7_75t_L g13781 ( 
.A1(n_11937),
.A2(n_5763),
.B(n_5762),
.Y(n_13781)
);

OAI22xp5_ASAP7_75t_L g13782 ( 
.A1(n_12155),
.A2(n_1129),
.B1(n_1126),
.B2(n_1127),
.Y(n_13782)
);

OAI22xp5_ASAP7_75t_L g13783 ( 
.A1(n_12155),
.A2(n_1131),
.B1(n_1129),
.B2(n_1130),
.Y(n_13783)
);

BUFx2_ASAP7_75t_L g13784 ( 
.A(n_12638),
.Y(n_13784)
);

HB1xp67_ASAP7_75t_L g13785 ( 
.A(n_12761),
.Y(n_13785)
);

INVx2_ASAP7_75t_L g13786 ( 
.A(n_12400),
.Y(n_13786)
);

NAND2xp5_ASAP7_75t_L g13787 ( 
.A(n_12761),
.B(n_1130),
.Y(n_13787)
);

NAND2xp5_ASAP7_75t_L g13788 ( 
.A(n_12761),
.B(n_1132),
.Y(n_13788)
);

BUFx2_ASAP7_75t_L g13789 ( 
.A(n_12638),
.Y(n_13789)
);

NOR2xp67_ASAP7_75t_L g13790 ( 
.A(n_12153),
.B(n_1132),
.Y(n_13790)
);

AND2x4_ASAP7_75t_L g13791 ( 
.A(n_12638),
.B(n_5764),
.Y(n_13791)
);

AND2x4_ASAP7_75t_L g13792 ( 
.A(n_12638),
.B(n_5765),
.Y(n_13792)
);

AOI21xp5_ASAP7_75t_L g13793 ( 
.A1(n_11937),
.A2(n_5767),
.B(n_5766),
.Y(n_13793)
);

NAND2xp5_ASAP7_75t_SL g13794 ( 
.A(n_11937),
.B(n_5768),
.Y(n_13794)
);

INVx2_ASAP7_75t_L g13795 ( 
.A(n_12400),
.Y(n_13795)
);

A2O1A1Ixp33_ASAP7_75t_L g13796 ( 
.A1(n_11937),
.A2(n_1135),
.B(n_1133),
.C(n_1134),
.Y(n_13796)
);

OAI22xp5_ASAP7_75t_L g13797 ( 
.A1(n_12155),
.A2(n_1136),
.B1(n_1133),
.B2(n_1135),
.Y(n_13797)
);

OAI22x1_ASAP7_75t_L g13798 ( 
.A1(n_12012),
.A2(n_1139),
.B1(n_1137),
.B2(n_1138),
.Y(n_13798)
);

OAI21xp5_ASAP7_75t_L g13799 ( 
.A1(n_11937),
.A2(n_5770),
.B(n_5769),
.Y(n_13799)
);

INVx2_ASAP7_75t_L g13800 ( 
.A(n_12400),
.Y(n_13800)
);

NOR2xp33_ASAP7_75t_L g13801 ( 
.A(n_12098),
.B(n_1137),
.Y(n_13801)
);

AOI21xp5_ASAP7_75t_L g13802 ( 
.A1(n_11937),
.A2(n_5772),
.B(n_5771),
.Y(n_13802)
);

NAND2xp5_ASAP7_75t_SL g13803 ( 
.A(n_11937),
.B(n_5773),
.Y(n_13803)
);

INVx2_ASAP7_75t_L g13804 ( 
.A(n_12400),
.Y(n_13804)
);

INVx2_ASAP7_75t_L g13805 ( 
.A(n_12400),
.Y(n_13805)
);

BUFx2_ASAP7_75t_L g13806 ( 
.A(n_12638),
.Y(n_13806)
);

AOI21xp5_ASAP7_75t_L g13807 ( 
.A1(n_11937),
.A2(n_5776),
.B(n_5774),
.Y(n_13807)
);

AO32x2_ASAP7_75t_L g13808 ( 
.A1(n_12491),
.A2(n_1140),
.A3(n_1138),
.B1(n_1139),
.B2(n_1141),
.Y(n_13808)
);

BUFx6f_ASAP7_75t_L g13809 ( 
.A(n_11999),
.Y(n_13809)
);

AOI21xp5_ASAP7_75t_L g13810 ( 
.A1(n_11937),
.A2(n_5778),
.B(n_5777),
.Y(n_13810)
);

INVx1_ASAP7_75t_L g13811 ( 
.A(n_12185),
.Y(n_13811)
);

AND2x4_ASAP7_75t_L g13812 ( 
.A(n_12638),
.B(n_5781),
.Y(n_13812)
);

NAND2xp5_ASAP7_75t_L g13813 ( 
.A(n_12761),
.B(n_1140),
.Y(n_13813)
);

O2A1O1Ixp33_ASAP7_75t_L g13814 ( 
.A1(n_12749),
.A2(n_1143),
.B(n_1141),
.C(n_1142),
.Y(n_13814)
);

INVx2_ASAP7_75t_SL g13815 ( 
.A(n_12167),
.Y(n_13815)
);

AOI21xp5_ASAP7_75t_L g13816 ( 
.A1(n_11937),
.A2(n_5783),
.B(n_5782),
.Y(n_13816)
);

AND2x2_ASAP7_75t_L g13817 ( 
.A(n_12302),
.B(n_1142),
.Y(n_13817)
);

AND2x2_ASAP7_75t_L g13818 ( 
.A(n_12302),
.B(n_1143),
.Y(n_13818)
);

NAND2xp5_ASAP7_75t_L g13819 ( 
.A(n_12761),
.B(n_1144),
.Y(n_13819)
);

AOI21x1_ASAP7_75t_L g13820 ( 
.A1(n_11952),
.A2(n_1144),
.B(n_1145),
.Y(n_13820)
);

INVx2_ASAP7_75t_L g13821 ( 
.A(n_12400),
.Y(n_13821)
);

A2O1A1Ixp33_ASAP7_75t_L g13822 ( 
.A1(n_11937),
.A2(n_1147),
.B(n_1145),
.C(n_1146),
.Y(n_13822)
);

NOR2xp33_ASAP7_75t_L g13823 ( 
.A(n_12098),
.B(n_1146),
.Y(n_13823)
);

NAND2xp5_ASAP7_75t_SL g13824 ( 
.A(n_11937),
.B(n_5784),
.Y(n_13824)
);

AOI21xp5_ASAP7_75t_L g13825 ( 
.A1(n_11937),
.A2(n_5787),
.B(n_5785),
.Y(n_13825)
);

NAND2xp5_ASAP7_75t_SL g13826 ( 
.A(n_11937),
.B(n_5791),
.Y(n_13826)
);

CKINVDCx11_ASAP7_75t_R g13827 ( 
.A(n_12072),
.Y(n_13827)
);

NAND2xp5_ASAP7_75t_SL g13828 ( 
.A(n_11937),
.B(n_5792),
.Y(n_13828)
);

INVx2_ASAP7_75t_L g13829 ( 
.A(n_12400),
.Y(n_13829)
);

AND2x2_ASAP7_75t_SL g13830 ( 
.A(n_12326),
.B(n_1147),
.Y(n_13830)
);

AOI21xp5_ASAP7_75t_L g13831 ( 
.A1(n_11937),
.A2(n_5794),
.B(n_5793),
.Y(n_13831)
);

AOI22xp5_ASAP7_75t_L g13832 ( 
.A1(n_12749),
.A2(n_1150),
.B1(n_1148),
.B2(n_1149),
.Y(n_13832)
);

O2A1O1Ixp33_ASAP7_75t_L g13833 ( 
.A1(n_12749),
.A2(n_1150),
.B(n_1148),
.C(n_1149),
.Y(n_13833)
);

NOR2xp33_ASAP7_75t_SL g13834 ( 
.A(n_12072),
.B(n_5795),
.Y(n_13834)
);

NAND2xp33_ASAP7_75t_L g13835 ( 
.A(n_12561),
.B(n_1151),
.Y(n_13835)
);

INVx3_ASAP7_75t_L g13836 ( 
.A(n_12097),
.Y(n_13836)
);

AOI21xp5_ASAP7_75t_L g13837 ( 
.A1(n_11937),
.A2(n_5797),
.B(n_5796),
.Y(n_13837)
);

AOI22xp33_ASAP7_75t_L g13838 ( 
.A1(n_12749),
.A2(n_1153),
.B1(n_1151),
.B2(n_1152),
.Y(n_13838)
);

AOI21xp5_ASAP7_75t_L g13839 ( 
.A1(n_11937),
.A2(n_5799),
.B(n_5798),
.Y(n_13839)
);

INVx2_ASAP7_75t_L g13840 ( 
.A(n_12400),
.Y(n_13840)
);

NAND2xp5_ASAP7_75t_L g13841 ( 
.A(n_12761),
.B(n_1152),
.Y(n_13841)
);

INVx1_ASAP7_75t_L g13842 ( 
.A(n_12185),
.Y(n_13842)
);

AOI21xp5_ASAP7_75t_L g13843 ( 
.A1(n_11937),
.A2(n_5801),
.B(n_5800),
.Y(n_13843)
);

NAND2xp5_ASAP7_75t_L g13844 ( 
.A(n_12761),
.B(n_1153),
.Y(n_13844)
);

OR2x6_ASAP7_75t_SL g13845 ( 
.A(n_12396),
.B(n_1154),
.Y(n_13845)
);

NAND2xp5_ASAP7_75t_SL g13846 ( 
.A(n_11937),
.B(n_5802),
.Y(n_13846)
);

OAI22xp5_ASAP7_75t_L g13847 ( 
.A1(n_12155),
.A2(n_1156),
.B1(n_1154),
.B2(n_1155),
.Y(n_13847)
);

O2A1O1Ixp5_ASAP7_75t_L g13848 ( 
.A1(n_11937),
.A2(n_1157),
.B(n_1155),
.C(n_1156),
.Y(n_13848)
);

NAND2x1p5_ASAP7_75t_L g13849 ( 
.A(n_12304),
.B(n_5803),
.Y(n_13849)
);

BUFx2_ASAP7_75t_L g13850 ( 
.A(n_12638),
.Y(n_13850)
);

INVx1_ASAP7_75t_L g13851 ( 
.A(n_12185),
.Y(n_13851)
);

A2O1A1Ixp33_ASAP7_75t_L g13852 ( 
.A1(n_11937),
.A2(n_1159),
.B(n_1157),
.C(n_1158),
.Y(n_13852)
);

NAND2xp5_ASAP7_75t_L g13853 ( 
.A(n_12761),
.B(n_1158),
.Y(n_13853)
);

AOI21xp5_ASAP7_75t_L g13854 ( 
.A1(n_11937),
.A2(n_5805),
.B(n_5804),
.Y(n_13854)
);

BUFx3_ASAP7_75t_L g13855 ( 
.A(n_11999),
.Y(n_13855)
);

AOI21xp5_ASAP7_75t_L g13856 ( 
.A1(n_11937),
.A2(n_5807),
.B(n_5806),
.Y(n_13856)
);

NAND2xp5_ASAP7_75t_L g13857 ( 
.A(n_12761),
.B(n_1159),
.Y(n_13857)
);

NAND2xp33_ASAP7_75t_L g13858 ( 
.A(n_12561),
.B(n_1160),
.Y(n_13858)
);

NAND2xp5_ASAP7_75t_L g13859 ( 
.A(n_12761),
.B(n_1160),
.Y(n_13859)
);

NAND2xp5_ASAP7_75t_SL g13860 ( 
.A(n_11937),
.B(n_5808),
.Y(n_13860)
);

INVx2_ASAP7_75t_L g13861 ( 
.A(n_12400),
.Y(n_13861)
);

AOI21x1_ASAP7_75t_L g13862 ( 
.A1(n_11952),
.A2(n_1161),
.B(n_1162),
.Y(n_13862)
);

A2O1A1Ixp33_ASAP7_75t_L g13863 ( 
.A1(n_11937),
.A2(n_1163),
.B(n_1161),
.C(n_1162),
.Y(n_13863)
);

NAND2xp5_ASAP7_75t_L g13864 ( 
.A(n_12761),
.B(n_1163),
.Y(n_13864)
);

INVx2_ASAP7_75t_L g13865 ( 
.A(n_12400),
.Y(n_13865)
);

INVx2_ASAP7_75t_L g13866 ( 
.A(n_12400),
.Y(n_13866)
);

INVx1_ASAP7_75t_L g13867 ( 
.A(n_12185),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_12185),
.Y(n_13868)
);

AOI21xp5_ASAP7_75t_L g13869 ( 
.A1(n_11937),
.A2(n_5810),
.B(n_5809),
.Y(n_13869)
);

OAI21xp5_ASAP7_75t_L g13870 ( 
.A1(n_11937),
.A2(n_5813),
.B(n_5811),
.Y(n_13870)
);

AOI21xp5_ASAP7_75t_L g13871 ( 
.A1(n_11937),
.A2(n_5815),
.B(n_5814),
.Y(n_13871)
);

BUFx2_ASAP7_75t_L g13872 ( 
.A(n_12638),
.Y(n_13872)
);

AOI22xp5_ASAP7_75t_L g13873 ( 
.A1(n_12749),
.A2(n_1166),
.B1(n_1164),
.B2(n_1165),
.Y(n_13873)
);

NAND2xp5_ASAP7_75t_L g13874 ( 
.A(n_12761),
.B(n_1164),
.Y(n_13874)
);

AOI22xp33_ASAP7_75t_L g13875 ( 
.A1(n_12749),
.A2(n_1167),
.B1(n_1165),
.B2(n_1166),
.Y(n_13875)
);

NAND2x1_ASAP7_75t_L g13876 ( 
.A(n_12189),
.B(n_5816),
.Y(n_13876)
);

AO21x2_ASAP7_75t_L g13877 ( 
.A1(n_11952),
.A2(n_1167),
.B(n_1168),
.Y(n_13877)
);

NAND2xp5_ASAP7_75t_L g13878 ( 
.A(n_12761),
.B(n_1168),
.Y(n_13878)
);

NOR2xp33_ASAP7_75t_L g13879 ( 
.A(n_12098),
.B(n_1169),
.Y(n_13879)
);

NAND2xp5_ASAP7_75t_L g13880 ( 
.A(n_12761),
.B(n_1169),
.Y(n_13880)
);

NAND2x1p5_ASAP7_75t_L g13881 ( 
.A(n_12304),
.B(n_5817),
.Y(n_13881)
);

NAND2xp5_ASAP7_75t_SL g13882 ( 
.A(n_11937),
.B(n_5818),
.Y(n_13882)
);

AOI22xp5_ASAP7_75t_L g13883 ( 
.A1(n_12749),
.A2(n_1172),
.B1(n_1170),
.B2(n_1171),
.Y(n_13883)
);

INVx2_ASAP7_75t_L g13884 ( 
.A(n_12400),
.Y(n_13884)
);

AOI22xp5_ASAP7_75t_L g13885 ( 
.A1(n_12749),
.A2(n_1173),
.B1(n_1171),
.B2(n_1172),
.Y(n_13885)
);

NAND2xp5_ASAP7_75t_L g13886 ( 
.A(n_12761),
.B(n_1173),
.Y(n_13886)
);

BUFx4f_ASAP7_75t_L g13887 ( 
.A(n_12303),
.Y(n_13887)
);

OAI22xp5_ASAP7_75t_L g13888 ( 
.A1(n_12155),
.A2(n_1176),
.B1(n_1174),
.B2(n_1175),
.Y(n_13888)
);

BUFx8_ASAP7_75t_L g13889 ( 
.A(n_12303),
.Y(n_13889)
);

CKINVDCx20_ASAP7_75t_R g13890 ( 
.A(n_12632),
.Y(n_13890)
);

NAND2xp5_ASAP7_75t_SL g13891 ( 
.A(n_11937),
.B(n_5820),
.Y(n_13891)
);

AOI22xp33_ASAP7_75t_L g13892 ( 
.A1(n_12749),
.A2(n_1177),
.B1(n_1174),
.B2(n_1175),
.Y(n_13892)
);

CKINVDCx14_ASAP7_75t_R g13893 ( 
.A(n_12396),
.Y(n_13893)
);

AOI21xp5_ASAP7_75t_L g13894 ( 
.A1(n_11937),
.A2(n_5822),
.B(n_5821),
.Y(n_13894)
);

CKINVDCx16_ASAP7_75t_R g13895 ( 
.A(n_12303),
.Y(n_13895)
);

A2O1A1Ixp33_ASAP7_75t_L g13896 ( 
.A1(n_11937),
.A2(n_1180),
.B(n_1177),
.C(n_1179),
.Y(n_13896)
);

OAI22xp5_ASAP7_75t_L g13897 ( 
.A1(n_12155),
.A2(n_1181),
.B1(n_1179),
.B2(n_1180),
.Y(n_13897)
);

NAND2xp5_ASAP7_75t_L g13898 ( 
.A(n_12761),
.B(n_1181),
.Y(n_13898)
);

AOI21xp5_ASAP7_75t_L g13899 ( 
.A1(n_11937),
.A2(n_5824),
.B(n_5823),
.Y(n_13899)
);

NAND2xp5_ASAP7_75t_L g13900 ( 
.A(n_12761),
.B(n_1182),
.Y(n_13900)
);

NOR2xp33_ASAP7_75t_L g13901 ( 
.A(n_12098),
.B(n_1182),
.Y(n_13901)
);

CKINVDCx5p33_ASAP7_75t_R g13902 ( 
.A(n_13635),
.Y(n_13902)
);

AOI22xp33_ASAP7_75t_L g13903 ( 
.A1(n_13115),
.A2(n_1185),
.B1(n_1183),
.B2(n_1184),
.Y(n_13903)
);

INVx2_ASAP7_75t_L g13904 ( 
.A(n_12863),
.Y(n_13904)
);

NAND2x1p5_ASAP7_75t_L g13905 ( 
.A(n_12793),
.B(n_5825),
.Y(n_13905)
);

INVx1_ASAP7_75t_L g13906 ( 
.A(n_12898),
.Y(n_13906)
);

NAND2xp5_ASAP7_75t_L g13907 ( 
.A(n_13091),
.B(n_1183),
.Y(n_13907)
);

AND2x2_ASAP7_75t_L g13908 ( 
.A(n_13609),
.B(n_1186),
.Y(n_13908)
);

AND2x2_ASAP7_75t_L g13909 ( 
.A(n_13665),
.B(n_1186),
.Y(n_13909)
);

AND2x2_ASAP7_75t_L g13910 ( 
.A(n_13706),
.B(n_1187),
.Y(n_13910)
);

INVx2_ASAP7_75t_L g13911 ( 
.A(n_12881),
.Y(n_13911)
);

AOI21xp33_ASAP7_75t_L g13912 ( 
.A1(n_12827),
.A2(n_13858),
.B(n_13835),
.Y(n_13912)
);

CKINVDCx5p33_ASAP7_75t_R g13913 ( 
.A(n_13827),
.Y(n_13913)
);

INVx2_ASAP7_75t_L g13914 ( 
.A(n_12892),
.Y(n_13914)
);

A2O1A1Ixp33_ASAP7_75t_SL g13915 ( 
.A1(n_13127),
.A2(n_1189),
.B(n_1187),
.C(n_1188),
.Y(n_13915)
);

AOI22xp5_ASAP7_75t_SL g13916 ( 
.A1(n_13318),
.A2(n_1192),
.B1(n_1190),
.B2(n_1191),
.Y(n_13916)
);

CKINVDCx16_ASAP7_75t_R g13917 ( 
.A(n_13895),
.Y(n_13917)
);

NAND2xp5_ASAP7_75t_L g13918 ( 
.A(n_13597),
.B(n_1191),
.Y(n_13918)
);

NAND3xp33_ASAP7_75t_SL g13919 ( 
.A(n_12890),
.B(n_1193),
.C(n_1194),
.Y(n_13919)
);

NAND2xp5_ASAP7_75t_L g13920 ( 
.A(n_13595),
.B(n_1193),
.Y(n_13920)
);

HB1xp67_ASAP7_75t_L g13921 ( 
.A(n_13683),
.Y(n_13921)
);

NAND2xp5_ASAP7_75t_L g13922 ( 
.A(n_13687),
.B(n_1195),
.Y(n_13922)
);

INVx2_ASAP7_75t_L g13923 ( 
.A(n_12893),
.Y(n_13923)
);

NAND2xp5_ASAP7_75t_L g13924 ( 
.A(n_13785),
.B(n_1195),
.Y(n_13924)
);

INVx4_ASAP7_75t_L g13925 ( 
.A(n_13264),
.Y(n_13925)
);

NAND2xp5_ASAP7_75t_L g13926 ( 
.A(n_13617),
.B(n_1196),
.Y(n_13926)
);

INVx1_ASAP7_75t_L g13927 ( 
.A(n_12909),
.Y(n_13927)
);

INVxp67_ASAP7_75t_L g13928 ( 
.A(n_12852),
.Y(n_13928)
);

NAND2xp5_ASAP7_75t_SL g13929 ( 
.A(n_12793),
.B(n_5826),
.Y(n_13929)
);

NAND2xp5_ASAP7_75t_L g13930 ( 
.A(n_13699),
.B(n_1196),
.Y(n_13930)
);

NAND2xp5_ASAP7_75t_L g13931 ( 
.A(n_13052),
.B(n_1197),
.Y(n_13931)
);

AND2x2_ASAP7_75t_L g13932 ( 
.A(n_13719),
.B(n_1197),
.Y(n_13932)
);

INVx2_ASAP7_75t_L g13933 ( 
.A(n_12920),
.Y(n_13933)
);

HB1xp67_ASAP7_75t_L g13934 ( 
.A(n_12807),
.Y(n_13934)
);

INVxp33_ASAP7_75t_SL g13935 ( 
.A(n_13077),
.Y(n_13935)
);

NAND2xp5_ASAP7_75t_L g13936 ( 
.A(n_13066),
.B(n_1198),
.Y(n_13936)
);

BUFx2_ASAP7_75t_L g13937 ( 
.A(n_13784),
.Y(n_13937)
);

INVx1_ASAP7_75t_L g13938 ( 
.A(n_12910),
.Y(n_13938)
);

AND2x2_ASAP7_75t_L g13939 ( 
.A(n_13789),
.B(n_1198),
.Y(n_13939)
);

OAI22xp5_ASAP7_75t_SL g13940 ( 
.A1(n_13386),
.A2(n_1201),
.B1(n_1199),
.B2(n_1200),
.Y(n_13940)
);

AND2x2_ASAP7_75t_L g13941 ( 
.A(n_13806),
.B(n_1199),
.Y(n_13941)
);

INVx2_ASAP7_75t_L g13942 ( 
.A(n_12935),
.Y(n_13942)
);

NAND2xp5_ASAP7_75t_L g13943 ( 
.A(n_13078),
.B(n_1200),
.Y(n_13943)
);

CKINVDCx5p33_ASAP7_75t_R g13944 ( 
.A(n_13890),
.Y(n_13944)
);

AOI22xp5_ASAP7_75t_L g13945 ( 
.A1(n_13191),
.A2(n_1203),
.B1(n_1201),
.B2(n_1202),
.Y(n_13945)
);

BUFx2_ASAP7_75t_L g13946 ( 
.A(n_13850),
.Y(n_13946)
);

AND3x1_ASAP7_75t_SL g13947 ( 
.A(n_13712),
.B(n_1202),
.C(n_1204),
.Y(n_13947)
);

NAND2xp5_ASAP7_75t_L g13948 ( 
.A(n_13089),
.B(n_1204),
.Y(n_13948)
);

INVx1_ASAP7_75t_L g13949 ( 
.A(n_12914),
.Y(n_13949)
);

INVx1_ASAP7_75t_L g13950 ( 
.A(n_12928),
.Y(n_13950)
);

INVx5_ASAP7_75t_L g13951 ( 
.A(n_13599),
.Y(n_13951)
);

OAI22xp5_ASAP7_75t_L g13952 ( 
.A1(n_13606),
.A2(n_1207),
.B1(n_1205),
.B2(n_1206),
.Y(n_13952)
);

INVx1_ASAP7_75t_L g13953 ( 
.A(n_12934),
.Y(n_13953)
);

CKINVDCx5p33_ASAP7_75t_R g13954 ( 
.A(n_12811),
.Y(n_13954)
);

AND2x2_ASAP7_75t_L g13955 ( 
.A(n_13872),
.B(n_1205),
.Y(n_13955)
);

INVx4_ASAP7_75t_L g13956 ( 
.A(n_13376),
.Y(n_13956)
);

BUFx2_ASAP7_75t_L g13957 ( 
.A(n_12895),
.Y(n_13957)
);

INVx1_ASAP7_75t_L g13958 ( 
.A(n_12973),
.Y(n_13958)
);

BUFx3_ASAP7_75t_L g13959 ( 
.A(n_13855),
.Y(n_13959)
);

BUFx6f_ASAP7_75t_L g13960 ( 
.A(n_12797),
.Y(n_13960)
);

BUFx2_ASAP7_75t_L g13961 ( 
.A(n_13152),
.Y(n_13961)
);

CKINVDCx16_ASAP7_75t_R g13962 ( 
.A(n_12916),
.Y(n_13962)
);

AOI22xp33_ASAP7_75t_L g13963 ( 
.A1(n_13353),
.A2(n_1208),
.B1(n_1206),
.B2(n_1207),
.Y(n_13963)
);

INVx2_ASAP7_75t_L g13964 ( 
.A(n_12982),
.Y(n_13964)
);

INVx1_ASAP7_75t_L g13965 ( 
.A(n_12983),
.Y(n_13965)
);

AND2x2_ASAP7_75t_L g13966 ( 
.A(n_12924),
.B(n_1208),
.Y(n_13966)
);

INVx1_ASAP7_75t_L g13967 ( 
.A(n_12987),
.Y(n_13967)
);

CKINVDCx5p33_ASAP7_75t_R g13968 ( 
.A(n_13752),
.Y(n_13968)
);

OAI22xp5_ASAP7_75t_SL g13969 ( 
.A1(n_13150),
.A2(n_1211),
.B1(n_1209),
.B2(n_1210),
.Y(n_13969)
);

CKINVDCx5p33_ASAP7_75t_R g13970 ( 
.A(n_12867),
.Y(n_13970)
);

BUFx6f_ASAP7_75t_L g13971 ( 
.A(n_12797),
.Y(n_13971)
);

INVx3_ASAP7_75t_L g13972 ( 
.A(n_12889),
.Y(n_13972)
);

NAND2xp5_ASAP7_75t_L g13973 ( 
.A(n_13303),
.B(n_1209),
.Y(n_13973)
);

INVx3_ASAP7_75t_L g13974 ( 
.A(n_12889),
.Y(n_13974)
);

NAND2xp5_ASAP7_75t_L g13975 ( 
.A(n_13456),
.B(n_1210),
.Y(n_13975)
);

INVx2_ASAP7_75t_L g13976 ( 
.A(n_12985),
.Y(n_13976)
);

INVx1_ASAP7_75t_L g13977 ( 
.A(n_12989),
.Y(n_13977)
);

INVx2_ASAP7_75t_L g13978 ( 
.A(n_12834),
.Y(n_13978)
);

NAND2xp5_ASAP7_75t_L g13979 ( 
.A(n_13220),
.B(n_1211),
.Y(n_13979)
);

AOI22xp5_ASAP7_75t_L g13980 ( 
.A1(n_12915),
.A2(n_1214),
.B1(n_1212),
.B2(n_1213),
.Y(n_13980)
);

AND2x2_ASAP7_75t_L g13981 ( 
.A(n_13045),
.B(n_1213),
.Y(n_13981)
);

AOI22xp33_ASAP7_75t_L g13982 ( 
.A1(n_13256),
.A2(n_1216),
.B1(n_1214),
.B2(n_1215),
.Y(n_13982)
);

BUFx6f_ASAP7_75t_L g13983 ( 
.A(n_13631),
.Y(n_13983)
);

NOR2xp33_ASAP7_75t_SL g13984 ( 
.A(n_13126),
.B(n_5829),
.Y(n_13984)
);

OR2x2_ASAP7_75t_L g13985 ( 
.A(n_12808),
.B(n_1217),
.Y(n_13985)
);

HB1xp67_ASAP7_75t_L g13986 ( 
.A(n_12854),
.Y(n_13986)
);

HB1xp67_ASAP7_75t_L g13987 ( 
.A(n_13644),
.Y(n_13987)
);

NAND2xp5_ASAP7_75t_L g13988 ( 
.A(n_13158),
.B(n_1217),
.Y(n_13988)
);

AND2x2_ASAP7_75t_L g13989 ( 
.A(n_13005),
.B(n_1218),
.Y(n_13989)
);

NOR2xp33_ASAP7_75t_L g13990 ( 
.A(n_13439),
.B(n_1218),
.Y(n_13990)
);

NAND2xp5_ASAP7_75t_L g13991 ( 
.A(n_13160),
.B(n_1219),
.Y(n_13991)
);

BUFx6f_ASAP7_75t_L g13992 ( 
.A(n_13631),
.Y(n_13992)
);

INVx2_ASAP7_75t_L g13993 ( 
.A(n_13600),
.Y(n_13993)
);

INVx2_ASAP7_75t_L g13994 ( 
.A(n_13618),
.Y(n_13994)
);

NAND2xp5_ASAP7_75t_SL g13995 ( 
.A(n_12793),
.B(n_5830),
.Y(n_13995)
);

NOR2xp67_ASAP7_75t_L g13996 ( 
.A(n_13539),
.B(n_1219),
.Y(n_13996)
);

NAND2xp5_ASAP7_75t_L g13997 ( 
.A(n_13272),
.B(n_1220),
.Y(n_13997)
);

NAND2xp5_ASAP7_75t_SL g13998 ( 
.A(n_13270),
.B(n_5832),
.Y(n_13998)
);

AOI22xp5_ASAP7_75t_L g13999 ( 
.A1(n_13374),
.A2(n_1223),
.B1(n_1220),
.B2(n_1222),
.Y(n_13999)
);

NOR2xp33_ASAP7_75t_L g14000 ( 
.A(n_12826),
.B(n_1222),
.Y(n_14000)
);

AOI22xp5_ASAP7_75t_L g14001 ( 
.A1(n_13141),
.A2(n_1225),
.B1(n_1223),
.B2(n_1224),
.Y(n_14001)
);

NAND2xp5_ASAP7_75t_L g14002 ( 
.A(n_13295),
.B(n_13307),
.Y(n_14002)
);

INVx1_ASAP7_75t_L g14003 ( 
.A(n_13008),
.Y(n_14003)
);

INVx2_ASAP7_75t_L g14004 ( 
.A(n_13657),
.Y(n_14004)
);

CKINVDCx11_ASAP7_75t_R g14005 ( 
.A(n_12823),
.Y(n_14005)
);

NAND2xp5_ASAP7_75t_L g14006 ( 
.A(n_13650),
.B(n_1224),
.Y(n_14006)
);

NAND2xp5_ASAP7_75t_L g14007 ( 
.A(n_13656),
.B(n_1225),
.Y(n_14007)
);

OAI21xp5_ASAP7_75t_L g14008 ( 
.A1(n_12795),
.A2(n_1226),
.B(n_1227),
.Y(n_14008)
);

NAND2xp5_ASAP7_75t_SL g14009 ( 
.A(n_13270),
.B(n_5833),
.Y(n_14009)
);

NOR2xp33_ASAP7_75t_R g14010 ( 
.A(n_13893),
.B(n_1226),
.Y(n_14010)
);

INVx3_ASAP7_75t_L g14011 ( 
.A(n_12926),
.Y(n_14011)
);

CKINVDCx5p33_ASAP7_75t_R g14012 ( 
.A(n_13365),
.Y(n_14012)
);

CKINVDCx5p33_ASAP7_75t_R g14013 ( 
.A(n_12812),
.Y(n_14013)
);

NAND2xp5_ASAP7_75t_L g14014 ( 
.A(n_13676),
.B(n_13689),
.Y(n_14014)
);

AND2x2_ASAP7_75t_L g14015 ( 
.A(n_13041),
.B(n_1227),
.Y(n_14015)
);

AND3x1_ASAP7_75t_SL g14016 ( 
.A(n_13151),
.B(n_1228),
.C(n_1229),
.Y(n_14016)
);

CKINVDCx5p33_ASAP7_75t_R g14017 ( 
.A(n_13750),
.Y(n_14017)
);

BUFx10_ASAP7_75t_L g14018 ( 
.A(n_13674),
.Y(n_14018)
);

CKINVDCx5p33_ASAP7_75t_R g14019 ( 
.A(n_13765),
.Y(n_14019)
);

INVx2_ASAP7_75t_L g14020 ( 
.A(n_13698),
.Y(n_14020)
);

OAI22xp5_ASAP7_75t_SL g14021 ( 
.A1(n_13162),
.A2(n_13104),
.B1(n_13090),
.B2(n_13621),
.Y(n_14021)
);

INVx2_ASAP7_75t_SL g14022 ( 
.A(n_13140),
.Y(n_14022)
);

INVx1_ASAP7_75t_L g14023 ( 
.A(n_13697),
.Y(n_14023)
);

AOI21xp5_ASAP7_75t_L g14024 ( 
.A1(n_12970),
.A2(n_1228),
.B(n_1229),
.Y(n_14024)
);

NAND2xp5_ASAP7_75t_L g14025 ( 
.A(n_13731),
.B(n_1230),
.Y(n_14025)
);

BUFx4f_ASAP7_75t_L g14026 ( 
.A(n_13674),
.Y(n_14026)
);

INVx2_ASAP7_75t_L g14027 ( 
.A(n_13767),
.Y(n_14027)
);

AND2x2_ASAP7_75t_L g14028 ( 
.A(n_13040),
.B(n_1230),
.Y(n_14028)
);

AND2x2_ASAP7_75t_L g14029 ( 
.A(n_12955),
.B(n_1231),
.Y(n_14029)
);

HB1xp67_ASAP7_75t_L g14030 ( 
.A(n_13732),
.Y(n_14030)
);

BUFx2_ASAP7_75t_L g14031 ( 
.A(n_13114),
.Y(n_14031)
);

AOI22xp5_ASAP7_75t_L g14032 ( 
.A1(n_12996),
.A2(n_1233),
.B1(n_1231),
.B2(n_1232),
.Y(n_14032)
);

INVx4_ASAP7_75t_L g14033 ( 
.A(n_13054),
.Y(n_14033)
);

AND2x2_ASAP7_75t_L g14034 ( 
.A(n_13564),
.B(n_1232),
.Y(n_14034)
);

AND2x2_ASAP7_75t_L g14035 ( 
.A(n_13733),
.B(n_1233),
.Y(n_14035)
);

NAND2xp5_ASAP7_75t_L g14036 ( 
.A(n_13743),
.B(n_1234),
.Y(n_14036)
);

BUFx6f_ASAP7_75t_L g14037 ( 
.A(n_13682),
.Y(n_14037)
);

INVx1_ASAP7_75t_L g14038 ( 
.A(n_13763),
.Y(n_14038)
);

INVx1_ASAP7_75t_L g14039 ( 
.A(n_13773),
.Y(n_14039)
);

INVx2_ASAP7_75t_L g14040 ( 
.A(n_13786),
.Y(n_14040)
);

INVx2_ASAP7_75t_L g14041 ( 
.A(n_13795),
.Y(n_14041)
);

NAND2xp5_ASAP7_75t_L g14042 ( 
.A(n_13811),
.B(n_1234),
.Y(n_14042)
);

BUFx2_ASAP7_75t_L g14043 ( 
.A(n_13186),
.Y(n_14043)
);

OR2x6_ASAP7_75t_L g14044 ( 
.A(n_13599),
.B(n_5835),
.Y(n_14044)
);

INVx1_ASAP7_75t_L g14045 ( 
.A(n_13842),
.Y(n_14045)
);

INVx1_ASAP7_75t_L g14046 ( 
.A(n_13851),
.Y(n_14046)
);

CKINVDCx5p33_ASAP7_75t_R g14047 ( 
.A(n_13087),
.Y(n_14047)
);

AND2x2_ASAP7_75t_L g14048 ( 
.A(n_13867),
.B(n_1235),
.Y(n_14048)
);

NOR2xp33_ASAP7_75t_L g14049 ( 
.A(n_13230),
.B(n_1235),
.Y(n_14049)
);

INVx2_ASAP7_75t_SL g14050 ( 
.A(n_12995),
.Y(n_14050)
);

INVx1_ASAP7_75t_L g14051 ( 
.A(n_13868),
.Y(n_14051)
);

INVx1_ASAP7_75t_L g14052 ( 
.A(n_12876),
.Y(n_14052)
);

NOR2xp67_ASAP7_75t_L g14053 ( 
.A(n_13410),
.B(n_1236),
.Y(n_14053)
);

NAND2xp5_ASAP7_75t_L g14054 ( 
.A(n_13800),
.B(n_1237),
.Y(n_14054)
);

A2O1A1Ixp33_ASAP7_75t_L g14055 ( 
.A1(n_13605),
.A2(n_1239),
.B(n_1237),
.C(n_1238),
.Y(n_14055)
);

INVx1_ASAP7_75t_L g14056 ( 
.A(n_13804),
.Y(n_14056)
);

INVx2_ASAP7_75t_L g14057 ( 
.A(n_13805),
.Y(n_14057)
);

CKINVDCx6p67_ASAP7_75t_R g14058 ( 
.A(n_13144),
.Y(n_14058)
);

INVx2_ASAP7_75t_L g14059 ( 
.A(n_13821),
.Y(n_14059)
);

NAND2xp5_ASAP7_75t_SL g14060 ( 
.A(n_13270),
.B(n_5837),
.Y(n_14060)
);

NAND2xp5_ASAP7_75t_L g14061 ( 
.A(n_13829),
.B(n_1238),
.Y(n_14061)
);

AND2x2_ASAP7_75t_L g14062 ( 
.A(n_13655),
.B(n_1239),
.Y(n_14062)
);

HB1xp67_ASAP7_75t_L g14063 ( 
.A(n_13840),
.Y(n_14063)
);

BUFx2_ASAP7_75t_L g14064 ( 
.A(n_13298),
.Y(n_14064)
);

NAND2xp5_ASAP7_75t_SL g14065 ( 
.A(n_12847),
.B(n_5838),
.Y(n_14065)
);

CKINVDCx8_ASAP7_75t_R g14066 ( 
.A(n_13682),
.Y(n_14066)
);

BUFx3_ASAP7_75t_L g14067 ( 
.A(n_13225),
.Y(n_14067)
);

NAND2xp5_ASAP7_75t_L g14068 ( 
.A(n_13861),
.B(n_1240),
.Y(n_14068)
);

INVx1_ASAP7_75t_L g14069 ( 
.A(n_13865),
.Y(n_14069)
);

INVx1_ASAP7_75t_L g14070 ( 
.A(n_13866),
.Y(n_14070)
);

NOR2xp67_ASAP7_75t_L g14071 ( 
.A(n_13410),
.B(n_1240),
.Y(n_14071)
);

BUFx3_ASAP7_75t_L g14072 ( 
.A(n_13700),
.Y(n_14072)
);

INVx1_ASAP7_75t_L g14073 ( 
.A(n_13884),
.Y(n_14073)
);

CKINVDCx5p33_ASAP7_75t_R g14074 ( 
.A(n_13889),
.Y(n_14074)
);

NAND2xp5_ASAP7_75t_L g14075 ( 
.A(n_13422),
.B(n_1241),
.Y(n_14075)
);

INVx1_ASAP7_75t_L g14076 ( 
.A(n_13013),
.Y(n_14076)
);

NAND2x1p5_ASAP7_75t_L g14077 ( 
.A(n_13395),
.B(n_5840),
.Y(n_14077)
);

OAI31xp33_ASAP7_75t_SL g14078 ( 
.A1(n_13246),
.A2(n_13038),
.A3(n_13741),
.B(n_12792),
.Y(n_14078)
);

INVx1_ASAP7_75t_L g14079 ( 
.A(n_13018),
.Y(n_14079)
);

NAND2xp5_ASAP7_75t_L g14080 ( 
.A(n_13445),
.B(n_1241),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_13455),
.B(n_1242),
.Y(n_14081)
);

AOI22x1_ASAP7_75t_L g14082 ( 
.A1(n_12851),
.A2(n_1245),
.B1(n_1243),
.B2(n_1244),
.Y(n_14082)
);

NAND2xp5_ASAP7_75t_SL g14083 ( 
.A(n_13520),
.B(n_5841),
.Y(n_14083)
);

INVx1_ASAP7_75t_L g14084 ( 
.A(n_13086),
.Y(n_14084)
);

NAND2xp5_ASAP7_75t_L g14085 ( 
.A(n_13175),
.B(n_1243),
.Y(n_14085)
);

NAND2xp5_ASAP7_75t_L g14086 ( 
.A(n_13248),
.B(n_1244),
.Y(n_14086)
);

NAND2xp5_ASAP7_75t_L g14087 ( 
.A(n_13269),
.B(n_13278),
.Y(n_14087)
);

AOI22x1_ASAP7_75t_L g14088 ( 
.A1(n_12904),
.A2(n_1247),
.B1(n_1245),
.B2(n_1246),
.Y(n_14088)
);

AND2x2_ASAP7_75t_L g14089 ( 
.A(n_13715),
.B(n_1246),
.Y(n_14089)
);

INVx2_ASAP7_75t_SL g14090 ( 
.A(n_12926),
.Y(n_14090)
);

NOR2xp67_ASAP7_75t_L g14091 ( 
.A(n_13410),
.B(n_1247),
.Y(n_14091)
);

A2O1A1Ixp33_ASAP7_75t_L g14092 ( 
.A1(n_13616),
.A2(n_13638),
.B(n_13661),
.C(n_13643),
.Y(n_14092)
);

INVx2_ASAP7_75t_L g14093 ( 
.A(n_12842),
.Y(n_14093)
);

INVx2_ASAP7_75t_L g14094 ( 
.A(n_13111),
.Y(n_14094)
);

BUFx2_ASAP7_75t_L g14095 ( 
.A(n_13377),
.Y(n_14095)
);

INVx3_ASAP7_75t_L g14096 ( 
.A(n_12969),
.Y(n_14096)
);

CKINVDCx14_ASAP7_75t_R g14097 ( 
.A(n_13401),
.Y(n_14097)
);

INVx2_ASAP7_75t_L g14098 ( 
.A(n_13132),
.Y(n_14098)
);

INVxp67_ASAP7_75t_L g14099 ( 
.A(n_13499),
.Y(n_14099)
);

NAND2xp5_ASAP7_75t_L g14100 ( 
.A(n_13321),
.B(n_1248),
.Y(n_14100)
);

CKINVDCx12_ASAP7_75t_R g14101 ( 
.A(n_13578),
.Y(n_14101)
);

INVx1_ASAP7_75t_L g14102 ( 
.A(n_13048),
.Y(n_14102)
);

NAND2xp5_ASAP7_75t_L g14103 ( 
.A(n_13335),
.B(n_1248),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_13062),
.Y(n_14104)
);

AND3x1_ASAP7_75t_SL g14105 ( 
.A(n_13468),
.B(n_1249),
.C(n_1250),
.Y(n_14105)
);

AND2x2_ASAP7_75t_L g14106 ( 
.A(n_13735),
.B(n_13747),
.Y(n_14106)
);

NAND2xp5_ASAP7_75t_L g14107 ( 
.A(n_13345),
.B(n_1250),
.Y(n_14107)
);

NAND2xp5_ASAP7_75t_L g14108 ( 
.A(n_13354),
.B(n_1251),
.Y(n_14108)
);

NAND2xp5_ASAP7_75t_L g14109 ( 
.A(n_13369),
.B(n_1252),
.Y(n_14109)
);

AND2x2_ASAP7_75t_L g14110 ( 
.A(n_13155),
.B(n_1252),
.Y(n_14110)
);

INVx1_ASAP7_75t_L g14111 ( 
.A(n_13068),
.Y(n_14111)
);

NAND2xp5_ASAP7_75t_L g14112 ( 
.A(n_13458),
.B(n_1253),
.Y(n_14112)
);

INVx3_ASAP7_75t_L g14113 ( 
.A(n_12969),
.Y(n_14113)
);

INVx1_ASAP7_75t_L g14114 ( 
.A(n_13084),
.Y(n_14114)
);

CKINVDCx16_ASAP7_75t_R g14115 ( 
.A(n_13080),
.Y(n_14115)
);

INVx1_ASAP7_75t_SL g14116 ( 
.A(n_13477),
.Y(n_14116)
);

INVx1_ASAP7_75t_L g14117 ( 
.A(n_13092),
.Y(n_14117)
);

INVx2_ASAP7_75t_L g14118 ( 
.A(n_13122),
.Y(n_14118)
);

AND2x2_ASAP7_75t_L g14119 ( 
.A(n_12813),
.B(n_1253),
.Y(n_14119)
);

INVxp67_ASAP7_75t_L g14120 ( 
.A(n_13555),
.Y(n_14120)
);

INVx2_ASAP7_75t_L g14121 ( 
.A(n_13125),
.Y(n_14121)
);

OAI22xp5_ASAP7_75t_SL g14122 ( 
.A1(n_13130),
.A2(n_1256),
.B1(n_1254),
.B2(n_1255),
.Y(n_14122)
);

AND2x4_ASAP7_75t_SL g14123 ( 
.A(n_13171),
.B(n_5842),
.Y(n_14123)
);

NAND2xp5_ASAP7_75t_L g14124 ( 
.A(n_13530),
.B(n_1254),
.Y(n_14124)
);

AND2x2_ASAP7_75t_L g14125 ( 
.A(n_13314),
.B(n_1255),
.Y(n_14125)
);

INVx1_ASAP7_75t_L g14126 ( 
.A(n_12971),
.Y(n_14126)
);

AND2x2_ASAP7_75t_L g14127 ( 
.A(n_13450),
.B(n_1256),
.Y(n_14127)
);

NAND2xp5_ASAP7_75t_L g14128 ( 
.A(n_13538),
.B(n_1257),
.Y(n_14128)
);

INVx1_ASAP7_75t_L g14129 ( 
.A(n_13042),
.Y(n_14129)
);

INVx1_ASAP7_75t_L g14130 ( 
.A(n_13145),
.Y(n_14130)
);

BUFx3_ASAP7_75t_L g14131 ( 
.A(n_13700),
.Y(n_14131)
);

OR2x2_ASAP7_75t_L g14132 ( 
.A(n_13182),
.B(n_1258),
.Y(n_14132)
);

INVx1_ASAP7_75t_L g14133 ( 
.A(n_13427),
.Y(n_14133)
);

INVx2_ASAP7_75t_L g14134 ( 
.A(n_13324),
.Y(n_14134)
);

AOI22xp33_ASAP7_75t_L g14135 ( 
.A1(n_12836),
.A2(n_13033),
.B1(n_13074),
.B2(n_13060),
.Y(n_14135)
);

BUFx2_ASAP7_75t_L g14136 ( 
.A(n_13395),
.Y(n_14136)
);

INVx2_ASAP7_75t_L g14137 ( 
.A(n_13326),
.Y(n_14137)
);

NAND2x1p5_ASAP7_75t_L g14138 ( 
.A(n_13395),
.B(n_5843),
.Y(n_14138)
);

A2O1A1Ixp33_ASAP7_75t_L g14139 ( 
.A1(n_13675),
.A2(n_1260),
.B(n_1258),
.C(n_1259),
.Y(n_14139)
);

INVx3_ASAP7_75t_L g14140 ( 
.A(n_13408),
.Y(n_14140)
);

A2O1A1Ixp33_ASAP7_75t_L g14141 ( 
.A1(n_13738),
.A2(n_1262),
.B(n_1259),
.C(n_1261),
.Y(n_14141)
);

NAND2xp5_ASAP7_75t_L g14142 ( 
.A(n_13543),
.B(n_13556),
.Y(n_14142)
);

INVx2_ASAP7_75t_L g14143 ( 
.A(n_13333),
.Y(n_14143)
);

NOR2xp33_ASAP7_75t_L g14144 ( 
.A(n_13267),
.B(n_1261),
.Y(n_14144)
);

AND2x2_ASAP7_75t_L g14145 ( 
.A(n_13557),
.B(n_13208),
.Y(n_14145)
);

CKINVDCx5p33_ASAP7_75t_R g14146 ( 
.A(n_13192),
.Y(n_14146)
);

AND2x2_ASAP7_75t_L g14147 ( 
.A(n_13233),
.B(n_1263),
.Y(n_14147)
);

NAND2xp5_ASAP7_75t_L g14148 ( 
.A(n_13339),
.B(n_1263),
.Y(n_14148)
);

BUFx2_ASAP7_75t_SL g14149 ( 
.A(n_12859),
.Y(n_14149)
);

CKINVDCx11_ASAP7_75t_R g14150 ( 
.A(n_13611),
.Y(n_14150)
);

NAND2xp5_ASAP7_75t_L g14151 ( 
.A(n_13364),
.B(n_1264),
.Y(n_14151)
);

NAND2xp5_ASAP7_75t_L g14152 ( 
.A(n_13391),
.B(n_1264),
.Y(n_14152)
);

XNOR2x1_ASAP7_75t_L g14153 ( 
.A(n_13487),
.B(n_13118),
.Y(n_14153)
);

BUFx12f_ASAP7_75t_L g14154 ( 
.A(n_13721),
.Y(n_14154)
);

OAI22xp5_ASAP7_75t_L g14155 ( 
.A1(n_13615),
.A2(n_1267),
.B1(n_1265),
.B2(n_1266),
.Y(n_14155)
);

INVx2_ASAP7_75t_L g14156 ( 
.A(n_13393),
.Y(n_14156)
);

INVx1_ASAP7_75t_L g14157 ( 
.A(n_13438),
.Y(n_14157)
);

NAND2xp5_ASAP7_75t_L g14158 ( 
.A(n_13247),
.B(n_1265),
.Y(n_14158)
);

NAND2xp5_ASAP7_75t_L g14159 ( 
.A(n_13301),
.B(n_1266),
.Y(n_14159)
);

AND2x2_ASAP7_75t_L g14160 ( 
.A(n_13310),
.B(n_1267),
.Y(n_14160)
);

AND2x4_ASAP7_75t_SL g14161 ( 
.A(n_13477),
.B(n_5844),
.Y(n_14161)
);

AOI22xp33_ASAP7_75t_L g14162 ( 
.A1(n_13830),
.A2(n_12841),
.B1(n_12922),
.B2(n_12903),
.Y(n_14162)
);

INVxp67_ASAP7_75t_L g14163 ( 
.A(n_13565),
.Y(n_14163)
);

NAND2xp5_ASAP7_75t_L g14164 ( 
.A(n_13474),
.B(n_1268),
.Y(n_14164)
);

INVx1_ASAP7_75t_L g14165 ( 
.A(n_13488),
.Y(n_14165)
);

NAND2xp5_ASAP7_75t_L g14166 ( 
.A(n_13480),
.B(n_1269),
.Y(n_14166)
);

AND2x2_ASAP7_75t_L g14167 ( 
.A(n_12864),
.B(n_1269),
.Y(n_14167)
);

INVx2_ASAP7_75t_L g14168 ( 
.A(n_13000),
.Y(n_14168)
);

INVx4_ASAP7_75t_L g14169 ( 
.A(n_12993),
.Y(n_14169)
);

INVx2_ASAP7_75t_L g14170 ( 
.A(n_13294),
.Y(n_14170)
);

CKINVDCx11_ASAP7_75t_R g14171 ( 
.A(n_13623),
.Y(n_14171)
);

AND2x2_ASAP7_75t_L g14172 ( 
.A(n_13478),
.B(n_1270),
.Y(n_14172)
);

AND2x2_ASAP7_75t_L g14173 ( 
.A(n_13392),
.B(n_1270),
.Y(n_14173)
);

NOR2x1_ASAP7_75t_L g14174 ( 
.A(n_12805),
.B(n_1271),
.Y(n_14174)
);

INVx1_ASAP7_75t_L g14175 ( 
.A(n_13593),
.Y(n_14175)
);

NOR2xp33_ASAP7_75t_L g14176 ( 
.A(n_13061),
.B(n_1271),
.Y(n_14176)
);

AND3x1_ASAP7_75t_SL g14177 ( 
.A(n_13274),
.B(n_1272),
.C(n_1273),
.Y(n_14177)
);

AND2x2_ASAP7_75t_L g14178 ( 
.A(n_13110),
.B(n_1272),
.Y(n_14178)
);

INVx2_ASAP7_75t_L g14179 ( 
.A(n_13313),
.Y(n_14179)
);

NAND2xp5_ASAP7_75t_L g14180 ( 
.A(n_13510),
.B(n_1273),
.Y(n_14180)
);

INVx1_ASAP7_75t_L g14181 ( 
.A(n_13577),
.Y(n_14181)
);

AND2x2_ASAP7_75t_L g14182 ( 
.A(n_13203),
.B(n_13237),
.Y(n_14182)
);

AND2x2_ASAP7_75t_L g14183 ( 
.A(n_12819),
.B(n_1274),
.Y(n_14183)
);

NAND2xp5_ASAP7_75t_L g14184 ( 
.A(n_12835),
.B(n_1274),
.Y(n_14184)
);

NAND2xp5_ASAP7_75t_L g14185 ( 
.A(n_12818),
.B(n_1275),
.Y(n_14185)
);

INVxp67_ASAP7_75t_L g14186 ( 
.A(n_13073),
.Y(n_14186)
);

INVx1_ASAP7_75t_L g14187 ( 
.A(n_13571),
.Y(n_14187)
);

INVx1_ASAP7_75t_L g14188 ( 
.A(n_13165),
.Y(n_14188)
);

NOR2xp33_ASAP7_75t_L g14189 ( 
.A(n_13421),
.B(n_1275),
.Y(n_14189)
);

NOR2xp33_ASAP7_75t_L g14190 ( 
.A(n_12800),
.B(n_1276),
.Y(n_14190)
);

NAND2xp5_ASAP7_75t_L g14191 ( 
.A(n_12885),
.B(n_1276),
.Y(n_14191)
);

NAND2xp5_ASAP7_75t_L g14192 ( 
.A(n_12940),
.B(n_1277),
.Y(n_14192)
);

BUFx3_ASAP7_75t_L g14193 ( 
.A(n_13721),
.Y(n_14193)
);

INVx1_ASAP7_75t_L g14194 ( 
.A(n_13749),
.Y(n_14194)
);

INVx2_ASAP7_75t_L g14195 ( 
.A(n_13137),
.Y(n_14195)
);

INVx3_ASAP7_75t_L g14196 ( 
.A(n_13408),
.Y(n_14196)
);

NAND2xp5_ASAP7_75t_L g14197 ( 
.A(n_12853),
.B(n_1278),
.Y(n_14197)
);

INVx1_ASAP7_75t_L g14198 ( 
.A(n_12952),
.Y(n_14198)
);

BUFx10_ASAP7_75t_L g14199 ( 
.A(n_13726),
.Y(n_14199)
);

AOI22xp33_ASAP7_75t_L g14200 ( 
.A1(n_12923),
.A2(n_12943),
.B1(n_13755),
.B2(n_13281),
.Y(n_14200)
);

AND2x6_ASAP7_75t_L g14201 ( 
.A(n_12849),
.B(n_5845),
.Y(n_14201)
);

INVx1_ASAP7_75t_L g14202 ( 
.A(n_12954),
.Y(n_14202)
);

NAND2xp5_ASAP7_75t_L g14203 ( 
.A(n_12855),
.B(n_1278),
.Y(n_14203)
);

NAND2xp5_ASAP7_75t_L g14204 ( 
.A(n_12880),
.B(n_1279),
.Y(n_14204)
);

BUFx2_ASAP7_75t_L g14205 ( 
.A(n_13304),
.Y(n_14205)
);

NAND2xp5_ASAP7_75t_L g14206 ( 
.A(n_12883),
.B(n_1279),
.Y(n_14206)
);

NAND2xp5_ASAP7_75t_L g14207 ( 
.A(n_12810),
.B(n_1280),
.Y(n_14207)
);

INVx2_ASAP7_75t_L g14208 ( 
.A(n_12822),
.Y(n_14208)
);

NAND2xp5_ASAP7_75t_SL g14209 ( 
.A(n_13570),
.B(n_5846),
.Y(n_14209)
);

OAI22xp5_ASAP7_75t_SL g14210 ( 
.A1(n_13148),
.A2(n_1282),
.B1(n_1280),
.B2(n_1281),
.Y(n_14210)
);

AND3x1_ASAP7_75t_SL g14211 ( 
.A(n_13031),
.B(n_1281),
.C(n_1282),
.Y(n_14211)
);

INVx1_ASAP7_75t_L g14212 ( 
.A(n_12962),
.Y(n_14212)
);

INVx1_ASAP7_75t_L g14213 ( 
.A(n_12964),
.Y(n_14213)
);

AND2x6_ASAP7_75t_L g14214 ( 
.A(n_13121),
.B(n_5847),
.Y(n_14214)
);

INVxp67_ASAP7_75t_L g14215 ( 
.A(n_12846),
.Y(n_14215)
);

INVx1_ASAP7_75t_L g14216 ( 
.A(n_12977),
.Y(n_14216)
);

INVx1_ASAP7_75t_L g14217 ( 
.A(n_12950),
.Y(n_14217)
);

INVxp67_ASAP7_75t_SL g14218 ( 
.A(n_13651),
.Y(n_14218)
);

BUFx3_ASAP7_75t_L g14219 ( 
.A(n_13726),
.Y(n_14219)
);

BUFx6f_ASAP7_75t_L g14220 ( 
.A(n_13809),
.Y(n_14220)
);

OR2x2_ASAP7_75t_L g14221 ( 
.A(n_13900),
.B(n_1283),
.Y(n_14221)
);

AND2x2_ASAP7_75t_L g14222 ( 
.A(n_13646),
.B(n_1283),
.Y(n_14222)
);

INVx1_ASAP7_75t_L g14223 ( 
.A(n_12967),
.Y(n_14223)
);

NAND2xp5_ASAP7_75t_L g14224 ( 
.A(n_12815),
.B(n_1285),
.Y(n_14224)
);

INVx6_ASAP7_75t_L g14225 ( 
.A(n_13809),
.Y(n_14225)
);

NAND2xp5_ASAP7_75t_L g14226 ( 
.A(n_13622),
.B(n_1286),
.Y(n_14226)
);

INVx1_ASAP7_75t_L g14227 ( 
.A(n_12976),
.Y(n_14227)
);

INVx2_ASAP7_75t_L g14228 ( 
.A(n_12913),
.Y(n_14228)
);

NAND2xp5_ASAP7_75t_L g14229 ( 
.A(n_13624),
.B(n_1286),
.Y(n_14229)
);

NAND2xp5_ASAP7_75t_L g14230 ( 
.A(n_13626),
.B(n_1287),
.Y(n_14230)
);

NAND2xp5_ASAP7_75t_L g14231 ( 
.A(n_13629),
.B(n_1287),
.Y(n_14231)
);

CKINVDCx5p33_ASAP7_75t_R g14232 ( 
.A(n_13010),
.Y(n_14232)
);

INVx2_ASAP7_75t_L g14233 ( 
.A(n_12936),
.Y(n_14233)
);

NAND2xp5_ASAP7_75t_L g14234 ( 
.A(n_13632),
.B(n_1288),
.Y(n_14234)
);

INVx1_ASAP7_75t_L g14235 ( 
.A(n_12986),
.Y(n_14235)
);

CKINVDCx20_ASAP7_75t_R g14236 ( 
.A(n_12981),
.Y(n_14236)
);

CKINVDCx5p33_ASAP7_75t_R g14237 ( 
.A(n_13290),
.Y(n_14237)
);

NOR2xp33_ASAP7_75t_L g14238 ( 
.A(n_13604),
.B(n_1288),
.Y(n_14238)
);

INVx2_ASAP7_75t_L g14239 ( 
.A(n_12991),
.Y(n_14239)
);

INVx1_ASAP7_75t_L g14240 ( 
.A(n_12990),
.Y(n_14240)
);

CKINVDCx11_ASAP7_75t_R g14241 ( 
.A(n_13845),
.Y(n_14241)
);

INVx1_ASAP7_75t_L g14242 ( 
.A(n_12999),
.Y(n_14242)
);

NAND2xp5_ASAP7_75t_L g14243 ( 
.A(n_13634),
.B(n_1289),
.Y(n_14243)
);

INVx1_ASAP7_75t_L g14244 ( 
.A(n_13007),
.Y(n_14244)
);

AND2x2_ASAP7_75t_L g14245 ( 
.A(n_13678),
.B(n_1289),
.Y(n_14245)
);

INVx1_ASAP7_75t_L g14246 ( 
.A(n_13016),
.Y(n_14246)
);

INVx1_ASAP7_75t_L g14247 ( 
.A(n_13017),
.Y(n_14247)
);

NAND2xp5_ASAP7_75t_L g14248 ( 
.A(n_13637),
.B(n_1290),
.Y(n_14248)
);

INVx1_ASAP7_75t_L g14249 ( 
.A(n_13024),
.Y(n_14249)
);

AOI211xp5_ASAP7_75t_L g14250 ( 
.A1(n_13426),
.A2(n_1292),
.B(n_1290),
.C(n_1291),
.Y(n_14250)
);

INVx4_ASAP7_75t_L g14251 ( 
.A(n_12993),
.Y(n_14251)
);

INVx3_ASAP7_75t_L g14252 ( 
.A(n_13012),
.Y(n_14252)
);

NAND2xp5_ASAP7_75t_L g14253 ( 
.A(n_13640),
.B(n_1291),
.Y(n_14253)
);

NAND2xp5_ASAP7_75t_L g14254 ( 
.A(n_13654),
.B(n_1292),
.Y(n_14254)
);

INVx4_ASAP7_75t_L g14255 ( 
.A(n_13012),
.Y(n_14255)
);

INVx1_ASAP7_75t_L g14256 ( 
.A(n_13026),
.Y(n_14256)
);

HB1xp67_ASAP7_75t_L g14257 ( 
.A(n_13356),
.Y(n_14257)
);

NAND2xp5_ASAP7_75t_L g14258 ( 
.A(n_13659),
.B(n_1293),
.Y(n_14258)
);

NAND2xp5_ASAP7_75t_L g14259 ( 
.A(n_13664),
.B(n_1293),
.Y(n_14259)
);

NAND2xp5_ASAP7_75t_L g14260 ( 
.A(n_13667),
.B(n_1294),
.Y(n_14260)
);

NAND2xp5_ASAP7_75t_L g14261 ( 
.A(n_13668),
.B(n_1294),
.Y(n_14261)
);

INVx2_ASAP7_75t_L g14262 ( 
.A(n_13019),
.Y(n_14262)
);

INVx1_ASAP7_75t_L g14263 ( 
.A(n_13030),
.Y(n_14263)
);

NAND2xp5_ASAP7_75t_SL g14264 ( 
.A(n_13399),
.B(n_5849),
.Y(n_14264)
);

AND2x2_ASAP7_75t_L g14265 ( 
.A(n_13684),
.B(n_1295),
.Y(n_14265)
);

NAND2xp5_ASAP7_75t_SL g14266 ( 
.A(n_12828),
.B(n_5851),
.Y(n_14266)
);

INVx2_ASAP7_75t_L g14267 ( 
.A(n_13607),
.Y(n_14267)
);

INVx1_ASAP7_75t_L g14268 ( 
.A(n_13032),
.Y(n_14268)
);

AND2x4_ASAP7_75t_L g14269 ( 
.A(n_13547),
.B(n_5852),
.Y(n_14269)
);

NAND2xp5_ASAP7_75t_L g14270 ( 
.A(n_13673),
.B(n_13677),
.Y(n_14270)
);

AND2x2_ASAP7_75t_L g14271 ( 
.A(n_13742),
.B(n_1295),
.Y(n_14271)
);

INVx1_ASAP7_75t_L g14272 ( 
.A(n_13044),
.Y(n_14272)
);

AND2x2_ASAP7_75t_L g14273 ( 
.A(n_13753),
.B(n_1296),
.Y(n_14273)
);

BUFx2_ASAP7_75t_L g14274 ( 
.A(n_13639),
.Y(n_14274)
);

INVx2_ASAP7_75t_L g14275 ( 
.A(n_13716),
.Y(n_14275)
);

INVx2_ASAP7_75t_L g14276 ( 
.A(n_13730),
.Y(n_14276)
);

AND3x1_ASAP7_75t_SL g14277 ( 
.A(n_12845),
.B(n_1297),
.C(n_1298),
.Y(n_14277)
);

AND2x6_ASAP7_75t_L g14278 ( 
.A(n_13688),
.B(n_5853),
.Y(n_14278)
);

OAI21x1_ASAP7_75t_L g14279 ( 
.A1(n_13009),
.A2(n_5856),
.B(n_5855),
.Y(n_14279)
);

NAND2xp5_ASAP7_75t_L g14280 ( 
.A(n_13680),
.B(n_1297),
.Y(n_14280)
);

CKINVDCx20_ASAP7_75t_R g14281 ( 
.A(n_13710),
.Y(n_14281)
);

INVxp67_ASAP7_75t_L g14282 ( 
.A(n_12848),
.Y(n_14282)
);

INVx4_ASAP7_75t_L g14283 ( 
.A(n_13184),
.Y(n_14283)
);

AND2x4_ASAP7_75t_L g14284 ( 
.A(n_12862),
.B(n_13836),
.Y(n_14284)
);

INVx2_ASAP7_75t_L g14285 ( 
.A(n_13083),
.Y(n_14285)
);

INVx1_ASAP7_75t_L g14286 ( 
.A(n_13050),
.Y(n_14286)
);

INVx2_ASAP7_75t_L g14287 ( 
.A(n_13136),
.Y(n_14287)
);

INVx2_ASAP7_75t_L g14288 ( 
.A(n_13157),
.Y(n_14288)
);

AND2x2_ASAP7_75t_L g14289 ( 
.A(n_13817),
.B(n_13818),
.Y(n_14289)
);

AND2x2_ASAP7_75t_L g14290 ( 
.A(n_13430),
.B(n_1298),
.Y(n_14290)
);

NOR2xp33_ASAP7_75t_R g14291 ( 
.A(n_13887),
.B(n_1299),
.Y(n_14291)
);

AOI22xp5_ASAP7_75t_L g14292 ( 
.A1(n_13357),
.A2(n_12821),
.B1(n_13213),
.B2(n_12799),
.Y(n_14292)
);

NAND2xp5_ASAP7_75t_L g14293 ( 
.A(n_13694),
.B(n_1299),
.Y(n_14293)
);

INVx1_ASAP7_75t_L g14294 ( 
.A(n_13058),
.Y(n_14294)
);

NAND2xp5_ASAP7_75t_L g14295 ( 
.A(n_13696),
.B(n_1300),
.Y(n_14295)
);

INVx2_ASAP7_75t_L g14296 ( 
.A(n_13209),
.Y(n_14296)
);

NAND2xp5_ASAP7_75t_L g14297 ( 
.A(n_13717),
.B(n_1301),
.Y(n_14297)
);

NAND2xp5_ASAP7_75t_L g14298 ( 
.A(n_13737),
.B(n_1301),
.Y(n_14298)
);

INVx2_ASAP7_75t_L g14299 ( 
.A(n_13271),
.Y(n_14299)
);

OAI22xp33_ASAP7_75t_L g14300 ( 
.A1(n_12869),
.A2(n_1304),
.B1(n_1302),
.B2(n_1303),
.Y(n_14300)
);

NAND2xp5_ASAP7_75t_L g14301 ( 
.A(n_13744),
.B(n_1302),
.Y(n_14301)
);

BUFx2_ASAP7_75t_L g14302 ( 
.A(n_13285),
.Y(n_14302)
);

AND3x1_ASAP7_75t_SL g14303 ( 
.A(n_12901),
.B(n_1305),
.C(n_1306),
.Y(n_14303)
);

NAND2xp5_ASAP7_75t_L g14304 ( 
.A(n_13760),
.B(n_1305),
.Y(n_14304)
);

INVx3_ASAP7_75t_L g14305 ( 
.A(n_13184),
.Y(n_14305)
);

AND2x2_ASAP7_75t_L g14306 ( 
.A(n_13081),
.B(n_1306),
.Y(n_14306)
);

BUFx6f_ASAP7_75t_L g14307 ( 
.A(n_13250),
.Y(n_14307)
);

BUFx6f_ASAP7_75t_L g14308 ( 
.A(n_13250),
.Y(n_14308)
);

NAND2xp5_ASAP7_75t_SL g14309 ( 
.A(n_13695),
.B(n_5857),
.Y(n_14309)
);

INVx1_ASAP7_75t_L g14310 ( 
.A(n_13063),
.Y(n_14310)
);

NAND2xp5_ASAP7_75t_SL g14311 ( 
.A(n_13149),
.B(n_13193),
.Y(n_14311)
);

INVx1_ASAP7_75t_L g14312 ( 
.A(n_13067),
.Y(n_14312)
);

NAND2xp5_ASAP7_75t_L g14313 ( 
.A(n_13761),
.B(n_1307),
.Y(n_14313)
);

INVx2_ASAP7_75t_L g14314 ( 
.A(n_13338),
.Y(n_14314)
);

INVx2_ASAP7_75t_L g14315 ( 
.A(n_13308),
.Y(n_14315)
);

AND2x2_ASAP7_75t_SL g14316 ( 
.A(n_13567),
.B(n_1307),
.Y(n_14316)
);

INVx2_ASAP7_75t_L g14317 ( 
.A(n_13331),
.Y(n_14317)
);

INVx3_ASAP7_75t_L g14318 ( 
.A(n_13331),
.Y(n_14318)
);

INVx1_ASAP7_75t_L g14319 ( 
.A(n_13071),
.Y(n_14319)
);

AND2x2_ASAP7_75t_L g14320 ( 
.A(n_12894),
.B(n_1308),
.Y(n_14320)
);

NAND2xp5_ASAP7_75t_L g14321 ( 
.A(n_13766),
.B(n_1308),
.Y(n_14321)
);

NAND2xp5_ASAP7_75t_L g14322 ( 
.A(n_13779),
.B(n_1309),
.Y(n_14322)
);

CKINVDCx16_ASAP7_75t_R g14323 ( 
.A(n_13370),
.Y(n_14323)
);

INVx2_ASAP7_75t_L g14324 ( 
.A(n_13787),
.Y(n_14324)
);

INVx2_ASAP7_75t_L g14325 ( 
.A(n_13788),
.Y(n_14325)
);

BUFx2_ASAP7_75t_L g14326 ( 
.A(n_13505),
.Y(n_14326)
);

CKINVDCx5p33_ASAP7_75t_R g14327 ( 
.A(n_13388),
.Y(n_14327)
);

NOR2xp33_ASAP7_75t_L g14328 ( 
.A(n_13660),
.B(n_1309),
.Y(n_14328)
);

NAND2xp5_ASAP7_75t_L g14329 ( 
.A(n_13813),
.B(n_1310),
.Y(n_14329)
);

INVx1_ASAP7_75t_L g14330 ( 
.A(n_13097),
.Y(n_14330)
);

NAND2xp5_ASAP7_75t_L g14331 ( 
.A(n_13819),
.B(n_1310),
.Y(n_14331)
);

AND2x2_ASAP7_75t_L g14332 ( 
.A(n_13525),
.B(n_1311),
.Y(n_14332)
);

AND2x2_ASAP7_75t_L g14333 ( 
.A(n_13841),
.B(n_1311),
.Y(n_14333)
);

NAND2xp5_ASAP7_75t_L g14334 ( 
.A(n_13844),
.B(n_13853),
.Y(n_14334)
);

NOR2xp33_ASAP7_75t_R g14335 ( 
.A(n_13195),
.B(n_1312),
.Y(n_14335)
);

CKINVDCx20_ASAP7_75t_R g14336 ( 
.A(n_13454),
.Y(n_14336)
);

INVx2_ASAP7_75t_L g14337 ( 
.A(n_13857),
.Y(n_14337)
);

OAI22xp5_ASAP7_75t_SL g14338 ( 
.A1(n_13390),
.A2(n_1314),
.B1(n_1312),
.B2(n_1313),
.Y(n_14338)
);

HB1xp67_ASAP7_75t_L g14339 ( 
.A(n_13729),
.Y(n_14339)
);

AOI22xp33_ASAP7_75t_L g14340 ( 
.A1(n_13360),
.A2(n_1316),
.B1(n_1313),
.B2(n_1315),
.Y(n_14340)
);

INVx1_ASAP7_75t_SL g14341 ( 
.A(n_13431),
.Y(n_14341)
);

AO22x1_ASAP7_75t_L g14342 ( 
.A1(n_13318),
.A2(n_1317),
.B1(n_1315),
.B2(n_1316),
.Y(n_14342)
);

NAND2xp5_ASAP7_75t_SL g14343 ( 
.A(n_13153),
.B(n_5858),
.Y(n_14343)
);

INVx1_ASAP7_75t_L g14344 ( 
.A(n_13099),
.Y(n_14344)
);

INVx1_ASAP7_75t_L g14345 ( 
.A(n_13108),
.Y(n_14345)
);

AND2x2_ASAP7_75t_L g14346 ( 
.A(n_13859),
.B(n_1317),
.Y(n_14346)
);

INVx2_ASAP7_75t_L g14347 ( 
.A(n_13864),
.Y(n_14347)
);

A2O1A1Ixp33_ASAP7_75t_L g14348 ( 
.A1(n_13758),
.A2(n_1320),
.B(n_1318),
.C(n_1319),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_13129),
.Y(n_14349)
);

CKINVDCx5p33_ASAP7_75t_R g14350 ( 
.A(n_13490),
.Y(n_14350)
);

AND2x2_ASAP7_75t_L g14351 ( 
.A(n_13874),
.B(n_1318),
.Y(n_14351)
);

AND2x2_ASAP7_75t_L g14352 ( 
.A(n_13878),
.B(n_13880),
.Y(n_14352)
);

AOI22xp5_ASAP7_75t_L g14353 ( 
.A1(n_12966),
.A2(n_1321),
.B1(n_1319),
.B2(n_1320),
.Y(n_14353)
);

AND2x2_ASAP7_75t_L g14354 ( 
.A(n_13886),
.B(n_1321),
.Y(n_14354)
);

AND2x2_ASAP7_75t_L g14355 ( 
.A(n_13898),
.B(n_1322),
.Y(n_14355)
);

INVx3_ASAP7_75t_SL g14356 ( 
.A(n_13046),
.Y(n_14356)
);

INVx1_ASAP7_75t_L g14357 ( 
.A(n_13131),
.Y(n_14357)
);

CKINVDCx11_ASAP7_75t_R g14358 ( 
.A(n_13119),
.Y(n_14358)
);

NAND2xp5_ASAP7_75t_SL g14359 ( 
.A(n_12838),
.B(n_5860),
.Y(n_14359)
);

NAND2xp5_ASAP7_75t_L g14360 ( 
.A(n_13670),
.B(n_13671),
.Y(n_14360)
);

INVx2_ASAP7_75t_L g14361 ( 
.A(n_13135),
.Y(n_14361)
);

AND2x2_ASAP7_75t_L g14362 ( 
.A(n_13625),
.B(n_1323),
.Y(n_14362)
);

INVx1_ASAP7_75t_L g14363 ( 
.A(n_13142),
.Y(n_14363)
);

AND2x2_ASAP7_75t_L g14364 ( 
.A(n_13691),
.B(n_1323),
.Y(n_14364)
);

INVx2_ASAP7_75t_L g14365 ( 
.A(n_13143),
.Y(n_14365)
);

BUFx12f_ASAP7_75t_L g14366 ( 
.A(n_13754),
.Y(n_14366)
);

AND2x4_ASAP7_75t_L g14367 ( 
.A(n_13434),
.B(n_13470),
.Y(n_14367)
);

INVx1_ASAP7_75t_L g14368 ( 
.A(n_12900),
.Y(n_14368)
);

INVx1_ASAP7_75t_L g14369 ( 
.A(n_12912),
.Y(n_14369)
);

NAND2xp5_ASAP7_75t_L g14370 ( 
.A(n_13686),
.B(n_1324),
.Y(n_14370)
);

NAND2x1p5_ASAP7_75t_L g14371 ( 
.A(n_13036),
.B(n_5861),
.Y(n_14371)
);

NAND2xp5_ASAP7_75t_L g14372 ( 
.A(n_13707),
.B(n_1324),
.Y(n_14372)
);

INVx1_ASAP7_75t_L g14373 ( 
.A(n_12831),
.Y(n_14373)
);

NAND2xp5_ASAP7_75t_L g14374 ( 
.A(n_13709),
.B(n_1325),
.Y(n_14374)
);

AND2x2_ASAP7_75t_L g14375 ( 
.A(n_13722),
.B(n_1325),
.Y(n_14375)
);

NAND2x1p5_ASAP7_75t_L g14376 ( 
.A(n_13630),
.B(n_5862),
.Y(n_14376)
);

CKINVDCx6p67_ASAP7_75t_R g14377 ( 
.A(n_13494),
.Y(n_14377)
);

INVx1_ASAP7_75t_L g14378 ( 
.A(n_12933),
.Y(n_14378)
);

NAND2xp5_ASAP7_75t_L g14379 ( 
.A(n_13724),
.B(n_1326),
.Y(n_14379)
);

INVx1_ASAP7_75t_L g14380 ( 
.A(n_12930),
.Y(n_14380)
);

NAND2xp5_ASAP7_75t_SL g14381 ( 
.A(n_13790),
.B(n_5863),
.Y(n_14381)
);

INVx1_ASAP7_75t_L g14382 ( 
.A(n_12941),
.Y(n_14382)
);

NAND2xp5_ASAP7_75t_L g14383 ( 
.A(n_13736),
.B(n_1326),
.Y(n_14383)
);

BUFx3_ASAP7_75t_L g14384 ( 
.A(n_13431),
.Y(n_14384)
);

NAND2x1p5_ASAP7_75t_L g14385 ( 
.A(n_13720),
.B(n_5864),
.Y(n_14385)
);

AND2x2_ASAP7_75t_L g14386 ( 
.A(n_13815),
.B(n_1327),
.Y(n_14386)
);

INVx1_ASAP7_75t_SL g14387 ( 
.A(n_13432),
.Y(n_14387)
);

HB1xp67_ASAP7_75t_L g14388 ( 
.A(n_13170),
.Y(n_14388)
);

OAI22xp5_ASAP7_75t_SL g14389 ( 
.A1(n_13210),
.A2(n_1330),
.B1(n_1328),
.B2(n_1329),
.Y(n_14389)
);

AND2x2_ASAP7_75t_L g14390 ( 
.A(n_12884),
.B(n_1328),
.Y(n_14390)
);

NAND2xp33_ASAP7_75t_L g14391 ( 
.A(n_12829),
.B(n_13448),
.Y(n_14391)
);

AOI22xp5_ASAP7_75t_L g14392 ( 
.A1(n_13693),
.A2(n_1331),
.B1(n_1329),
.B2(n_1330),
.Y(n_14392)
);

AND2x2_ASAP7_75t_L g14393 ( 
.A(n_13123),
.B(n_1331),
.Y(n_14393)
);

INVx1_ASAP7_75t_L g14394 ( 
.A(n_12953),
.Y(n_14394)
);

INVx3_ASAP7_75t_L g14395 ( 
.A(n_13432),
.Y(n_14395)
);

AND2x2_ASAP7_75t_L g14396 ( 
.A(n_13133),
.B(n_1332),
.Y(n_14396)
);

NAND2xp5_ASAP7_75t_SL g14397 ( 
.A(n_13166),
.B(n_5866),
.Y(n_14397)
);

NAND2xp5_ASAP7_75t_L g14398 ( 
.A(n_13801),
.B(n_1332),
.Y(n_14398)
);

INVx1_ASAP7_75t_L g14399 ( 
.A(n_12861),
.Y(n_14399)
);

INVx1_ASAP7_75t_L g14400 ( 
.A(n_12877),
.Y(n_14400)
);

OAI22xp5_ASAP7_75t_SL g14401 ( 
.A1(n_13088),
.A2(n_1335),
.B1(n_1333),
.B2(n_1334),
.Y(n_14401)
);

NAND2xp5_ASAP7_75t_L g14402 ( 
.A(n_13823),
.B(n_1333),
.Y(n_14402)
);

OAI22xp5_ASAP7_75t_L g14403 ( 
.A1(n_13725),
.A2(n_1336),
.B1(n_1334),
.B2(n_1335),
.Y(n_14403)
);

AOI22xp33_ASAP7_75t_L g14404 ( 
.A1(n_12873),
.A2(n_1338),
.B1(n_1336),
.B2(n_1337),
.Y(n_14404)
);

BUFx12f_ASAP7_75t_L g14405 ( 
.A(n_13494),
.Y(n_14405)
);

CKINVDCx5p33_ASAP7_75t_R g14406 ( 
.A(n_13146),
.Y(n_14406)
);

INVx1_ASAP7_75t_L g14407 ( 
.A(n_12958),
.Y(n_14407)
);

INVx1_ASAP7_75t_L g14408 ( 
.A(n_13177),
.Y(n_14408)
);

BUFx2_ASAP7_75t_L g14409 ( 
.A(n_13774),
.Y(n_14409)
);

INVx1_ASAP7_75t_SL g14410 ( 
.A(n_12858),
.Y(n_14410)
);

INVx1_ASAP7_75t_L g14411 ( 
.A(n_13589),
.Y(n_14411)
);

INVx1_ASAP7_75t_L g14412 ( 
.A(n_13053),
.Y(n_14412)
);

AND2x2_ASAP7_75t_L g14413 ( 
.A(n_13167),
.B(n_1337),
.Y(n_14413)
);

NAND2xp5_ASAP7_75t_L g14414 ( 
.A(n_13879),
.B(n_1338),
.Y(n_14414)
);

INVx1_ASAP7_75t_L g14415 ( 
.A(n_13219),
.Y(n_14415)
);

INVx1_ASAP7_75t_L g14416 ( 
.A(n_12872),
.Y(n_14416)
);

INVx1_ASAP7_75t_L g14417 ( 
.A(n_12839),
.Y(n_14417)
);

INVx1_ASAP7_75t_L g14418 ( 
.A(n_12896),
.Y(n_14418)
);

INVx2_ASAP7_75t_SL g14419 ( 
.A(n_13552),
.Y(n_14419)
);

INVx2_ASAP7_75t_L g14420 ( 
.A(n_12902),
.Y(n_14420)
);

AOI22xp33_ASAP7_75t_L g14421 ( 
.A1(n_13279),
.A2(n_1341),
.B1(n_1339),
.B2(n_1340),
.Y(n_14421)
);

INVx2_ASAP7_75t_L g14422 ( 
.A(n_12929),
.Y(n_14422)
);

INVx2_ASAP7_75t_L g14423 ( 
.A(n_13877),
.Y(n_14423)
);

HB1xp67_ASAP7_75t_L g14424 ( 
.A(n_13358),
.Y(n_14424)
);

INVx1_ASAP7_75t_L g14425 ( 
.A(n_13069),
.Y(n_14425)
);

AND2x4_ASAP7_75t_L g14426 ( 
.A(n_12804),
.B(n_13759),
.Y(n_14426)
);

NAND2xp5_ASAP7_75t_SL g14427 ( 
.A(n_13579),
.B(n_5867),
.Y(n_14427)
);

INVx1_ASAP7_75t_L g14428 ( 
.A(n_13679),
.Y(n_14428)
);

OR2x6_ASAP7_75t_L g14429 ( 
.A(n_13774),
.B(n_5869),
.Y(n_14429)
);

NAND2xp5_ASAP7_75t_L g14430 ( 
.A(n_13901),
.B(n_13173),
.Y(n_14430)
);

AND2x2_ASAP7_75t_L g14431 ( 
.A(n_13189),
.B(n_1339),
.Y(n_14431)
);

AND2x2_ASAP7_75t_L g14432 ( 
.A(n_13224),
.B(n_1340),
.Y(n_14432)
);

INVx2_ASAP7_75t_SL g14433 ( 
.A(n_13552),
.Y(n_14433)
);

BUFx2_ASAP7_75t_L g14434 ( 
.A(n_13791),
.Y(n_14434)
);

AND2x2_ASAP7_75t_L g14435 ( 
.A(n_13275),
.B(n_1341),
.Y(n_14435)
);

CKINVDCx5p33_ASAP7_75t_R g14436 ( 
.A(n_13234),
.Y(n_14436)
);

CKINVDCx5p33_ASAP7_75t_R g14437 ( 
.A(n_13299),
.Y(n_14437)
);

HB1xp67_ASAP7_75t_L g14438 ( 
.A(n_13587),
.Y(n_14438)
);

AND2x2_ASAP7_75t_L g14439 ( 
.A(n_13297),
.B(n_1342),
.Y(n_14439)
);

INVx1_ASAP7_75t_L g14440 ( 
.A(n_13820),
.Y(n_14440)
);

NAND2xp5_ASAP7_75t_SL g14441 ( 
.A(n_12907),
.B(n_5870),
.Y(n_14441)
);

HB1xp67_ASAP7_75t_L g14442 ( 
.A(n_13425),
.Y(n_14442)
);

OR2x2_ASAP7_75t_L g14443 ( 
.A(n_13194),
.B(n_1342),
.Y(n_14443)
);

NAND2xp5_ASAP7_75t_SL g14444 ( 
.A(n_12937),
.B(n_5871),
.Y(n_14444)
);

OAI21xp5_ASAP7_75t_L g14445 ( 
.A1(n_13190),
.A2(n_12832),
.B(n_13035),
.Y(n_14445)
);

INVx2_ASAP7_75t_L g14446 ( 
.A(n_13862),
.Y(n_14446)
);

BUFx2_ASAP7_75t_L g14447 ( 
.A(n_13792),
.Y(n_14447)
);

NAND2xp5_ASAP7_75t_L g14448 ( 
.A(n_13216),
.B(n_1344),
.Y(n_14448)
);

INVx2_ASAP7_75t_L g14449 ( 
.A(n_13572),
.Y(n_14449)
);

NAND2xp5_ASAP7_75t_L g14450 ( 
.A(n_13223),
.B(n_1344),
.Y(n_14450)
);

INVx2_ASAP7_75t_L g14451 ( 
.A(n_13812),
.Y(n_14451)
);

INVx2_ASAP7_75t_L g14452 ( 
.A(n_13259),
.Y(n_14452)
);

AND2x6_ASAP7_75t_L g14453 ( 
.A(n_13728),
.B(n_5872),
.Y(n_14453)
);

INVx1_ASAP7_75t_SL g14454 ( 
.A(n_12968),
.Y(n_14454)
);

INVx1_ASAP7_75t_L g14455 ( 
.A(n_13398),
.Y(n_14455)
);

AOI22xp5_ASAP7_75t_L g14456 ( 
.A1(n_13746),
.A2(n_1347),
.B1(n_1345),
.B2(n_1346),
.Y(n_14456)
);

HB1xp67_ASAP7_75t_L g14457 ( 
.A(n_12947),
.Y(n_14457)
);

OAI21xp5_ASAP7_75t_L g14458 ( 
.A1(n_13065),
.A2(n_1345),
.B(n_1347),
.Y(n_14458)
);

INVx1_ASAP7_75t_L g14459 ( 
.A(n_13590),
.Y(n_14459)
);

AOI22xp5_ASAP7_75t_L g14460 ( 
.A1(n_13832),
.A2(n_1350),
.B1(n_1348),
.B2(n_1349),
.Y(n_14460)
);

AND2x2_ASAP7_75t_SL g14461 ( 
.A(n_13227),
.B(n_1348),
.Y(n_14461)
);

INVx4_ASAP7_75t_L g14462 ( 
.A(n_12911),
.Y(n_14462)
);

CKINVDCx5p33_ASAP7_75t_R g14463 ( 
.A(n_13014),
.Y(n_14463)
);

OAI21xp5_ASAP7_75t_L g14464 ( 
.A1(n_13147),
.A2(n_1349),
.B(n_1350),
.Y(n_14464)
);

INVx1_ASAP7_75t_L g14465 ( 
.A(n_13159),
.Y(n_14465)
);

AND2x2_ASAP7_75t_L g14466 ( 
.A(n_13359),
.B(n_1351),
.Y(n_14466)
);

INVx2_ASAP7_75t_L g14467 ( 
.A(n_13215),
.Y(n_14467)
);

AOI22xp5_ASAP7_75t_L g14468 ( 
.A1(n_13873),
.A2(n_1354),
.B1(n_1351),
.B2(n_1352),
.Y(n_14468)
);

AND3x1_ASAP7_75t_SL g14469 ( 
.A(n_13228),
.B(n_13563),
.C(n_12921),
.Y(n_14469)
);

INVx2_ASAP7_75t_L g14470 ( 
.A(n_12917),
.Y(n_14470)
);

BUFx6f_ASAP7_75t_L g14471 ( 
.A(n_13179),
.Y(n_14471)
);

INVx2_ASAP7_75t_L g14472 ( 
.A(n_13508),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_13159),
.Y(n_14473)
);

BUFx12f_ASAP7_75t_L g14474 ( 
.A(n_13424),
.Y(n_14474)
);

NOR2xp33_ASAP7_75t_L g14475 ( 
.A(n_13252),
.B(n_1352),
.Y(n_14475)
);

AND2x4_ASAP7_75t_SL g14476 ( 
.A(n_12865),
.B(n_5873),
.Y(n_14476)
);

NAND2x1p5_ASAP7_75t_L g14477 ( 
.A(n_13876),
.B(n_5874),
.Y(n_14477)
);

NAND2xp5_ASAP7_75t_L g14478 ( 
.A(n_13235),
.B(n_1354),
.Y(n_14478)
);

INVx1_ASAP7_75t_L g14479 ( 
.A(n_13103),
.Y(n_14479)
);

NAND2xp5_ASAP7_75t_L g14480 ( 
.A(n_13236),
.B(n_1355),
.Y(n_14480)
);

INVx2_ASAP7_75t_L g14481 ( 
.A(n_13514),
.Y(n_14481)
);

NAND2x1p5_ASAP7_75t_L g14482 ( 
.A(n_13663),
.B(n_5875),
.Y(n_14482)
);

AND2x2_ASAP7_75t_L g14483 ( 
.A(n_13473),
.B(n_1355),
.Y(n_14483)
);

NAND2xp5_ASAP7_75t_L g14484 ( 
.A(n_13240),
.B(n_1356),
.Y(n_14484)
);

INVx1_ASAP7_75t_L g14485 ( 
.A(n_13103),
.Y(n_14485)
);

INVx2_ASAP7_75t_L g14486 ( 
.A(n_13528),
.Y(n_14486)
);

INVx1_ASAP7_75t_L g14487 ( 
.A(n_13808),
.Y(n_14487)
);

AOI22x1_ASAP7_75t_L g14488 ( 
.A1(n_13652),
.A2(n_1358),
.B1(n_1356),
.B2(n_1357),
.Y(n_14488)
);

NAND2xp5_ASAP7_75t_L g14489 ( 
.A(n_13254),
.B(n_1357),
.Y(n_14489)
);

BUFx6f_ASAP7_75t_L g14490 ( 
.A(n_13440),
.Y(n_14490)
);

NAND2xp5_ASAP7_75t_SL g14491 ( 
.A(n_13692),
.B(n_5876),
.Y(n_14491)
);

A2O1A1Ixp33_ASAP7_75t_L g14492 ( 
.A1(n_13814),
.A2(n_1360),
.B(n_1358),
.C(n_1359),
.Y(n_14492)
);

CKINVDCx5p33_ASAP7_75t_R g14493 ( 
.A(n_12825),
.Y(n_14493)
);

AND2x2_ASAP7_75t_L g14494 ( 
.A(n_13049),
.B(n_1359),
.Y(n_14494)
);

INVx1_ASAP7_75t_L g14495 ( 
.A(n_13808),
.Y(n_14495)
);

CKINVDCx5p33_ASAP7_75t_R g14496 ( 
.A(n_12997),
.Y(n_14496)
);

AND2x2_ASAP7_75t_L g14497 ( 
.A(n_13371),
.B(n_1360),
.Y(n_14497)
);

CKINVDCx5p33_ASAP7_75t_R g14498 ( 
.A(n_13479),
.Y(n_14498)
);

NAND2x1p5_ASAP7_75t_L g14499 ( 
.A(n_13666),
.B(n_5878),
.Y(n_14499)
);

INVx2_ASAP7_75t_L g14500 ( 
.A(n_13536),
.Y(n_14500)
);

INVx2_ASAP7_75t_L g14501 ( 
.A(n_13542),
.Y(n_14501)
);

AND2x2_ASAP7_75t_L g14502 ( 
.A(n_13527),
.B(n_1361),
.Y(n_14502)
);

INVx1_ASAP7_75t_L g14503 ( 
.A(n_13251),
.Y(n_14503)
);

NAND2xp5_ASAP7_75t_L g14504 ( 
.A(n_13276),
.B(n_1361),
.Y(n_14504)
);

AND2x2_ASAP7_75t_L g14505 ( 
.A(n_13291),
.B(n_1362),
.Y(n_14505)
);

NAND2xp5_ASAP7_75t_SL g14506 ( 
.A(n_13702),
.B(n_5879),
.Y(n_14506)
);

NAND2xp5_ASAP7_75t_L g14507 ( 
.A(n_13282),
.B(n_1363),
.Y(n_14507)
);

INVx1_ASAP7_75t_L g14508 ( 
.A(n_13251),
.Y(n_14508)
);

INVx2_ASAP7_75t_L g14509 ( 
.A(n_13546),
.Y(n_14509)
);

NAND2xp5_ASAP7_75t_L g14510 ( 
.A(n_13287),
.B(n_1363),
.Y(n_14510)
);

OAI22xp5_ASAP7_75t_SL g14511 ( 
.A1(n_13412),
.A2(n_1367),
.B1(n_1365),
.B2(n_1366),
.Y(n_14511)
);

NAND2xp5_ASAP7_75t_L g14512 ( 
.A(n_13289),
.B(n_1365),
.Y(n_14512)
);

INVx1_ASAP7_75t_L g14513 ( 
.A(n_13549),
.Y(n_14513)
);

INVx2_ASAP7_75t_L g14514 ( 
.A(n_13559),
.Y(n_14514)
);

AND2x4_ASAP7_75t_L g14515 ( 
.A(n_13055),
.B(n_5880),
.Y(n_14515)
);

BUFx6f_ASAP7_75t_L g14516 ( 
.A(n_13205),
.Y(n_14516)
);

OAI21xp5_ASAP7_75t_L g14517 ( 
.A1(n_13483),
.A2(n_1366),
.B(n_1367),
.Y(n_14517)
);

NAND2xp5_ASAP7_75t_L g14518 ( 
.A(n_13296),
.B(n_1368),
.Y(n_14518)
);

INVx2_ASAP7_75t_L g14519 ( 
.A(n_13560),
.Y(n_14519)
);

AND2x2_ASAP7_75t_L g14520 ( 
.A(n_13316),
.B(n_1368),
.Y(n_14520)
);

BUFx3_ASAP7_75t_L g14521 ( 
.A(n_13214),
.Y(n_14521)
);

INVx1_ASAP7_75t_L g14522 ( 
.A(n_13591),
.Y(n_14522)
);

INVx3_ASAP7_75t_SL g14523 ( 
.A(n_13423),
.Y(n_14523)
);

BUFx4f_ASAP7_75t_L g14524 ( 
.A(n_13849),
.Y(n_14524)
);

NAND2xp5_ASAP7_75t_L g14525 ( 
.A(n_13322),
.B(n_1369),
.Y(n_14525)
);

AND2x2_ASAP7_75t_L g14526 ( 
.A(n_12888),
.B(n_1370),
.Y(n_14526)
);

NAND2xp5_ASAP7_75t_SL g14527 ( 
.A(n_13834),
.B(n_5881),
.Y(n_14527)
);

NOR2xp33_ASAP7_75t_R g14528 ( 
.A(n_13292),
.B(n_1371),
.Y(n_14528)
);

OR2x2_ASAP7_75t_L g14529 ( 
.A(n_13325),
.B(n_13332),
.Y(n_14529)
);

NAND2xp5_ASAP7_75t_L g14530 ( 
.A(n_13352),
.B(n_1371),
.Y(n_14530)
);

NAND2xp5_ASAP7_75t_L g14531 ( 
.A(n_13366),
.B(n_1372),
.Y(n_14531)
);

AND2x2_ASAP7_75t_L g14532 ( 
.A(n_12942),
.B(n_1372),
.Y(n_14532)
);

INVx1_ASAP7_75t_L g14533 ( 
.A(n_13596),
.Y(n_14533)
);

INVx3_ASAP7_75t_L g14534 ( 
.A(n_13500),
.Y(n_14534)
);

INVx2_ASAP7_75t_L g14535 ( 
.A(n_12992),
.Y(n_14535)
);

NAND2xp5_ASAP7_75t_L g14536 ( 
.A(n_13367),
.B(n_1373),
.Y(n_14536)
);

AOI22xp5_ASAP7_75t_L g14537 ( 
.A1(n_13883),
.A2(n_1376),
.B1(n_1374),
.B2(n_1375),
.Y(n_14537)
);

A2O1A1Ixp33_ASAP7_75t_SL g14538 ( 
.A1(n_13437),
.A2(n_1376),
.B(n_1374),
.C(n_1375),
.Y(n_14538)
);

AOI22xp33_ASAP7_75t_L g14539 ( 
.A1(n_13021),
.A2(n_13284),
.B1(n_13318),
.B2(n_13034),
.Y(n_14539)
);

INVx4_ASAP7_75t_L g14540 ( 
.A(n_12865),
.Y(n_14540)
);

CKINVDCx20_ASAP7_75t_R g14541 ( 
.A(n_13317),
.Y(n_14541)
);

AND2x4_ASAP7_75t_L g14542 ( 
.A(n_13517),
.B(n_5883),
.Y(n_14542)
);

BUFx2_ASAP7_75t_L g14543 ( 
.A(n_12869),
.Y(n_14543)
);

INVx2_ASAP7_75t_L g14544 ( 
.A(n_13059),
.Y(n_14544)
);

INVx1_ASAP7_75t_L g14545 ( 
.A(n_13636),
.Y(n_14545)
);

NAND2xp5_ASAP7_75t_L g14546 ( 
.A(n_13382),
.B(n_1377),
.Y(n_14546)
);

NAND2xp5_ASAP7_75t_L g14547 ( 
.A(n_13387),
.B(n_1377),
.Y(n_14547)
);

NAND2x1_ASAP7_75t_L g14548 ( 
.A(n_13034),
.B(n_1378),
.Y(n_14548)
);

AND2x2_ASAP7_75t_L g14549 ( 
.A(n_12960),
.B(n_1378),
.Y(n_14549)
);

NAND2xp5_ASAP7_75t_SL g14550 ( 
.A(n_13452),
.B(n_5884),
.Y(n_14550)
);

BUFx3_ASAP7_75t_L g14551 ( 
.A(n_13302),
.Y(n_14551)
);

AOI22xp33_ASAP7_75t_L g14552 ( 
.A1(n_13001),
.A2(n_13384),
.B1(n_13187),
.B2(n_13176),
.Y(n_14552)
);

OR2x2_ASAP7_75t_L g14553 ( 
.A(n_13389),
.B(n_1379),
.Y(n_14553)
);

NAND3xp33_ASAP7_75t_SL g14554 ( 
.A(n_13833),
.B(n_1379),
.C(n_1380),
.Y(n_14554)
);

AND2x4_ASAP7_75t_L g14555 ( 
.A(n_13517),
.B(n_5885),
.Y(n_14555)
);

INVxp67_ASAP7_75t_L g14556 ( 
.A(n_13400),
.Y(n_14556)
);

CKINVDCx5p33_ASAP7_75t_R g14557 ( 
.A(n_13101),
.Y(n_14557)
);

INVx1_ASAP7_75t_L g14558 ( 
.A(n_13848),
.Y(n_14558)
);

CKINVDCx5p33_ASAP7_75t_R g14559 ( 
.A(n_13116),
.Y(n_14559)
);

CKINVDCx20_ASAP7_75t_R g14560 ( 
.A(n_13586),
.Y(n_14560)
);

BUFx6f_ASAP7_75t_L g14561 ( 
.A(n_13881),
.Y(n_14561)
);

NOR2xp67_ASAP7_75t_L g14562 ( 
.A(n_13402),
.B(n_1380),
.Y(n_14562)
);

INVx1_ASAP7_75t_L g14563 ( 
.A(n_12843),
.Y(n_14563)
);

INVx2_ASAP7_75t_L g14564 ( 
.A(n_13406),
.Y(n_14564)
);

OAI22xp5_ASAP7_75t_SL g14565 ( 
.A1(n_13100),
.A2(n_1383),
.B1(n_1381),
.B2(n_1382),
.Y(n_14565)
);

CKINVDCx20_ASAP7_75t_R g14566 ( 
.A(n_13355),
.Y(n_14566)
);

NAND2xp5_ASAP7_75t_L g14567 ( 
.A(n_13403),
.B(n_1382),
.Y(n_14567)
);

NAND2xp5_ASAP7_75t_L g14568 ( 
.A(n_13407),
.B(n_13415),
.Y(n_14568)
);

AND2x2_ASAP7_75t_L g14569 ( 
.A(n_13537),
.B(n_1383),
.Y(n_14569)
);

A2O1A1Ixp33_ASAP7_75t_SL g14570 ( 
.A1(n_12918),
.A2(n_1386),
.B(n_1384),
.C(n_1385),
.Y(n_14570)
);

INVx1_ASAP7_75t_L g14571 ( 
.A(n_12908),
.Y(n_14571)
);

AOI22xp5_ASAP7_75t_L g14572 ( 
.A1(n_13885),
.A2(n_13257),
.B1(n_12891),
.B2(n_12919),
.Y(n_14572)
);

AND3x1_ASAP7_75t_SL g14573 ( 
.A(n_12932),
.B(n_1384),
.C(n_1385),
.Y(n_14573)
);

CKINVDCx11_ASAP7_75t_R g14574 ( 
.A(n_12794),
.Y(n_14574)
);

INVx1_ASAP7_75t_L g14575 ( 
.A(n_13183),
.Y(n_14575)
);

AND2x2_ASAP7_75t_L g14576 ( 
.A(n_13441),
.B(n_1387),
.Y(n_14576)
);

NAND2xp5_ASAP7_75t_L g14577 ( 
.A(n_13433),
.B(n_1387),
.Y(n_14577)
);

NAND2xp5_ASAP7_75t_L g14578 ( 
.A(n_13446),
.B(n_1388),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_13449),
.Y(n_14579)
);

INVx1_ASAP7_75t_L g14580 ( 
.A(n_13451),
.Y(n_14580)
);

NAND2xp5_ASAP7_75t_L g14581 ( 
.A(n_13466),
.B(n_13489),
.Y(n_14581)
);

INVx1_ASAP7_75t_L g14582 ( 
.A(n_13496),
.Y(n_14582)
);

CKINVDCx5p33_ASAP7_75t_R g14583 ( 
.A(n_13211),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_13443),
.B(n_13453),
.Y(n_14584)
);

AOI22xp33_ASAP7_75t_SL g14585 ( 
.A1(n_13602),
.A2(n_1390),
.B1(n_1388),
.B2(n_1389),
.Y(n_14585)
);

NAND2xp5_ASAP7_75t_SL g14586 ( 
.A(n_12944),
.B(n_5886),
.Y(n_14586)
);

AND2x2_ASAP7_75t_L g14587 ( 
.A(n_13476),
.B(n_1389),
.Y(n_14587)
);

NOR2xp33_ASAP7_75t_L g14588 ( 
.A(n_13341),
.B(n_1390),
.Y(n_14588)
);

AND2x4_ASAP7_75t_L g14589 ( 
.A(n_13113),
.B(n_5887),
.Y(n_14589)
);

NAND2xp5_ASAP7_75t_SL g14590 ( 
.A(n_13023),
.B(n_5888),
.Y(n_14590)
);

INVx1_ASAP7_75t_L g14591 ( 
.A(n_13497),
.Y(n_14591)
);

INVx1_ASAP7_75t_L g14592 ( 
.A(n_13498),
.Y(n_14592)
);

INVx2_ASAP7_75t_L g14593 ( 
.A(n_12939),
.Y(n_14593)
);

INVx1_ASAP7_75t_L g14594 ( 
.A(n_13501),
.Y(n_14594)
);

NAND2xp5_ASAP7_75t_L g14595 ( 
.A(n_13253),
.B(n_1391),
.Y(n_14595)
);

INVxp67_ASAP7_75t_L g14596 ( 
.A(n_13217),
.Y(n_14596)
);

NAND2xp5_ASAP7_75t_SL g14597 ( 
.A(n_13610),
.B(n_13612),
.Y(n_14597)
);

CKINVDCx5p33_ASAP7_75t_R g14598 ( 
.A(n_13070),
.Y(n_14598)
);

NAND2xp5_ASAP7_75t_L g14599 ( 
.A(n_13280),
.B(n_1392),
.Y(n_14599)
);

NAND2xp5_ASAP7_75t_SL g14600 ( 
.A(n_13748),
.B(n_5889),
.Y(n_14600)
);

AOI22xp5_ASAP7_75t_L g14601 ( 
.A1(n_12899),
.A2(n_1394),
.B1(n_1392),
.B2(n_1393),
.Y(n_14601)
);

CKINVDCx5p33_ASAP7_75t_R g14602 ( 
.A(n_13491),
.Y(n_14602)
);

NAND2xp5_ASAP7_75t_SL g14603 ( 
.A(n_13799),
.B(n_13870),
.Y(n_14603)
);

HB1xp67_ASAP7_75t_L g14604 ( 
.A(n_12994),
.Y(n_14604)
);

AND2x2_ASAP7_75t_L g14605 ( 
.A(n_13513),
.B(n_1393),
.Y(n_14605)
);

AOI22xp5_ASAP7_75t_L g14606 ( 
.A1(n_13029),
.A2(n_1397),
.B1(n_1394),
.B2(n_1396),
.Y(n_14606)
);

NAND2xp5_ASAP7_75t_L g14607 ( 
.A(n_13288),
.B(n_13334),
.Y(n_14607)
);

INVx1_ASAP7_75t_L g14608 ( 
.A(n_13265),
.Y(n_14608)
);

INVx1_ASAP7_75t_L g14609 ( 
.A(n_13592),
.Y(n_14609)
);

AND3x1_ASAP7_75t_SL g14610 ( 
.A(n_13164),
.B(n_1396),
.C(n_1397),
.Y(n_14610)
);

NAND2xp5_ASAP7_75t_L g14611 ( 
.A(n_13566),
.B(n_1398),
.Y(n_14611)
);

BUFx3_ASAP7_75t_L g14612 ( 
.A(n_13529),
.Y(n_14612)
);

AND3x1_ASAP7_75t_SL g14613 ( 
.A(n_13309),
.B(n_1398),
.C(n_1399),
.Y(n_14613)
);

INVx2_ASAP7_75t_L g14614 ( 
.A(n_13619),
.Y(n_14614)
);

AND2x2_ASAP7_75t_L g14615 ( 
.A(n_13541),
.B(n_1399),
.Y(n_14615)
);

INVx2_ASAP7_75t_L g14616 ( 
.A(n_13798),
.Y(n_14616)
);

AND2x2_ASAP7_75t_L g14617 ( 
.A(n_13544),
.B(n_13562),
.Y(n_14617)
);

INVx2_ASAP7_75t_L g14618 ( 
.A(n_13608),
.Y(n_14618)
);

INVx1_ASAP7_75t_L g14619 ( 
.A(n_13522),
.Y(n_14619)
);

NAND2xp5_ASAP7_75t_L g14620 ( 
.A(n_13168),
.B(n_1400),
.Y(n_14620)
);

AOI22xp5_ASAP7_75t_L g14621 ( 
.A1(n_13156),
.A2(n_1402),
.B1(n_1400),
.B2(n_1401),
.Y(n_14621)
);

BUFx8_ASAP7_75t_L g14622 ( 
.A(n_13372),
.Y(n_14622)
);

NAND2xp5_ASAP7_75t_L g14623 ( 
.A(n_12961),
.B(n_1401),
.Y(n_14623)
);

AND2x2_ASAP7_75t_L g14624 ( 
.A(n_13117),
.B(n_1402),
.Y(n_14624)
);

INVx2_ASAP7_75t_L g14625 ( 
.A(n_13713),
.Y(n_14625)
);

BUFx12f_ASAP7_75t_L g14626 ( 
.A(n_13378),
.Y(n_14626)
);

INVx2_ASAP7_75t_L g14627 ( 
.A(n_12951),
.Y(n_14627)
);

AND2x2_ASAP7_75t_L g14628 ( 
.A(n_13524),
.B(n_1403),
.Y(n_14628)
);

AND2x2_ASAP7_75t_L g14629 ( 
.A(n_12959),
.B(n_1403),
.Y(n_14629)
);

INVx2_ASAP7_75t_L g14630 ( 
.A(n_12963),
.Y(n_14630)
);

AOI22xp5_ASAP7_75t_L g14631 ( 
.A1(n_13218),
.A2(n_1406),
.B1(n_1404),
.B2(n_1405),
.Y(n_14631)
);

NAND2xp5_ASAP7_75t_L g14632 ( 
.A(n_12931),
.B(n_1405),
.Y(n_14632)
);

CKINVDCx5p33_ASAP7_75t_R g14633 ( 
.A(n_13576),
.Y(n_14633)
);

NAND2xp5_ASAP7_75t_L g14634 ( 
.A(n_13102),
.B(n_1406),
.Y(n_14634)
);

AND2x2_ASAP7_75t_L g14635 ( 
.A(n_12965),
.B(n_1407),
.Y(n_14635)
);

BUFx2_ASAP7_75t_L g14636 ( 
.A(n_12837),
.Y(n_14636)
);

NAND2xp5_ASAP7_75t_L g14637 ( 
.A(n_13463),
.B(n_1407),
.Y(n_14637)
);

AND2x2_ASAP7_75t_L g14638 ( 
.A(n_13444),
.B(n_1408),
.Y(n_14638)
);

INVxp67_ASAP7_75t_L g14639 ( 
.A(n_12824),
.Y(n_14639)
);

CKINVDCx5p33_ASAP7_75t_R g14640 ( 
.A(n_13603),
.Y(n_14640)
);

INVx2_ASAP7_75t_L g14641 ( 
.A(n_12957),
.Y(n_14641)
);

AND2x2_ASAP7_75t_L g14642 ( 
.A(n_13201),
.B(n_13221),
.Y(n_14642)
);

NOR2xp33_ASAP7_75t_R g14643 ( 
.A(n_13594),
.B(n_1408),
.Y(n_14643)
);

AND3x1_ASAP7_75t_SL g14644 ( 
.A(n_13641),
.B(n_1409),
.C(n_1410),
.Y(n_14644)
);

NAND2xp5_ASAP7_75t_L g14645 ( 
.A(n_13464),
.B(n_1409),
.Y(n_14645)
);

INVx2_ASAP7_75t_L g14646 ( 
.A(n_12972),
.Y(n_14646)
);

INVx2_ASAP7_75t_L g14647 ( 
.A(n_13037),
.Y(n_14647)
);

AND2x2_ASAP7_75t_L g14648 ( 
.A(n_13222),
.B(n_1410),
.Y(n_14648)
);

OAI22xp5_ASAP7_75t_SL g14649 ( 
.A1(n_12809),
.A2(n_1413),
.B1(n_1411),
.B2(n_1412),
.Y(n_14649)
);

AO22x1_ASAP7_75t_L g14650 ( 
.A1(n_13558),
.A2(n_1413),
.B1(n_1411),
.B2(n_1412),
.Y(n_14650)
);

BUFx4f_ASAP7_75t_L g14651 ( 
.A(n_13580),
.Y(n_14651)
);

INVx3_ASAP7_75t_L g14652 ( 
.A(n_13107),
.Y(n_14652)
);

CKINVDCx5p33_ASAP7_75t_R g14653 ( 
.A(n_13645),
.Y(n_14653)
);

CKINVDCx6p67_ASAP7_75t_R g14654 ( 
.A(n_13561),
.Y(n_14654)
);

AOI22xp33_ASAP7_75t_L g14655 ( 
.A1(n_12975),
.A2(n_1416),
.B1(n_1414),
.B2(n_1415),
.Y(n_14655)
);

INVx1_ASAP7_75t_L g14656 ( 
.A(n_13569),
.Y(n_14656)
);

NAND2x1p5_ASAP7_75t_L g14657 ( 
.A(n_13739),
.B(n_5890),
.Y(n_14657)
);

INVxp67_ASAP7_75t_SL g14658 ( 
.A(n_13492),
.Y(n_14658)
);

CKINVDCx20_ASAP7_75t_R g14659 ( 
.A(n_13120),
.Y(n_14659)
);

BUFx6f_ASAP7_75t_L g14660 ( 
.A(n_13057),
.Y(n_14660)
);

BUFx3_ASAP7_75t_L g14661 ( 
.A(n_13533),
.Y(n_14661)
);

AOI22xp5_ASAP7_75t_L g14662 ( 
.A1(n_13312),
.A2(n_1416),
.B1(n_1414),
.B2(n_1415),
.Y(n_14662)
);

NAND2xp5_ASAP7_75t_L g14663 ( 
.A(n_13465),
.B(n_1417),
.Y(n_14663)
);

AND3x1_ASAP7_75t_SL g14664 ( 
.A(n_13690),
.B(n_1418),
.C(n_1419),
.Y(n_14664)
);

NAND2xp5_ASAP7_75t_L g14665 ( 
.A(n_13502),
.B(n_13535),
.Y(n_14665)
);

CKINVDCx5p33_ASAP7_75t_R g14666 ( 
.A(n_13711),
.Y(n_14666)
);

CKINVDCx5p33_ASAP7_75t_R g14667 ( 
.A(n_13751),
.Y(n_14667)
);

AND2x2_ASAP7_75t_L g14668 ( 
.A(n_12874),
.B(n_1419),
.Y(n_14668)
);

INVx1_ASAP7_75t_L g14669 ( 
.A(n_13181),
.Y(n_14669)
);

NOR2xp67_ASAP7_75t_L g14670 ( 
.A(n_12801),
.B(n_1420),
.Y(n_14670)
);

NOR2xp33_ASAP7_75t_L g14671 ( 
.A(n_13460),
.B(n_1420),
.Y(n_14671)
);

INVx3_ASAP7_75t_L g14672 ( 
.A(n_13093),
.Y(n_14672)
);

INVx1_ASAP7_75t_L g14673 ( 
.A(n_13350),
.Y(n_14673)
);

NAND2xp5_ASAP7_75t_L g14674 ( 
.A(n_13540),
.B(n_1421),
.Y(n_14674)
);

BUFx4f_ASAP7_75t_L g14675 ( 
.A(n_13363),
.Y(n_14675)
);

INVx8_ASAP7_75t_L g14676 ( 
.A(n_12796),
.Y(n_14676)
);

BUFx2_ASAP7_75t_L g14677 ( 
.A(n_13405),
.Y(n_14677)
);

NAND2xp5_ASAP7_75t_L g14678 ( 
.A(n_13413),
.B(n_1421),
.Y(n_14678)
);

INVx2_ASAP7_75t_L g14679 ( 
.A(n_12840),
.Y(n_14679)
);

NOR2xp33_ASAP7_75t_L g14680 ( 
.A(n_13461),
.B(n_1423),
.Y(n_14680)
);

INVx4_ASAP7_75t_L g14681 ( 
.A(n_12798),
.Y(n_14681)
);

INVx1_ASAP7_75t_L g14682 ( 
.A(n_13521),
.Y(n_14682)
);

CKINVDCx5p33_ASAP7_75t_R g14683 ( 
.A(n_13771),
.Y(n_14683)
);

INVxp33_ASAP7_75t_L g14684 ( 
.A(n_13022),
.Y(n_14684)
);

INVx2_ASAP7_75t_L g14685 ( 
.A(n_13503),
.Y(n_14685)
);

NAND2xp5_ASAP7_75t_SL g14686 ( 
.A(n_13249),
.B(n_5893),
.Y(n_14686)
);

INVx2_ASAP7_75t_L g14687 ( 
.A(n_13506),
.Y(n_14687)
);

AND2x2_ASAP7_75t_L g14688 ( 
.A(n_13006),
.B(n_1423),
.Y(n_14688)
);

NAND2xp5_ASAP7_75t_L g14689 ( 
.A(n_13457),
.B(n_1424),
.Y(n_14689)
);

NOR2xp33_ASAP7_75t_L g14690 ( 
.A(n_13025),
.B(n_1424),
.Y(n_14690)
);

NAND2xp5_ASAP7_75t_L g14691 ( 
.A(n_12882),
.B(n_1425),
.Y(n_14691)
);

INVx2_ASAP7_75t_L g14692 ( 
.A(n_13305),
.Y(n_14692)
);

NAND2xp5_ASAP7_75t_L g14693 ( 
.A(n_13411),
.B(n_1425),
.Y(n_14693)
);

AND2x2_ASAP7_75t_L g14694 ( 
.A(n_13015),
.B(n_1426),
.Y(n_14694)
);

INVx2_ASAP7_75t_L g14695 ( 
.A(n_13471),
.Y(n_14695)
);

BUFx3_ASAP7_75t_L g14696 ( 
.A(n_13545),
.Y(n_14696)
);

CKINVDCx20_ASAP7_75t_R g14697 ( 
.A(n_13283),
.Y(n_14697)
);

NAND2xp5_ASAP7_75t_L g14698 ( 
.A(n_13169),
.B(n_1426),
.Y(n_14698)
);

AND2x2_ASAP7_75t_L g14699 ( 
.A(n_13368),
.B(n_1427),
.Y(n_14699)
);

NAND2xp5_ASAP7_75t_SL g14700 ( 
.A(n_13315),
.B(n_5894),
.Y(n_14700)
);

AOI221x1_ASAP7_75t_L g14701 ( 
.A1(n_12806),
.A2(n_1429),
.B1(n_1427),
.B2(n_1428),
.C(n_1430),
.Y(n_14701)
);

INVx3_ASAP7_75t_L g14702 ( 
.A(n_13582),
.Y(n_14702)
);

INVx2_ASAP7_75t_L g14703 ( 
.A(n_13481),
.Y(n_14703)
);

INVx2_ASAP7_75t_L g14704 ( 
.A(n_13241),
.Y(n_14704)
);

OAI21xp5_ASAP7_75t_L g14705 ( 
.A1(n_13343),
.A2(n_1428),
.B(n_1429),
.Y(n_14705)
);

AOI22xp33_ASAP7_75t_L g14706 ( 
.A1(n_13161),
.A2(n_1432),
.B1(n_1430),
.B2(n_1431),
.Y(n_14706)
);

NAND2xp5_ASAP7_75t_L g14707 ( 
.A(n_13207),
.B(n_1431),
.Y(n_14707)
);

NAND2xp5_ASAP7_75t_L g14708 ( 
.A(n_13163),
.B(n_1432),
.Y(n_14708)
);

INVxp67_ASAP7_75t_L g14709 ( 
.A(n_13553),
.Y(n_14709)
);

NAND2xp5_ASAP7_75t_L g14710 ( 
.A(n_12925),
.B(n_1433),
.Y(n_14710)
);

NAND2xp5_ASAP7_75t_L g14711 ( 
.A(n_13459),
.B(n_1434),
.Y(n_14711)
);

OR2x2_ASAP7_75t_L g14712 ( 
.A(n_13258),
.B(n_13277),
.Y(n_14712)
);

HB1xp67_ASAP7_75t_L g14713 ( 
.A(n_13373),
.Y(n_14713)
);

INVx1_ASAP7_75t_L g14714 ( 
.A(n_13204),
.Y(n_14714)
);

AOI22xp5_ASAP7_75t_L g14715 ( 
.A1(n_13056),
.A2(n_1436),
.B1(n_1434),
.B2(n_1435),
.Y(n_14715)
);

INVx5_ASAP7_75t_L g14716 ( 
.A(n_13226),
.Y(n_14716)
);

INVx1_ASAP7_75t_L g14717 ( 
.A(n_13381),
.Y(n_14717)
);

AOI22xp5_ASAP7_75t_L g14718 ( 
.A1(n_13072),
.A2(n_1438),
.B1(n_1435),
.B2(n_1437),
.Y(n_14718)
);

AND2x2_ASAP7_75t_L g14719 ( 
.A(n_13428),
.B(n_1437),
.Y(n_14719)
);

NAND2xp5_ASAP7_75t_SL g14720 ( 
.A(n_13482),
.B(n_5895),
.Y(n_14720)
);

NAND2xp5_ASAP7_75t_L g14721 ( 
.A(n_13653),
.B(n_13704),
.Y(n_14721)
);

BUFx3_ASAP7_75t_L g14722 ( 
.A(n_13550),
.Y(n_14722)
);

INVx2_ASAP7_75t_L g14723 ( 
.A(n_13769),
.Y(n_14723)
);

NAND2xp5_ASAP7_75t_L g14724 ( 
.A(n_13723),
.B(n_1438),
.Y(n_14724)
);

NAND2xp5_ASAP7_75t_L g14725 ( 
.A(n_13768),
.B(n_1439),
.Y(n_14725)
);

INVx1_ASAP7_75t_L g14726 ( 
.A(n_13409),
.Y(n_14726)
);

NAND2xp5_ASAP7_75t_L g14727 ( 
.A(n_13796),
.B(n_1439),
.Y(n_14727)
);

NAND2xp5_ASAP7_75t_L g14728 ( 
.A(n_13822),
.B(n_1440),
.Y(n_14728)
);

A2O1A1Ixp33_ASAP7_75t_L g14729 ( 
.A1(n_12980),
.A2(n_1442),
.B(n_1440),
.C(n_1441),
.Y(n_14729)
);

INVx2_ASAP7_75t_L g14730 ( 
.A(n_13775),
.Y(n_14730)
);

INVx2_ASAP7_75t_L g14731 ( 
.A(n_13777),
.Y(n_14731)
);

AND3x1_ASAP7_75t_SL g14732 ( 
.A(n_13772),
.B(n_1441),
.C(n_1443),
.Y(n_14732)
);

INVx2_ASAP7_75t_L g14733 ( 
.A(n_13794),
.Y(n_14733)
);

BUFx6f_ASAP7_75t_L g14734 ( 
.A(n_13803),
.Y(n_14734)
);

NAND2xp5_ASAP7_75t_SL g14735 ( 
.A(n_13782),
.B(n_5896),
.Y(n_14735)
);

OAI22xp5_ASAP7_75t_L g14736 ( 
.A1(n_13601),
.A2(n_1445),
.B1(n_1443),
.B2(n_1444),
.Y(n_14736)
);

INVx1_ASAP7_75t_L g14737 ( 
.A(n_13462),
.Y(n_14737)
);

BUFx3_ASAP7_75t_L g14738 ( 
.A(n_13783),
.Y(n_14738)
);

NAND2xp5_ASAP7_75t_L g14739 ( 
.A(n_13852),
.B(n_13863),
.Y(n_14739)
);

INVxp67_ASAP7_75t_L g14740 ( 
.A(n_13824),
.Y(n_14740)
);

CKINVDCx11_ASAP7_75t_R g14741 ( 
.A(n_13797),
.Y(n_14741)
);

NAND2xp5_ASAP7_75t_L g14742 ( 
.A(n_13896),
.B(n_1444),
.Y(n_14742)
);

INVx2_ASAP7_75t_L g14743 ( 
.A(n_13826),
.Y(n_14743)
);

NAND2xp5_ASAP7_75t_L g14744 ( 
.A(n_12998),
.B(n_1446),
.Y(n_14744)
);

INVx1_ASAP7_75t_L g14745 ( 
.A(n_13574),
.Y(n_14745)
);

AND2x2_ASAP7_75t_L g14746 ( 
.A(n_13447),
.B(n_1447),
.Y(n_14746)
);

OAI21xp5_ASAP7_75t_L g14747 ( 
.A1(n_12879),
.A2(n_1447),
.B(n_1448),
.Y(n_14747)
);

AOI22xp5_ASAP7_75t_L g14748 ( 
.A1(n_13328),
.A2(n_1451),
.B1(n_1449),
.B2(n_1450),
.Y(n_14748)
);

INVx2_ASAP7_75t_SL g14749 ( 
.A(n_13828),
.Y(n_14749)
);

INVx3_ASAP7_75t_L g14750 ( 
.A(n_13846),
.Y(n_14750)
);

AND2x2_ASAP7_75t_L g14751 ( 
.A(n_13860),
.B(n_1449),
.Y(n_14751)
);

INVx1_ASAP7_75t_L g14752 ( 
.A(n_13551),
.Y(n_14752)
);

NAND2xp5_ASAP7_75t_L g14753 ( 
.A(n_13082),
.B(n_1450),
.Y(n_14753)
);

NAND2xp5_ASAP7_75t_SL g14754 ( 
.A(n_13847),
.B(n_5897),
.Y(n_14754)
);

NAND2xp5_ASAP7_75t_L g14755 ( 
.A(n_13633),
.B(n_1451),
.Y(n_14755)
);

OAI22xp5_ASAP7_75t_SL g14756 ( 
.A1(n_13197),
.A2(n_1454),
.B1(n_1452),
.B2(n_1453),
.Y(n_14756)
);

BUFx8_ASAP7_75t_L g14757 ( 
.A(n_13888),
.Y(n_14757)
);

INVx2_ASAP7_75t_L g14758 ( 
.A(n_13882),
.Y(n_14758)
);

BUFx2_ASAP7_75t_L g14759 ( 
.A(n_13286),
.Y(n_14759)
);

CKINVDCx5p33_ASAP7_75t_R g14760 ( 
.A(n_13897),
.Y(n_14760)
);

NAND2xp5_ASAP7_75t_L g14761 ( 
.A(n_13105),
.B(n_1452),
.Y(n_14761)
);

INVx1_ASAP7_75t_L g14762 ( 
.A(n_13348),
.Y(n_14762)
);

OR2x2_ASAP7_75t_L g14763 ( 
.A(n_13891),
.B(n_1453),
.Y(n_14763)
);

INVx1_ASAP7_75t_L g14764 ( 
.A(n_13361),
.Y(n_14764)
);

OAI22xp5_ASAP7_75t_L g14765 ( 
.A1(n_13669),
.A2(n_1457),
.B1(n_1455),
.B2(n_1456),
.Y(n_14765)
);

OAI22xp5_ASAP7_75t_L g14766 ( 
.A1(n_13703),
.A2(n_13875),
.B1(n_13892),
.B2(n_13838),
.Y(n_14766)
);

BUFx3_ASAP7_75t_L g14767 ( 
.A(n_13134),
.Y(n_14767)
);

INVx1_ASAP7_75t_L g14768 ( 
.A(n_13418),
.Y(n_14768)
);

NAND2xp5_ASAP7_75t_L g14769 ( 
.A(n_13429),
.B(n_1456),
.Y(n_14769)
);

INVx2_ASAP7_75t_L g14770 ( 
.A(n_13573),
.Y(n_14770)
);

CKINVDCx5p33_ASAP7_75t_R g14771 ( 
.A(n_13531),
.Y(n_14771)
);

INVxp33_ASAP7_75t_L g14772 ( 
.A(n_13584),
.Y(n_14772)
);

INVx2_ASAP7_75t_L g14773 ( 
.A(n_13583),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_13266),
.Y(n_14774)
);

CKINVDCx20_ASAP7_75t_R g14775 ( 
.A(n_13231),
.Y(n_14775)
);

NAND2xp5_ASAP7_75t_L g14776 ( 
.A(n_13516),
.B(n_1458),
.Y(n_14776)
);

NAND2xp5_ASAP7_75t_L g14777 ( 
.A(n_13196),
.B(n_1458),
.Y(n_14777)
);

BUFx6f_ASAP7_75t_L g14778 ( 
.A(n_13188),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_13548),
.Y(n_14779)
);

AND3x1_ASAP7_75t_SL g14780 ( 
.A(n_13518),
.B(n_1459),
.C(n_1460),
.Y(n_14780)
);

INVx2_ASAP7_75t_L g14781 ( 
.A(n_13375),
.Y(n_14781)
);

CKINVDCx14_ASAP7_75t_R g14782 ( 
.A(n_13138),
.Y(n_14782)
);

NAND2xp5_ASAP7_75t_L g14783 ( 
.A(n_13098),
.B(n_13261),
.Y(n_14783)
);

INVx1_ASAP7_75t_L g14784 ( 
.A(n_13229),
.Y(n_14784)
);

AND3x1_ASAP7_75t_SL g14785 ( 
.A(n_12803),
.B(n_1459),
.C(n_1460),
.Y(n_14785)
);

AOI22xp33_ASAP7_75t_L g14786 ( 
.A1(n_13180),
.A2(n_1463),
.B1(n_1461),
.B2(n_1462),
.Y(n_14786)
);

INVxp67_ASAP7_75t_L g14787 ( 
.A(n_13420),
.Y(n_14787)
);

INVx3_ASAP7_75t_L g14788 ( 
.A(n_13198),
.Y(n_14788)
);

AND2x2_ASAP7_75t_L g14789 ( 
.A(n_13585),
.B(n_1461),
.Y(n_14789)
);

HB1xp67_ASAP7_75t_L g14790 ( 
.A(n_13588),
.Y(n_14790)
);

INVx1_ASAP7_75t_L g14791 ( 
.A(n_12820),
.Y(n_14791)
);

INVx1_ASAP7_75t_L g14792 ( 
.A(n_12833),
.Y(n_14792)
);

NAND2xp5_ASAP7_75t_L g14793 ( 
.A(n_13306),
.B(n_1462),
.Y(n_14793)
);

CKINVDCx11_ASAP7_75t_R g14794 ( 
.A(n_13519),
.Y(n_14794)
);

OAI22xp5_ASAP7_75t_L g14795 ( 
.A1(n_13336),
.A2(n_1465),
.B1(n_1463),
.B2(n_1464),
.Y(n_14795)
);

BUFx6f_ASAP7_75t_L g14796 ( 
.A(n_13243),
.Y(n_14796)
);

INVx1_ASAP7_75t_L g14797 ( 
.A(n_12905),
.Y(n_14797)
);

AND2x2_ASAP7_75t_L g14798 ( 
.A(n_13598),
.B(n_1465),
.Y(n_14798)
);

INVx2_ASAP7_75t_L g14799 ( 
.A(n_13383),
.Y(n_14799)
);

AOI22xp33_ASAP7_75t_L g14800 ( 
.A1(n_13200),
.A2(n_13202),
.B1(n_13419),
.B2(n_13416),
.Y(n_14800)
);

NAND2xp5_ASAP7_75t_L g14801 ( 
.A(n_13342),
.B(n_1466),
.Y(n_14801)
);

OAI22xp5_ASAP7_75t_SL g14802 ( 
.A1(n_13385),
.A2(n_1468),
.B1(n_1466),
.B2(n_1467),
.Y(n_14802)
);

NAND2xp5_ASAP7_75t_L g14803 ( 
.A(n_13396),
.B(n_1468),
.Y(n_14803)
);

INVx1_ASAP7_75t_L g14804 ( 
.A(n_13051),
.Y(n_14804)
);

NOR2xp33_ASAP7_75t_L g14805 ( 
.A(n_13255),
.B(n_1469),
.Y(n_14805)
);

INVx2_ASAP7_75t_L g14806 ( 
.A(n_13414),
.Y(n_14806)
);

INVx4_ASAP7_75t_L g14807 ( 
.A(n_13185),
.Y(n_14807)
);

NOR2xp33_ASAP7_75t_L g14808 ( 
.A(n_13515),
.B(n_1469),
.Y(n_14808)
);

INVx1_ASAP7_75t_L g14809 ( 
.A(n_13095),
.Y(n_14809)
);

INVx2_ASAP7_75t_L g14810 ( 
.A(n_12850),
.Y(n_14810)
);

AOI22xp5_ASAP7_75t_L g14811 ( 
.A1(n_13003),
.A2(n_1472),
.B1(n_1470),
.B2(n_1471),
.Y(n_14811)
);

NAND2xp5_ASAP7_75t_L g14812 ( 
.A(n_13495),
.B(n_1470),
.Y(n_14812)
);

AND2x2_ASAP7_75t_L g14813 ( 
.A(n_13613),
.B(n_13614),
.Y(n_14813)
);

INVx1_ASAP7_75t_L g14814 ( 
.A(n_13232),
.Y(n_14814)
);

NOR2xp33_ASAP7_75t_L g14815 ( 
.A(n_13486),
.B(n_1471),
.Y(n_14815)
);

NAND2xp5_ASAP7_75t_L g14816 ( 
.A(n_13511),
.B(n_1472),
.Y(n_14816)
);

AOI22xp5_ASAP7_75t_L g14817 ( 
.A1(n_13064),
.A2(n_1475),
.B1(n_1473),
.B2(n_1474),
.Y(n_14817)
);

NAND2xp5_ASAP7_75t_L g14818 ( 
.A(n_12886),
.B(n_1473),
.Y(n_14818)
);

INVx1_ASAP7_75t_L g14819 ( 
.A(n_12887),
.Y(n_14819)
);

NAND2xp5_ASAP7_75t_L g14820 ( 
.A(n_12906),
.B(n_1474),
.Y(n_14820)
);

NOR2xp33_ASAP7_75t_L g14821 ( 
.A(n_12860),
.B(n_1475),
.Y(n_14821)
);

INVxp33_ASAP7_75t_SL g14822 ( 
.A(n_12897),
.Y(n_14822)
);

INVx2_ASAP7_75t_L g14823 ( 
.A(n_12927),
.Y(n_14823)
);

NAND2xp5_ASAP7_75t_L g14824 ( 
.A(n_12938),
.B(n_1476),
.Y(n_14824)
);

NAND2xp5_ASAP7_75t_L g14825 ( 
.A(n_13320),
.B(n_1476),
.Y(n_14825)
);

AND2x2_ASAP7_75t_SL g14826 ( 
.A(n_13620),
.B(n_1477),
.Y(n_14826)
);

AOI22xp33_ASAP7_75t_L g14827 ( 
.A1(n_12945),
.A2(n_1479),
.B1(n_1477),
.B2(n_1478),
.Y(n_14827)
);

A2O1A1Ixp33_ASAP7_75t_L g14828 ( 
.A1(n_12946),
.A2(n_1480),
.B(n_1478),
.C(n_1479),
.Y(n_14828)
);

NAND2xp5_ASAP7_75t_L g14829 ( 
.A(n_13627),
.B(n_1480),
.Y(n_14829)
);

INVx1_ASAP7_75t_L g14830 ( 
.A(n_12802),
.Y(n_14830)
);

NAND2xp5_ASAP7_75t_L g14831 ( 
.A(n_13628),
.B(n_1481),
.Y(n_14831)
);

INVx2_ASAP7_75t_L g14832 ( 
.A(n_12814),
.Y(n_14832)
);

CKINVDCx5p33_ASAP7_75t_R g14833 ( 
.A(n_13239),
.Y(n_14833)
);

AND2x2_ASAP7_75t_L g14834 ( 
.A(n_13642),
.B(n_1481),
.Y(n_14834)
);

NAND2xp5_ASAP7_75t_L g14835 ( 
.A(n_13647),
.B(n_1482),
.Y(n_14835)
);

INVx1_ASAP7_75t_L g14836 ( 
.A(n_12816),
.Y(n_14836)
);

O2A1O1Ixp33_ASAP7_75t_L g14837 ( 
.A1(n_13648),
.A2(n_1484),
.B(n_1482),
.C(n_1483),
.Y(n_14837)
);

INVx2_ASAP7_75t_L g14838 ( 
.A(n_12830),
.Y(n_14838)
);

NAND2xp33_ASAP7_75t_SL g14839 ( 
.A(n_13649),
.B(n_1483),
.Y(n_14839)
);

NAND2xp5_ASAP7_75t_L g14840 ( 
.A(n_13658),
.B(n_13662),
.Y(n_14840)
);

INVx1_ASAP7_75t_L g14841 ( 
.A(n_13672),
.Y(n_14841)
);

INVx1_ASAP7_75t_L g14842 ( 
.A(n_13681),
.Y(n_14842)
);

INVx2_ASAP7_75t_L g14843 ( 
.A(n_13685),
.Y(n_14843)
);

INVx1_ASAP7_75t_L g14844 ( 
.A(n_13701),
.Y(n_14844)
);

INVxp67_ASAP7_75t_L g14845 ( 
.A(n_13705),
.Y(n_14845)
);

AO22x1_ASAP7_75t_L g14846 ( 
.A1(n_13708),
.A2(n_1486),
.B1(n_1484),
.B2(n_1485),
.Y(n_14846)
);

INVx1_ASAP7_75t_L g14847 ( 
.A(n_13714),
.Y(n_14847)
);

INVx1_ASAP7_75t_L g14848 ( 
.A(n_13718),
.Y(n_14848)
);

HB1xp67_ASAP7_75t_L g14849 ( 
.A(n_13727),
.Y(n_14849)
);

INVx2_ASAP7_75t_L g14850 ( 
.A(n_13734),
.Y(n_14850)
);

INVxp67_ASAP7_75t_L g14851 ( 
.A(n_13740),
.Y(n_14851)
);

BUFx2_ASAP7_75t_L g14852 ( 
.A(n_13899),
.Y(n_14852)
);

BUFx3_ASAP7_75t_L g14853 ( 
.A(n_13238),
.Y(n_14853)
);

INVx2_ASAP7_75t_L g14854 ( 
.A(n_13745),
.Y(n_14854)
);

INVx1_ASAP7_75t_L g14855 ( 
.A(n_13756),
.Y(n_14855)
);

NAND2xp5_ASAP7_75t_L g14856 ( 
.A(n_13757),
.B(n_1487),
.Y(n_14856)
);

INVx2_ASAP7_75t_L g14857 ( 
.A(n_13762),
.Y(n_14857)
);

HB1xp67_ASAP7_75t_L g14858 ( 
.A(n_13764),
.Y(n_14858)
);

INVx2_ASAP7_75t_L g14859 ( 
.A(n_13770),
.Y(n_14859)
);

CKINVDCx20_ASAP7_75t_R g14860 ( 
.A(n_12844),
.Y(n_14860)
);

INVx1_ASAP7_75t_L g14861 ( 
.A(n_13776),
.Y(n_14861)
);

AND2x2_ASAP7_75t_L g14862 ( 
.A(n_13778),
.B(n_13780),
.Y(n_14862)
);

NAND2xp5_ASAP7_75t_L g14863 ( 
.A(n_14188),
.B(n_14126),
.Y(n_14863)
);

BUFx6f_ASAP7_75t_SL g14864 ( 
.A(n_14067),
.Y(n_14864)
);

OAI22x1_ASAP7_75t_L g14865 ( 
.A1(n_13957),
.A2(n_13793),
.B1(n_13802),
.B2(n_13781),
.Y(n_14865)
);

A2O1A1Ixp33_ASAP7_75t_L g14866 ( 
.A1(n_13912),
.A2(n_12949),
.B(n_12956),
.C(n_12948),
.Y(n_14866)
);

AOI21xp5_ASAP7_75t_L g14867 ( 
.A1(n_14445),
.A2(n_12978),
.B(n_12974),
.Y(n_14867)
);

NAND2xp5_ASAP7_75t_L g14868 ( 
.A(n_14129),
.B(n_13807),
.Y(n_14868)
);

NOR2xp67_ASAP7_75t_L g14869 ( 
.A(n_14608),
.B(n_13810),
.Y(n_14869)
);

NAND2xp5_ASAP7_75t_L g14870 ( 
.A(n_13921),
.B(n_13816),
.Y(n_14870)
);

OAI22xp5_ASAP7_75t_L g14871 ( 
.A1(n_14539),
.A2(n_13831),
.B1(n_13837),
.B2(n_13825),
.Y(n_14871)
);

HB1xp67_ASAP7_75t_L g14872 ( 
.A(n_14063),
.Y(n_14872)
);

AO31x2_ASAP7_75t_L g14873 ( 
.A1(n_14416),
.A2(n_12984),
.A3(n_12988),
.B(n_12979),
.Y(n_14873)
);

NAND2xp5_ASAP7_75t_L g14874 ( 
.A(n_14002),
.B(n_13839),
.Y(n_14874)
);

CKINVDCx20_ASAP7_75t_R g14875 ( 
.A(n_14236),
.Y(n_14875)
);

INVx2_ASAP7_75t_L g14876 ( 
.A(n_13961),
.Y(n_14876)
);

NOR2xp33_ASAP7_75t_L g14877 ( 
.A(n_13917),
.B(n_13843),
.Y(n_14877)
);

AOI21xp5_ASAP7_75t_L g14878 ( 
.A1(n_14597),
.A2(n_13004),
.B(n_13002),
.Y(n_14878)
);

OAI21xp5_ASAP7_75t_L g14879 ( 
.A1(n_14458),
.A2(n_13242),
.B(n_13244),
.Y(n_14879)
);

BUFx3_ASAP7_75t_L g14880 ( 
.A(n_14012),
.Y(n_14880)
);

NAND2xp5_ASAP7_75t_SL g14881 ( 
.A(n_13951),
.B(n_14540),
.Y(n_14881)
);

OA21x2_ASAP7_75t_L g14882 ( 
.A1(n_14411),
.A2(n_14130),
.B(n_14175),
.Y(n_14882)
);

INVx2_ASAP7_75t_L g14883 ( 
.A(n_14134),
.Y(n_14883)
);

CKINVDCx5p33_ASAP7_75t_R g14884 ( 
.A(n_13944),
.Y(n_14884)
);

INVx6_ASAP7_75t_L g14885 ( 
.A(n_14018),
.Y(n_14885)
);

OAI21x1_ASAP7_75t_L g14886 ( 
.A1(n_14420),
.A2(n_13856),
.B(n_13854),
.Y(n_14886)
);

NOR2xp67_ASAP7_75t_SL g14887 ( 
.A(n_13951),
.B(n_13869),
.Y(n_14887)
);

AO32x2_ASAP7_75t_L g14888 ( 
.A1(n_14021),
.A2(n_13894),
.A3(n_13871),
.B1(n_13027),
.B2(n_13028),
.Y(n_14888)
);

OAI21xp5_ASAP7_75t_L g14889 ( 
.A1(n_14464),
.A2(n_13020),
.B(n_13011),
.Y(n_14889)
);

NOR2xp33_ASAP7_75t_L g14890 ( 
.A(n_14186),
.B(n_13380),
.Y(n_14890)
);

O2A1O1Ixp33_ASAP7_75t_L g14891 ( 
.A1(n_14391),
.A2(n_13043),
.B(n_13047),
.C(n_13039),
.Y(n_14891)
);

AND2x4_ASAP7_75t_L g14892 ( 
.A(n_14031),
.B(n_13532),
.Y(n_14892)
);

A2O1A1Ixp33_ASAP7_75t_L g14893 ( 
.A1(n_14078),
.A2(n_13076),
.B(n_13079),
.C(n_13075),
.Y(n_14893)
);

AOI22xp33_ASAP7_75t_L g14894 ( 
.A1(n_14677),
.A2(n_13085),
.B1(n_13096),
.B2(n_13094),
.Y(n_14894)
);

AOI21xp5_ASAP7_75t_L g14895 ( 
.A1(n_14603),
.A2(n_13109),
.B(n_13106),
.Y(n_14895)
);

INVxp67_ASAP7_75t_L g14896 ( 
.A(n_14388),
.Y(n_14896)
);

AOI21x1_ASAP7_75t_L g14897 ( 
.A1(n_14311),
.A2(n_13575),
.B(n_13568),
.Y(n_14897)
);

INVx2_ASAP7_75t_L g14898 ( 
.A(n_14137),
.Y(n_14898)
);

A2O1A1Ixp33_ASAP7_75t_L g14899 ( 
.A1(n_13916),
.A2(n_13124),
.B(n_13128),
.C(n_13112),
.Y(n_14899)
);

BUFx3_ASAP7_75t_L g14900 ( 
.A(n_14154),
.Y(n_14900)
);

INVx1_ASAP7_75t_L g14901 ( 
.A(n_14052),
.Y(n_14901)
);

INVx1_ASAP7_75t_L g14902 ( 
.A(n_13906),
.Y(n_14902)
);

A2O1A1Ixp33_ASAP7_75t_L g14903 ( 
.A1(n_14092),
.A2(n_13154),
.B(n_13139),
.C(n_13172),
.Y(n_14903)
);

O2A1O1Ixp33_ASAP7_75t_SL g14904 ( 
.A1(n_14250),
.A2(n_12856),
.B(n_12866),
.C(n_12857),
.Y(n_14904)
);

INVx1_ASAP7_75t_L g14905 ( 
.A(n_13927),
.Y(n_14905)
);

BUFx2_ASAP7_75t_L g14906 ( 
.A(n_14136),
.Y(n_14906)
);

NAND2xp5_ASAP7_75t_L g14907 ( 
.A(n_14099),
.B(n_14120),
.Y(n_14907)
);

AOI221x1_ASAP7_75t_L g14908 ( 
.A1(n_13969),
.A2(n_13245),
.B1(n_13263),
.B2(n_13262),
.C(n_13260),
.Y(n_14908)
);

AO31x2_ASAP7_75t_L g14909 ( 
.A1(n_14423),
.A2(n_13273),
.A3(n_13293),
.B(n_13268),
.Y(n_14909)
);

OAI21xp5_ASAP7_75t_L g14910 ( 
.A1(n_14705),
.A2(n_13311),
.B(n_13300),
.Y(n_14910)
);

AOI21xp5_ASAP7_75t_L g14911 ( 
.A1(n_14840),
.A2(n_13323),
.B(n_13319),
.Y(n_14911)
);

OAI21xp5_ASAP7_75t_L g14912 ( 
.A1(n_14024),
.A2(n_13329),
.B(n_13327),
.Y(n_14912)
);

NAND2xp5_ASAP7_75t_L g14913 ( 
.A(n_14163),
.B(n_13199),
.Y(n_14913)
);

AOI221xp5_ASAP7_75t_L g14914 ( 
.A1(n_14656),
.A2(n_13178),
.B1(n_13174),
.B2(n_13337),
.C(n_13330),
.Y(n_14914)
);

AOI21xp5_ASAP7_75t_L g14915 ( 
.A1(n_14600),
.A2(n_13344),
.B(n_13340),
.Y(n_14915)
);

INVx1_ASAP7_75t_L g14916 ( 
.A(n_13938),
.Y(n_14916)
);

HB1xp67_ASAP7_75t_L g14917 ( 
.A(n_13934),
.Y(n_14917)
);

OAI21x1_ASAP7_75t_L g14918 ( 
.A1(n_14422),
.A2(n_13206),
.B(n_13346),
.Y(n_14918)
);

NAND2xp5_ASAP7_75t_L g14919 ( 
.A(n_14438),
.B(n_13347),
.Y(n_14919)
);

OAI22xp5_ASAP7_75t_L g14920 ( 
.A1(n_14135),
.A2(n_12868),
.B1(n_12871),
.B2(n_12870),
.Y(n_14920)
);

OAI21xp33_ASAP7_75t_L g14921 ( 
.A1(n_14353),
.A2(n_13351),
.B(n_13349),
.Y(n_14921)
);

OAI22x1_ASAP7_75t_L g14922 ( 
.A1(n_14616),
.A2(n_1489),
.B1(n_1487),
.B2(n_1488),
.Y(n_14922)
);

NAND3xp33_ASAP7_75t_SL g14923 ( 
.A(n_14008),
.B(n_13379),
.C(n_13362),
.Y(n_14923)
);

NAND2xp5_ASAP7_75t_L g14924 ( 
.A(n_14143),
.B(n_13475),
.Y(n_14924)
);

AOI31xp67_ASAP7_75t_L g14925 ( 
.A1(n_14679),
.A2(n_1490),
.A3(n_1488),
.B(n_1489),
.Y(n_14925)
);

OAI21xp5_ASAP7_75t_SL g14926 ( 
.A1(n_14292),
.A2(n_12878),
.B(n_12875),
.Y(n_14926)
);

OR2x2_ASAP7_75t_L g14927 ( 
.A(n_14014),
.B(n_13484),
.Y(n_14927)
);

O2A1O1Ixp33_ASAP7_75t_L g14928 ( 
.A1(n_14729),
.A2(n_13512),
.B(n_13435),
.C(n_13436),
.Y(n_14928)
);

INVx2_ASAP7_75t_SL g14929 ( 
.A(n_14326),
.Y(n_14929)
);

BUFx3_ASAP7_75t_L g14930 ( 
.A(n_14405),
.Y(n_14930)
);

AOI21xp5_ASAP7_75t_L g14931 ( 
.A1(n_14586),
.A2(n_13581),
.B(n_13212),
.Y(n_14931)
);

NAND3xp33_ASAP7_75t_L g14932 ( 
.A(n_14713),
.B(n_14455),
.C(n_14619),
.Y(n_14932)
);

AO32x2_ASAP7_75t_L g14933 ( 
.A1(n_14122),
.A2(n_13404),
.A3(n_13417),
.B1(n_13397),
.B2(n_13394),
.Y(n_14933)
);

AOI21xp5_ASAP7_75t_L g14934 ( 
.A1(n_14550),
.A2(n_13467),
.B(n_13442),
.Y(n_14934)
);

AOI21xp5_ASAP7_75t_L g14935 ( 
.A1(n_14700),
.A2(n_13472),
.B(n_13469),
.Y(n_14935)
);

OR2x2_ASAP7_75t_SL g14936 ( 
.A(n_14323),
.B(n_13962),
.Y(n_14936)
);

NOR4xp25_ASAP7_75t_L g14937 ( 
.A(n_13919),
.B(n_1493),
.C(n_1491),
.D(n_1492),
.Y(n_14937)
);

AOI21xp5_ASAP7_75t_L g14938 ( 
.A1(n_14720),
.A2(n_13526),
.B(n_13523),
.Y(n_14938)
);

INVx1_ASAP7_75t_L g14939 ( 
.A(n_13949),
.Y(n_14939)
);

A2O1A1Ixp33_ASAP7_75t_L g14940 ( 
.A1(n_14572),
.A2(n_14759),
.B(n_14768),
.C(n_14764),
.Y(n_14940)
);

BUFx2_ASAP7_75t_L g14941 ( 
.A(n_14043),
.Y(n_14941)
);

OAI21x1_ASAP7_75t_L g14942 ( 
.A1(n_14452),
.A2(n_13554),
.B(n_13534),
.Y(n_14942)
);

AND2x2_ASAP7_75t_L g14943 ( 
.A(n_13937),
.B(n_13485),
.Y(n_14943)
);

INVx2_ASAP7_75t_L g14944 ( 
.A(n_14156),
.Y(n_14944)
);

AOI21xp5_ASAP7_75t_L g14945 ( 
.A1(n_14686),
.A2(n_13504),
.B(n_13493),
.Y(n_14945)
);

INVx1_ASAP7_75t_L g14946 ( 
.A(n_13950),
.Y(n_14946)
);

A2O1A1Ixp33_ASAP7_75t_L g14947 ( 
.A1(n_14762),
.A2(n_12817),
.B(n_13509),
.C(n_13507),
.Y(n_14947)
);

INVx8_ASAP7_75t_L g14948 ( 
.A(n_14366),
.Y(n_14948)
);

AND2x4_ASAP7_75t_L g14949 ( 
.A(n_14064),
.B(n_1493),
.Y(n_14949)
);

AOI21xp5_ASAP7_75t_L g14950 ( 
.A1(n_14441),
.A2(n_5899),
.B(n_5898),
.Y(n_14950)
);

CKINVDCx5p33_ASAP7_75t_R g14951 ( 
.A(n_13954),
.Y(n_14951)
);

AOI21xp5_ASAP7_75t_L g14952 ( 
.A1(n_14444),
.A2(n_5901),
.B(n_5900),
.Y(n_14952)
);

AND2x2_ASAP7_75t_L g14953 ( 
.A(n_13946),
.B(n_1494),
.Y(n_14953)
);

NOR2xp67_ASAP7_75t_L g14954 ( 
.A(n_14716),
.B(n_1495),
.Y(n_14954)
);

AOI221xp5_ASAP7_75t_L g14955 ( 
.A1(n_14511),
.A2(n_1497),
.B1(n_1495),
.B2(n_1496),
.C(n_1498),
.Y(n_14955)
);

NOR2x1_ASAP7_75t_SL g14956 ( 
.A(n_13951),
.B(n_1496),
.Y(n_14956)
);

OAI21x1_ASAP7_75t_L g14957 ( 
.A1(n_14467),
.A2(n_1497),
.B(n_1498),
.Y(n_14957)
);

OA21x2_ASAP7_75t_L g14958 ( 
.A1(n_14133),
.A2(n_1499),
.B(n_1500),
.Y(n_14958)
);

INVx2_ASAP7_75t_L g14959 ( 
.A(n_13953),
.Y(n_14959)
);

INVx1_ASAP7_75t_L g14960 ( 
.A(n_13958),
.Y(n_14960)
);

INVx1_ASAP7_75t_L g14961 ( 
.A(n_13965),
.Y(n_14961)
);

OAI22xp33_ASAP7_75t_L g14962 ( 
.A1(n_14609),
.A2(n_1501),
.B1(n_1499),
.B2(n_1500),
.Y(n_14962)
);

O2A1O1Ixp5_ASAP7_75t_SL g14963 ( 
.A1(n_14408),
.A2(n_14412),
.B(n_14424),
.C(n_14442),
.Y(n_14963)
);

OAI21x1_ASAP7_75t_SL g14964 ( 
.A1(n_14620),
.A2(n_1502),
.B(n_1503),
.Y(n_14964)
);

OAI22xp5_ASAP7_75t_L g14965 ( 
.A1(n_14200),
.A2(n_1505),
.B1(n_1502),
.B2(n_1504),
.Y(n_14965)
);

INVx2_ASAP7_75t_SL g14966 ( 
.A(n_14058),
.Y(n_14966)
);

OAI21x1_ASAP7_75t_L g14967 ( 
.A1(n_14382),
.A2(n_1504),
.B(n_1505),
.Y(n_14967)
);

AOI221x1_ASAP7_75t_L g14968 ( 
.A1(n_14632),
.A2(n_1508),
.B1(n_1506),
.B2(n_1507),
.C(n_1509),
.Y(n_14968)
);

NAND2xp5_ASAP7_75t_L g14969 ( 
.A(n_13986),
.B(n_1506),
.Y(n_14969)
);

AO31x2_ASAP7_75t_L g14970 ( 
.A1(n_14394),
.A2(n_1511),
.A3(n_1508),
.B(n_1510),
.Y(n_14970)
);

OAI21xp5_ASAP7_75t_L g14971 ( 
.A1(n_14747),
.A2(n_1510),
.B(n_1511),
.Y(n_14971)
);

BUFx4f_ASAP7_75t_L g14972 ( 
.A(n_13960),
.Y(n_14972)
);

AND2x2_ASAP7_75t_L g14973 ( 
.A(n_14095),
.B(n_1512),
.Y(n_14973)
);

OAI21x1_ASAP7_75t_L g14974 ( 
.A1(n_14417),
.A2(n_1512),
.B(n_1513),
.Y(n_14974)
);

NAND2xp33_ASAP7_75t_L g14975 ( 
.A(n_14528),
.B(n_1513),
.Y(n_14975)
);

NAND2xp5_ASAP7_75t_L g14976 ( 
.A(n_13987),
.B(n_1514),
.Y(n_14976)
);

OAI21x1_ASAP7_75t_L g14977 ( 
.A1(n_14418),
.A2(n_1514),
.B(n_1515),
.Y(n_14977)
);

HB1xp67_ASAP7_75t_L g14978 ( 
.A(n_14030),
.Y(n_14978)
);

AOI21xp5_ASAP7_75t_L g14979 ( 
.A1(n_14397),
.A2(n_5903),
.B(n_5902),
.Y(n_14979)
);

O2A1O1Ixp33_ASAP7_75t_L g14980 ( 
.A1(n_14055),
.A2(n_1517),
.B(n_1515),
.C(n_1516),
.Y(n_14980)
);

BUFx6f_ASAP7_75t_L g14981 ( 
.A(n_14307),
.Y(n_14981)
);

AOI221x1_ASAP7_75t_L g14982 ( 
.A1(n_14127),
.A2(n_1518),
.B1(n_1516),
.B2(n_1517),
.C(n_1519),
.Y(n_14982)
);

INVx1_ASAP7_75t_SL g14983 ( 
.A(n_14149),
.Y(n_14983)
);

BUFx3_ASAP7_75t_L g14984 ( 
.A(n_14336),
.Y(n_14984)
);

OAI22xp5_ASAP7_75t_L g14985 ( 
.A1(n_14782),
.A2(n_1520),
.B1(n_1518),
.B2(n_1519),
.Y(n_14985)
);

OAI21xp5_ASAP7_75t_SL g14986 ( 
.A1(n_14001),
.A2(n_1520),
.B(n_1521),
.Y(n_14986)
);

AO32x2_ASAP7_75t_L g14987 ( 
.A1(n_14389),
.A2(n_1523),
.A3(n_1521),
.B1(n_1522),
.B2(n_1524),
.Y(n_14987)
);

INVx4_ASAP7_75t_L g14988 ( 
.A(n_13968),
.Y(n_14988)
);

INVx1_ASAP7_75t_L g14989 ( 
.A(n_13967),
.Y(n_14989)
);

AOI21xp5_ASAP7_75t_L g14990 ( 
.A1(n_14839),
.A2(n_5908),
.B(n_5906),
.Y(n_14990)
);

OAI21x1_ASAP7_75t_L g14991 ( 
.A1(n_14425),
.A2(n_1522),
.B(n_1523),
.Y(n_14991)
);

AO21x1_ASAP7_75t_L g14992 ( 
.A1(n_14479),
.A2(n_14487),
.B(n_14485),
.Y(n_14992)
);

INVx1_ASAP7_75t_L g14993 ( 
.A(n_13977),
.Y(n_14993)
);

OAI21xp5_ASAP7_75t_L g14994 ( 
.A1(n_14845),
.A2(n_1525),
.B(n_1526),
.Y(n_14994)
);

AND2x2_ASAP7_75t_L g14995 ( 
.A(n_13928),
.B(n_13976),
.Y(n_14995)
);

INVx2_ASAP7_75t_L g14996 ( 
.A(n_14003),
.Y(n_14996)
);

NOR2xp33_ASAP7_75t_L g14997 ( 
.A(n_14556),
.B(n_1525),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_14076),
.Y(n_14998)
);

INVx1_ASAP7_75t_L g14999 ( 
.A(n_14079),
.Y(n_14999)
);

O2A1O1Ixp33_ASAP7_75t_L g15000 ( 
.A1(n_14139),
.A2(n_1528),
.B(n_1526),
.C(n_1527),
.Y(n_15000)
);

OAI21xp5_ASAP7_75t_L g15001 ( 
.A1(n_14851),
.A2(n_1527),
.B(n_1529),
.Y(n_15001)
);

AOI21xp5_ASAP7_75t_L g15002 ( 
.A1(n_14858),
.A2(n_5910),
.B(n_5909),
.Y(n_15002)
);

OAI21x1_ASAP7_75t_L g15003 ( 
.A1(n_14535),
.A2(n_1529),
.B(n_1530),
.Y(n_15003)
);

NAND3xp33_ASAP7_75t_SL g15004 ( 
.A(n_14406),
.B(n_1530),
.C(n_1531),
.Y(n_15004)
);

BUFx6f_ASAP7_75t_L g15005 ( 
.A(n_14307),
.Y(n_15005)
);

OAI21x1_ASAP7_75t_L g15006 ( 
.A1(n_14544),
.A2(n_1531),
.B(n_1532),
.Y(n_15006)
);

NOR2xp33_ASAP7_75t_L g15007 ( 
.A(n_13925),
.B(n_1532),
.Y(n_15007)
);

INVx1_ASAP7_75t_L g15008 ( 
.A(n_14084),
.Y(n_15008)
);

INVx1_ASAP7_75t_L g15009 ( 
.A(n_14056),
.Y(n_15009)
);

O2A1O1Ixp33_ASAP7_75t_L g15010 ( 
.A1(n_14141),
.A2(n_1535),
.B(n_1533),
.C(n_1534),
.Y(n_15010)
);

BUFx6f_ASAP7_75t_L g15011 ( 
.A(n_14308),
.Y(n_15011)
);

A2O1A1Ixp33_ASAP7_75t_L g15012 ( 
.A1(n_14774),
.A2(n_1535),
.B(n_1533),
.C(n_1534),
.Y(n_15012)
);

BUFx2_ASAP7_75t_L g15013 ( 
.A(n_14274),
.Y(n_15013)
);

AOI21xp5_ASAP7_75t_L g15014 ( 
.A1(n_14849),
.A2(n_5912),
.B(n_5911),
.Y(n_15014)
);

AND2x2_ASAP7_75t_L g15015 ( 
.A(n_14205),
.B(n_1536),
.Y(n_15015)
);

AOI21xp5_ASAP7_75t_L g15016 ( 
.A1(n_14427),
.A2(n_5914),
.B(n_5913),
.Y(n_15016)
);

AO21x2_ASAP7_75t_L g15017 ( 
.A1(n_14522),
.A2(n_1536),
.B(n_1537),
.Y(n_15017)
);

A2O1A1Ixp33_ASAP7_75t_L g15018 ( 
.A1(n_14791),
.A2(n_1539),
.B(n_1537),
.C(n_1538),
.Y(n_15018)
);

AO21x2_ASAP7_75t_L g15019 ( 
.A1(n_14415),
.A2(n_1538),
.B(n_1539),
.Y(n_15019)
);

OAI21xp5_ASAP7_75t_L g15020 ( 
.A1(n_14745),
.A2(n_1540),
.B(n_1541),
.Y(n_15020)
);

BUFx12f_ASAP7_75t_L g15021 ( 
.A(n_14005),
.Y(n_15021)
);

AOI221x1_ASAP7_75t_L g15022 ( 
.A1(n_13940),
.A2(n_1542),
.B1(n_1540),
.B2(n_1541),
.C(n_1543),
.Y(n_15022)
);

CKINVDCx11_ASAP7_75t_R g15023 ( 
.A(n_14066),
.Y(n_15023)
);

INVxp67_ASAP7_75t_SL g15024 ( 
.A(n_14339),
.Y(n_15024)
);

AND2x2_ASAP7_75t_L g15025 ( 
.A(n_14257),
.B(n_1542),
.Y(n_15025)
);

AOI21xp5_ASAP7_75t_L g15026 ( 
.A1(n_14716),
.A2(n_5916),
.B(n_5915),
.Y(n_15026)
);

INVx1_ASAP7_75t_L g15027 ( 
.A(n_14069),
.Y(n_15027)
);

OAI21x1_ASAP7_75t_L g15028 ( 
.A1(n_14564),
.A2(n_1543),
.B(n_1544),
.Y(n_15028)
);

INVx1_ASAP7_75t_L g15029 ( 
.A(n_14070),
.Y(n_15029)
);

AO31x2_ASAP7_75t_L g15030 ( 
.A1(n_14465),
.A2(n_14473),
.A3(n_14440),
.B(n_14428),
.Y(n_15030)
);

AOI221xp5_ASAP7_75t_SL g15031 ( 
.A1(n_14495),
.A2(n_14503),
.B1(n_14508),
.B2(n_14210),
.C(n_14300),
.Y(n_15031)
);

INVx2_ASAP7_75t_L g15032 ( 
.A(n_14094),
.Y(n_15032)
);

NAND2xp5_ASAP7_75t_L g15033 ( 
.A(n_14145),
.B(n_1544),
.Y(n_15033)
);

INVx2_ASAP7_75t_L g15034 ( 
.A(n_14098),
.Y(n_15034)
);

OAI22xp5_ASAP7_75t_L g15035 ( 
.A1(n_14800),
.A2(n_1547),
.B1(n_1545),
.B2(n_1546),
.Y(n_15035)
);

NOR2xp33_ASAP7_75t_SL g15036 ( 
.A(n_13902),
.B(n_1545),
.Y(n_15036)
);

NAND2x1p5_ASAP7_75t_L g15037 ( 
.A(n_14716),
.B(n_5918),
.Y(n_15037)
);

NOR2xp33_ASAP7_75t_SL g15038 ( 
.A(n_13913),
.B(n_1546),
.Y(n_15038)
);

NAND2xp5_ASAP7_75t_SL g15039 ( 
.A(n_14681),
.B(n_1547),
.Y(n_15039)
);

NAND2xp5_ASAP7_75t_L g15040 ( 
.A(n_14361),
.B(n_1548),
.Y(n_15040)
);

OR2x2_ASAP7_75t_L g15041 ( 
.A(n_14023),
.B(n_1548),
.Y(n_15041)
);

O2A1O1Ixp33_ASAP7_75t_SL g15042 ( 
.A1(n_14548),
.A2(n_1551),
.B(n_1549),
.C(n_1550),
.Y(n_15042)
);

OAI21xp5_ASAP7_75t_L g15043 ( 
.A1(n_14828),
.A2(n_1549),
.B(n_1550),
.Y(n_15043)
);

BUFx12f_ASAP7_75t_L g15044 ( 
.A(n_14074),
.Y(n_15044)
);

INVx2_ASAP7_75t_SL g15045 ( 
.A(n_14384),
.Y(n_15045)
);

AO31x2_ASAP7_75t_L g15046 ( 
.A1(n_14446),
.A2(n_1553),
.A3(n_1551),
.B(n_1552),
.Y(n_15046)
);

NAND2xp5_ASAP7_75t_L g15047 ( 
.A(n_14365),
.B(n_1552),
.Y(n_15047)
);

AO32x2_ASAP7_75t_L g15048 ( 
.A1(n_14565),
.A2(n_1555),
.A3(n_1553),
.B1(n_1554),
.B2(n_1557),
.Y(n_15048)
);

OAI22xp5_ASAP7_75t_L g15049 ( 
.A1(n_14162),
.A2(n_1557),
.B1(n_1554),
.B2(n_1555),
.Y(n_15049)
);

NOR2x1_ASAP7_75t_L g15050 ( 
.A(n_14087),
.B(n_1558),
.Y(n_15050)
);

AOI21xp5_ASAP7_75t_L g15051 ( 
.A1(n_14650),
.A2(n_5920),
.B(n_5919),
.Y(n_15051)
);

A2O1A1Ixp33_ASAP7_75t_L g15052 ( 
.A1(n_14792),
.A2(n_1561),
.B(n_1559),
.C(n_1560),
.Y(n_15052)
);

OAI21xp5_ASAP7_75t_L g15053 ( 
.A1(n_14772),
.A2(n_1559),
.B(n_1560),
.Y(n_15053)
);

A2O1A1Ixp33_ASAP7_75t_L g15054 ( 
.A1(n_14797),
.A2(n_1563),
.B(n_1561),
.C(n_1562),
.Y(n_15054)
);

INVx2_ASAP7_75t_SL g15055 ( 
.A(n_14395),
.Y(n_15055)
);

NAND2xp5_ASAP7_75t_L g15056 ( 
.A(n_14324),
.B(n_14325),
.Y(n_15056)
);

AOI21xp5_ASAP7_75t_L g15057 ( 
.A1(n_14852),
.A2(n_5923),
.B(n_5921),
.Y(n_15057)
);

BUFx5_ASAP7_75t_L g15058 ( 
.A(n_14626),
.Y(n_15058)
);

CKINVDCx20_ASAP7_75t_R g15059 ( 
.A(n_14281),
.Y(n_15059)
);

CKINVDCx5p33_ASAP7_75t_R g15060 ( 
.A(n_14047),
.Y(n_15060)
);

AND2x2_ASAP7_75t_L g15061 ( 
.A(n_14106),
.B(n_14449),
.Y(n_15061)
);

OAI21x1_ASAP7_75t_L g15062 ( 
.A1(n_14593),
.A2(n_1562),
.B(n_1563),
.Y(n_15062)
);

AOI21xp5_ASAP7_75t_L g15063 ( 
.A1(n_14784),
.A2(n_5925),
.B(n_5924),
.Y(n_15063)
);

A2O1A1Ixp33_ASAP7_75t_L g15064 ( 
.A1(n_14804),
.A2(n_1566),
.B(n_1564),
.C(n_1565),
.Y(n_15064)
);

O2A1O1Ixp5_ASAP7_75t_L g15065 ( 
.A1(n_14342),
.A2(n_1567),
.B(n_1565),
.C(n_1566),
.Y(n_15065)
);

OAI21x1_ASAP7_75t_L g15066 ( 
.A1(n_14614),
.A2(n_1567),
.B(n_1568),
.Y(n_15066)
);

OAI21xp5_ASAP7_75t_L g15067 ( 
.A1(n_14809),
.A2(n_1568),
.B(n_1569),
.Y(n_15067)
);

OAI21x1_ASAP7_75t_L g15068 ( 
.A1(n_14187),
.A2(n_1569),
.B(n_1570),
.Y(n_15068)
);

OAI21x1_ASAP7_75t_L g15069 ( 
.A1(n_14830),
.A2(n_1570),
.B(n_1571),
.Y(n_15069)
);

AOI21xp5_ASAP7_75t_L g15070 ( 
.A1(n_14813),
.A2(n_5930),
.B(n_5928),
.Y(n_15070)
);

INVx1_ASAP7_75t_L g15071 ( 
.A(n_14073),
.Y(n_15071)
);

NAND2xp5_ASAP7_75t_SL g15072 ( 
.A(n_14778),
.B(n_14543),
.Y(n_15072)
);

INVx1_ASAP7_75t_L g15073 ( 
.A(n_13904),
.Y(n_15073)
);

OA21x2_ASAP7_75t_L g15074 ( 
.A1(n_14157),
.A2(n_1571),
.B(n_1572),
.Y(n_15074)
);

BUFx6f_ASAP7_75t_L g15075 ( 
.A(n_14308),
.Y(n_15075)
);

INVx3_ASAP7_75t_L g15076 ( 
.A(n_14284),
.Y(n_15076)
);

AOI21xp5_ASAP7_75t_L g15077 ( 
.A1(n_14862),
.A2(n_5932),
.B(n_5931),
.Y(n_15077)
);

INVx1_ASAP7_75t_L g15078 ( 
.A(n_13911),
.Y(n_15078)
);

NOR2xp33_ASAP7_75t_L g15079 ( 
.A(n_13956),
.B(n_1573),
.Y(n_15079)
);

INVx2_ASAP7_75t_L g15080 ( 
.A(n_13914),
.Y(n_15080)
);

AOI21xp5_ASAP7_75t_L g15081 ( 
.A1(n_13915),
.A2(n_14676),
.B(n_14554),
.Y(n_15081)
);

INVx2_ASAP7_75t_L g15082 ( 
.A(n_13923),
.Y(n_15082)
);

AOI31xp67_ASAP7_75t_L g15083 ( 
.A1(n_14641),
.A2(n_1576),
.A3(n_1573),
.B(n_1574),
.Y(n_15083)
);

OR2x2_ASAP7_75t_L g15084 ( 
.A(n_14038),
.B(n_1574),
.Y(n_15084)
);

A2O1A1Ixp33_ASAP7_75t_L g15085 ( 
.A1(n_14814),
.A2(n_1578),
.B(n_1576),
.C(n_1577),
.Y(n_15085)
);

INVx1_ASAP7_75t_L g15086 ( 
.A(n_13933),
.Y(n_15086)
);

AO31x2_ASAP7_75t_L g15087 ( 
.A1(n_14533),
.A2(n_1580),
.A3(n_1578),
.B(n_1579),
.Y(n_15087)
);

OAI21x1_ASAP7_75t_L g15088 ( 
.A1(n_14836),
.A2(n_1579),
.B(n_1580),
.Y(n_15088)
);

INVx6_ASAP7_75t_L g15089 ( 
.A(n_14199),
.Y(n_15089)
);

BUFx10_ASAP7_75t_L g15090 ( 
.A(n_14232),
.Y(n_15090)
);

INVx2_ASAP7_75t_L g15091 ( 
.A(n_13942),
.Y(n_15091)
);

INVx2_ASAP7_75t_L g15092 ( 
.A(n_13964),
.Y(n_15092)
);

O2A1O1Ixp5_ASAP7_75t_L g15093 ( 
.A1(n_14517),
.A2(n_1583),
.B(n_1581),
.C(n_1582),
.Y(n_15093)
);

NAND2x1p5_ASAP7_75t_L g15094 ( 
.A(n_14409),
.B(n_5934),
.Y(n_15094)
);

AO31x2_ASAP7_75t_L g15095 ( 
.A1(n_14545),
.A2(n_1586),
.A3(n_1582),
.B(n_1585),
.Y(n_15095)
);

AOI21x1_ASAP7_75t_L g15096 ( 
.A1(n_14604),
.A2(n_1585),
.B(n_1586),
.Y(n_15096)
);

INVx4_ASAP7_75t_L g15097 ( 
.A(n_13970),
.Y(n_15097)
);

OA21x2_ASAP7_75t_L g15098 ( 
.A1(n_14165),
.A2(n_1587),
.B(n_1588),
.Y(n_15098)
);

AOI21xp5_ASAP7_75t_L g15099 ( 
.A1(n_14676),
.A2(n_5936),
.B(n_5935),
.Y(n_15099)
);

AOI22xp5_ASAP7_75t_L g15100 ( 
.A1(n_14278),
.A2(n_1589),
.B1(n_1587),
.B2(n_1588),
.Y(n_15100)
);

AOI21xp5_ASAP7_75t_L g15101 ( 
.A1(n_14790),
.A2(n_5938),
.B(n_5937),
.Y(n_15101)
);

O2A1O1Ixp33_ASAP7_75t_SL g15102 ( 
.A1(n_14560),
.A2(n_1591),
.B(n_1589),
.C(n_1590),
.Y(n_15102)
);

AOI22xp5_ASAP7_75t_L g15103 ( 
.A1(n_14278),
.A2(n_1594),
.B1(n_1592),
.B2(n_1593),
.Y(n_15103)
);

AOI21xp5_ASAP7_75t_L g15104 ( 
.A1(n_14819),
.A2(n_5940),
.B(n_5939),
.Y(n_15104)
);

AO32x2_ASAP7_75t_L g15105 ( 
.A1(n_14022),
.A2(n_14401),
.A3(n_14802),
.B1(n_14338),
.B2(n_14649),
.Y(n_15105)
);

NAND2xp5_ASAP7_75t_L g15106 ( 
.A(n_14337),
.B(n_1592),
.Y(n_15106)
);

INVx3_ASAP7_75t_L g15107 ( 
.A(n_14255),
.Y(n_15107)
);

BUFx3_ASAP7_75t_L g15108 ( 
.A(n_13959),
.Y(n_15108)
);

AND2x4_ASAP7_75t_L g15109 ( 
.A(n_14302),
.B(n_1593),
.Y(n_15109)
);

OAI21x1_ASAP7_75t_L g15110 ( 
.A1(n_14832),
.A2(n_1594),
.B(n_1596),
.Y(n_15110)
);

AOI21xp5_ASAP7_75t_L g15111 ( 
.A1(n_14264),
.A2(n_5942),
.B(n_5941),
.Y(n_15111)
);

INVx2_ASAP7_75t_SL g15112 ( 
.A(n_14182),
.Y(n_15112)
);

NAND2xp5_ASAP7_75t_L g15113 ( 
.A(n_14347),
.B(n_14217),
.Y(n_15113)
);

NAND3xp33_ASAP7_75t_L g15114 ( 
.A(n_14815),
.B(n_1597),
.C(n_1598),
.Y(n_15114)
);

O2A1O1Ixp5_ASAP7_75t_L g15115 ( 
.A1(n_14846),
.A2(n_1599),
.B(n_1597),
.C(n_1598),
.Y(n_15115)
);

INVxp67_ASAP7_75t_L g15116 ( 
.A(n_13975),
.Y(n_15116)
);

AOI21x1_ASAP7_75t_L g15117 ( 
.A1(n_13907),
.A2(n_1599),
.B(n_1601),
.Y(n_15117)
);

CKINVDCx11_ASAP7_75t_R g15118 ( 
.A(n_14150),
.Y(n_15118)
);

BUFx2_ASAP7_75t_L g15119 ( 
.A(n_14367),
.Y(n_15119)
);

INVx1_ASAP7_75t_L g15120 ( 
.A(n_13978),
.Y(n_15120)
);

OAI21xp5_ASAP7_75t_L g15121 ( 
.A1(n_14818),
.A2(n_1601),
.B(n_1602),
.Y(n_15121)
);

AND2x2_ASAP7_75t_L g15122 ( 
.A(n_14168),
.B(n_1602),
.Y(n_15122)
);

AOI21xp5_ASAP7_75t_L g15123 ( 
.A1(n_14359),
.A2(n_5944),
.B(n_5943),
.Y(n_15123)
);

INVx5_ASAP7_75t_L g15124 ( 
.A(n_14214),
.Y(n_15124)
);

INVx3_ASAP7_75t_SL g15125 ( 
.A(n_14013),
.Y(n_15125)
);

AOI21xp5_ASAP7_75t_SL g15126 ( 
.A1(n_14044),
.A2(n_14429),
.B(n_13995),
.Y(n_15126)
);

NAND2xp5_ASAP7_75t_L g15127 ( 
.A(n_14223),
.B(n_1603),
.Y(n_15127)
);

AOI21xp5_ASAP7_75t_L g15128 ( 
.A1(n_14837),
.A2(n_14065),
.B(n_14044),
.Y(n_15128)
);

OAI22xp5_ASAP7_75t_L g15129 ( 
.A1(n_14552),
.A2(n_13903),
.B1(n_13980),
.B2(n_14348),
.Y(n_15129)
);

AOI22xp33_ASAP7_75t_L g15130 ( 
.A1(n_14278),
.A2(n_1605),
.B1(n_1603),
.B2(n_1604),
.Y(n_15130)
);

OAI21x1_ASAP7_75t_L g15131 ( 
.A1(n_14279),
.A2(n_1604),
.B(n_1605),
.Y(n_15131)
);

NAND3xp33_ASAP7_75t_L g15132 ( 
.A(n_14808),
.B(n_14717),
.C(n_14714),
.Y(n_15132)
);

OAI21x1_ASAP7_75t_L g15133 ( 
.A1(n_14788),
.A2(n_1606),
.B(n_1607),
.Y(n_15133)
);

INVx1_ASAP7_75t_L g15134 ( 
.A(n_13993),
.Y(n_15134)
);

AOI21xp5_ASAP7_75t_L g15135 ( 
.A1(n_14429),
.A2(n_5946),
.B(n_5945),
.Y(n_15135)
);

AO31x2_ASAP7_75t_L g15136 ( 
.A1(n_14558),
.A2(n_1608),
.A3(n_1606),
.B(n_1607),
.Y(n_15136)
);

O2A1O1Ixp5_ASAP7_75t_L g15137 ( 
.A1(n_14646),
.A2(n_14669),
.B(n_14575),
.C(n_14769),
.Y(n_15137)
);

AOI21xp5_ASAP7_75t_L g15138 ( 
.A1(n_14820),
.A2(n_5948),
.B(n_5947),
.Y(n_15138)
);

NOR2xp67_ASAP7_75t_SL g15139 ( 
.A(n_14778),
.B(n_1608),
.Y(n_15139)
);

AOI21xp5_ASAP7_75t_L g15140 ( 
.A1(n_14824),
.A2(n_5951),
.B(n_5950),
.Y(n_15140)
);

CKINVDCx8_ASAP7_75t_R g15141 ( 
.A(n_14115),
.Y(n_15141)
);

OA21x2_ASAP7_75t_L g15142 ( 
.A1(n_14181),
.A2(n_1609),
.B(n_1610),
.Y(n_15142)
);

BUFx6f_ASAP7_75t_L g15143 ( 
.A(n_13960),
.Y(n_15143)
);

INVx1_ASAP7_75t_L g15144 ( 
.A(n_13994),
.Y(n_15144)
);

BUFx6f_ASAP7_75t_L g15145 ( 
.A(n_13971),
.Y(n_15145)
);

INVx1_ASAP7_75t_L g15146 ( 
.A(n_14004),
.Y(n_15146)
);

CKINVDCx16_ASAP7_75t_R g15147 ( 
.A(n_14010),
.Y(n_15147)
);

AOI21xp5_ASAP7_75t_L g15148 ( 
.A1(n_14721),
.A2(n_14739),
.B(n_14492),
.Y(n_15148)
);

BUFx10_ASAP7_75t_L g15149 ( 
.A(n_14017),
.Y(n_15149)
);

OAI21x1_ASAP7_75t_L g15150 ( 
.A1(n_14838),
.A2(n_1609),
.B(n_1611),
.Y(n_15150)
);

AO31x2_ASAP7_75t_L g15151 ( 
.A1(n_14701),
.A2(n_1615),
.A3(n_1612),
.B(n_1614),
.Y(n_15151)
);

AOI221x1_ASAP7_75t_L g15152 ( 
.A1(n_14779),
.A2(n_1615),
.B1(n_1612),
.B2(n_1614),
.C(n_1616),
.Y(n_15152)
);

INVxp67_ASAP7_75t_SL g15153 ( 
.A(n_14142),
.Y(n_15153)
);

NAND2xp5_ASAP7_75t_L g15154 ( 
.A(n_14227),
.B(n_1616),
.Y(n_15154)
);

O2A1O1Ixp33_ASAP7_75t_SL g15155 ( 
.A1(n_14469),
.A2(n_1619),
.B(n_1617),
.C(n_1618),
.Y(n_15155)
);

A2O1A1Ixp33_ASAP7_75t_L g15156 ( 
.A1(n_14032),
.A2(n_14805),
.B(n_14821),
.C(n_14174),
.Y(n_15156)
);

OAI21x1_ASAP7_75t_L g15157 ( 
.A1(n_14842),
.A2(n_1617),
.B(n_1618),
.Y(n_15157)
);

AND2x2_ASAP7_75t_L g15158 ( 
.A(n_14039),
.B(n_1620),
.Y(n_15158)
);

BUFx3_ASAP7_75t_L g15159 ( 
.A(n_14225),
.Y(n_15159)
);

AO31x2_ASAP7_75t_L g15160 ( 
.A1(n_14563),
.A2(n_1623),
.A3(n_1621),
.B(n_1622),
.Y(n_15160)
);

AO31x2_ASAP7_75t_L g15161 ( 
.A1(n_14571),
.A2(n_1623),
.A3(n_1621),
.B(n_1622),
.Y(n_15161)
);

AOI221x1_ASAP7_75t_L g15162 ( 
.A1(n_14373),
.A2(n_1626),
.B1(n_1624),
.B2(n_1625),
.C(n_1627),
.Y(n_15162)
);

OAI21x1_ASAP7_75t_L g15163 ( 
.A1(n_14841),
.A2(n_1625),
.B(n_1626),
.Y(n_15163)
);

INVx1_ASAP7_75t_L g15164 ( 
.A(n_14020),
.Y(n_15164)
);

AOI21xp5_ASAP7_75t_L g15165 ( 
.A1(n_14844),
.A2(n_5953),
.B(n_5952),
.Y(n_15165)
);

AOI221xp5_ASAP7_75t_SL g15166 ( 
.A1(n_14636),
.A2(n_1630),
.B1(n_1628),
.B2(n_1629),
.C(n_1631),
.Y(n_15166)
);

AOI21x1_ASAP7_75t_L g15167 ( 
.A1(n_13973),
.A2(n_1628),
.B(n_1629),
.Y(n_15167)
);

AOI221x1_ASAP7_75t_L g15168 ( 
.A1(n_14235),
.A2(n_1633),
.B1(n_1631),
.B2(n_1632),
.C(n_1634),
.Y(n_15168)
);

NOR2x1_ASAP7_75t_L g15169 ( 
.A(n_14380),
.B(n_1632),
.Y(n_15169)
);

A2O1A1Ixp33_ASAP7_75t_L g15170 ( 
.A1(n_13945),
.A2(n_1635),
.B(n_1633),
.C(n_1634),
.Y(n_15170)
);

AND2x4_ASAP7_75t_L g15171 ( 
.A(n_14315),
.B(n_1635),
.Y(n_15171)
);

NOR2xp67_ASAP7_75t_L g15172 ( 
.A(n_14045),
.B(n_1636),
.Y(n_15172)
);

INVx2_ASAP7_75t_L g15173 ( 
.A(n_14027),
.Y(n_15173)
);

AOI21xp5_ASAP7_75t_L g15174 ( 
.A1(n_14847),
.A2(n_14855),
.B(n_14848),
.Y(n_15174)
);

AO22x2_ASAP7_75t_L g15175 ( 
.A1(n_14046),
.A2(n_1638),
.B1(n_1636),
.B2(n_1637),
.Y(n_15175)
);

OAI21xp5_ASAP7_75t_L g15176 ( 
.A1(n_14776),
.A2(n_1639),
.B(n_1640),
.Y(n_15176)
);

A2O1A1Ixp33_ASAP7_75t_L g15177 ( 
.A1(n_13999),
.A2(n_1641),
.B(n_1639),
.C(n_1640),
.Y(n_15177)
);

OAI21x1_ASAP7_75t_L g15178 ( 
.A1(n_14861),
.A2(n_1642),
.B(n_1643),
.Y(n_15178)
);

OAI21x1_ASAP7_75t_L g15179 ( 
.A1(n_14843),
.A2(n_1642),
.B(n_1643),
.Y(n_15179)
);

BUFx3_ASAP7_75t_L g15180 ( 
.A(n_14225),
.Y(n_15180)
);

O2A1O1Ixp33_ASAP7_75t_L g15181 ( 
.A1(n_14795),
.A2(n_1646),
.B(n_1644),
.C(n_1645),
.Y(n_15181)
);

A2O1A1Ixp33_ASAP7_75t_L g15182 ( 
.A1(n_14690),
.A2(n_14606),
.B(n_14601),
.C(n_14726),
.Y(n_15182)
);

NAND2x1p5_ASAP7_75t_L g15183 ( 
.A(n_14462),
.B(n_5955),
.Y(n_15183)
);

NAND2xp5_ASAP7_75t_L g15184 ( 
.A(n_14240),
.B(n_1644),
.Y(n_15184)
);

INVx2_ASAP7_75t_L g15185 ( 
.A(n_14040),
.Y(n_15185)
);

BUFx6f_ASAP7_75t_L g15186 ( 
.A(n_13971),
.Y(n_15186)
);

O2A1O1Ixp33_ASAP7_75t_L g15187 ( 
.A1(n_14753),
.A2(n_1647),
.B(n_1645),
.C(n_1646),
.Y(n_15187)
);

NAND2xp5_ASAP7_75t_L g15188 ( 
.A(n_14242),
.B(n_1648),
.Y(n_15188)
);

AO32x2_ASAP7_75t_L g15189 ( 
.A1(n_14090),
.A2(n_1650),
.A3(n_1648),
.B1(n_1649),
.B2(n_1651),
.Y(n_15189)
);

OAI21x1_ASAP7_75t_L g15190 ( 
.A1(n_14850),
.A2(n_1649),
.B(n_1650),
.Y(n_15190)
);

AOI21xp5_ASAP7_75t_L g15191 ( 
.A1(n_14570),
.A2(n_5957),
.B(n_5956),
.Y(n_15191)
);

NAND2xp5_ASAP7_75t_L g15192 ( 
.A(n_14244),
.B(n_1651),
.Y(n_15192)
);

AOI21xp5_ASAP7_75t_L g15193 ( 
.A1(n_14829),
.A2(n_5959),
.B(n_5958),
.Y(n_15193)
);

OAI21xp5_ASAP7_75t_L g15194 ( 
.A1(n_14826),
.A2(n_1652),
.B(n_1653),
.Y(n_15194)
);

AOI21xp5_ASAP7_75t_L g15195 ( 
.A1(n_14831),
.A2(n_5961),
.B(n_5960),
.Y(n_15195)
);

INVx3_ASAP7_75t_L g15196 ( 
.A(n_14283),
.Y(n_15196)
);

INVx3_ASAP7_75t_SL g15197 ( 
.A(n_14019),
.Y(n_15197)
);

AOI21xp5_ASAP7_75t_L g15198 ( 
.A1(n_14835),
.A2(n_14856),
.B(n_14506),
.Y(n_15198)
);

NAND2xp5_ASAP7_75t_L g15199 ( 
.A(n_14246),
.B(n_1652),
.Y(n_15199)
);

BUFx6f_ASAP7_75t_L g15200 ( 
.A(n_13983),
.Y(n_15200)
);

OA21x2_ASAP7_75t_L g15201 ( 
.A1(n_14051),
.A2(n_1654),
.B(n_1655),
.Y(n_15201)
);

OAI21xp5_ASAP7_75t_L g15202 ( 
.A1(n_14670),
.A2(n_1654),
.B(n_1655),
.Y(n_15202)
);

HB1xp67_ASAP7_75t_L g15203 ( 
.A(n_14041),
.Y(n_15203)
);

INVx2_ASAP7_75t_SL g15204 ( 
.A(n_14170),
.Y(n_15204)
);

OA21x2_ASAP7_75t_L g15205 ( 
.A1(n_14006),
.A2(n_1656),
.B(n_1657),
.Y(n_15205)
);

OAI21x1_ASAP7_75t_L g15206 ( 
.A1(n_14854),
.A2(n_1656),
.B(n_1658),
.Y(n_15206)
);

OAI22x1_ASAP7_75t_L g15207 ( 
.A1(n_14194),
.A2(n_1660),
.B1(n_1658),
.B2(n_1659),
.Y(n_15207)
);

OAI21xp5_ASAP7_75t_L g15208 ( 
.A1(n_14266),
.A2(n_1659),
.B(n_1661),
.Y(n_15208)
);

INVx3_ASAP7_75t_L g15209 ( 
.A(n_14169),
.Y(n_15209)
);

NAND2xp33_ASAP7_75t_L g15210 ( 
.A(n_14214),
.B(n_1661),
.Y(n_15210)
);

AO21x1_ASAP7_75t_L g15211 ( 
.A1(n_14368),
.A2(n_1662),
.B(n_1663),
.Y(n_15211)
);

A2O1A1Ixp33_ASAP7_75t_L g15212 ( 
.A1(n_14737),
.A2(n_1664),
.B(n_1662),
.C(n_1663),
.Y(n_15212)
);

A2O1A1Ixp33_ASAP7_75t_L g15213 ( 
.A1(n_14671),
.A2(n_1666),
.B(n_1664),
.C(n_1665),
.Y(n_15213)
);

NAND2xp5_ASAP7_75t_L g15214 ( 
.A(n_14247),
.B(n_1665),
.Y(n_15214)
);

AOI21xp5_ASAP7_75t_L g15215 ( 
.A1(n_14527),
.A2(n_5963),
.B(n_5962),
.Y(n_15215)
);

CKINVDCx8_ASAP7_75t_R g15216 ( 
.A(n_14350),
.Y(n_15216)
);

NAND3xp33_ASAP7_75t_SL g15217 ( 
.A(n_14335),
.B(n_1666),
.C(n_1667),
.Y(n_15217)
);

OR2x2_ASAP7_75t_L g15218 ( 
.A(n_14057),
.B(n_14059),
.Y(n_15218)
);

AOI221x1_ASAP7_75t_L g15219 ( 
.A1(n_14249),
.A2(n_1669),
.B1(n_1667),
.B2(n_1668),
.C(n_1670),
.Y(n_15219)
);

INVx1_ASAP7_75t_L g15220 ( 
.A(n_14102),
.Y(n_15220)
);

AO31x2_ASAP7_75t_L g15221 ( 
.A1(n_14459),
.A2(n_1671),
.A3(n_1668),
.B(n_1670),
.Y(n_15221)
);

AOI22xp33_ASAP7_75t_L g15222 ( 
.A1(n_14453),
.A2(n_14822),
.B1(n_14661),
.B2(n_14767),
.Y(n_15222)
);

INVx2_ASAP7_75t_L g15223 ( 
.A(n_14093),
.Y(n_15223)
);

OAI21xp5_ASAP7_75t_L g15224 ( 
.A1(n_14309),
.A2(n_1671),
.B(n_1672),
.Y(n_15224)
);

NAND2xp5_ASAP7_75t_L g15225 ( 
.A(n_14256),
.B(n_1672),
.Y(n_15225)
);

OAI21xp5_ASAP7_75t_L g15226 ( 
.A1(n_14665),
.A2(n_1673),
.B(n_1674),
.Y(n_15226)
);

AOI21xp5_ASAP7_75t_L g15227 ( 
.A1(n_14491),
.A2(n_5967),
.B(n_5966),
.Y(n_15227)
);

AOI21xp5_ASAP7_75t_L g15228 ( 
.A1(n_14538),
.A2(n_5970),
.B(n_5969),
.Y(n_15228)
);

INVx3_ASAP7_75t_L g15229 ( 
.A(n_14251),
.Y(n_15229)
);

AO31x2_ASAP7_75t_L g15230 ( 
.A1(n_14263),
.A2(n_1675),
.A3(n_1673),
.B(n_1674),
.Y(n_15230)
);

BUFx2_ASAP7_75t_SL g15231 ( 
.A(n_14033),
.Y(n_15231)
);

INVx1_ASAP7_75t_L g15232 ( 
.A(n_14104),
.Y(n_15232)
);

INVx2_ASAP7_75t_L g15233 ( 
.A(n_14118),
.Y(n_15233)
);

AND2x2_ASAP7_75t_L g15234 ( 
.A(n_14179),
.B(n_1675),
.Y(n_15234)
);

INVx2_ASAP7_75t_L g15235 ( 
.A(n_14121),
.Y(n_15235)
);

NOR2xp67_ASAP7_75t_SL g15236 ( 
.A(n_14796),
.B(n_1676),
.Y(n_15236)
);

O2A1O1Ixp33_ASAP7_75t_L g15237 ( 
.A1(n_14698),
.A2(n_1678),
.B(n_1676),
.C(n_1677),
.Y(n_15237)
);

BUFx2_ASAP7_75t_L g15238 ( 
.A(n_14195),
.Y(n_15238)
);

NOR2x1_ASAP7_75t_L g15239 ( 
.A(n_14378),
.B(n_1677),
.Y(n_15239)
);

OAI21xp5_ASAP7_75t_L g15240 ( 
.A1(n_14360),
.A2(n_1678),
.B(n_1679),
.Y(n_15240)
);

INVx2_ASAP7_75t_L g15241 ( 
.A(n_14111),
.Y(n_15241)
);

AOI21xp5_ASAP7_75t_L g15242 ( 
.A1(n_14857),
.A2(n_5973),
.B(n_5971),
.Y(n_15242)
);

NOR2x1_ASAP7_75t_SL g15243 ( 
.A(n_14132),
.B(n_1679),
.Y(n_15243)
);

AOI21xp5_ASAP7_75t_L g15244 ( 
.A1(n_14859),
.A2(n_5975),
.B(n_5974),
.Y(n_15244)
);

AOI21x1_ASAP7_75t_L g15245 ( 
.A1(n_13931),
.A2(n_1680),
.B(n_1681),
.Y(n_15245)
);

BUFx2_ASAP7_75t_L g15246 ( 
.A(n_14208),
.Y(n_15246)
);

NAND2xp5_ASAP7_75t_L g15247 ( 
.A(n_14268),
.B(n_1680),
.Y(n_15247)
);

NOR2xp33_ASAP7_75t_L g15248 ( 
.A(n_14568),
.B(n_14581),
.Y(n_15248)
);

AO32x2_ASAP7_75t_L g15249 ( 
.A1(n_14756),
.A2(n_1683),
.A3(n_1681),
.B1(n_1682),
.B2(n_1684),
.Y(n_15249)
);

AOI21xp5_ASAP7_75t_L g15250 ( 
.A1(n_14651),
.A2(n_5978),
.B(n_5976),
.Y(n_15250)
);

INVx3_ASAP7_75t_L g15251 ( 
.A(n_13972),
.Y(n_15251)
);

AO31x2_ASAP7_75t_L g15252 ( 
.A1(n_14272),
.A2(n_1684),
.A3(n_1682),
.B(n_1683),
.Y(n_15252)
);

OAI21x1_ASAP7_75t_L g15253 ( 
.A1(n_14647),
.A2(n_1685),
.B(n_1686),
.Y(n_15253)
);

AOI21xp5_ASAP7_75t_L g15254 ( 
.A1(n_14343),
.A2(n_5980),
.B(n_5979),
.Y(n_15254)
);

NOR2x1_ASAP7_75t_R g15255 ( 
.A(n_14171),
.B(n_1685),
.Y(n_15255)
);

INVx5_ASAP7_75t_L g15256 ( 
.A(n_14214),
.Y(n_15256)
);

NAND2xp5_ASAP7_75t_L g15257 ( 
.A(n_14286),
.B(n_1686),
.Y(n_15257)
);

OAI22xp5_ASAP7_75t_L g15258 ( 
.A1(n_13963),
.A2(n_1689),
.B1(n_1687),
.B2(n_1688),
.Y(n_15258)
);

NAND4xp25_ASAP7_75t_L g15259 ( 
.A(n_14634),
.B(n_1689),
.C(n_1687),
.D(n_1688),
.Y(n_15259)
);

A2O1A1Ixp33_ASAP7_75t_L g15260 ( 
.A1(n_14680),
.A2(n_1692),
.B(n_1690),
.C(n_1691),
.Y(n_15260)
);

O2A1O1Ixp5_ASAP7_75t_L g15261 ( 
.A1(n_14691),
.A2(n_1693),
.B(n_1691),
.C(n_1692),
.Y(n_15261)
);

NOR2xp33_ASAP7_75t_L g15262 ( 
.A(n_14215),
.B(n_1693),
.Y(n_15262)
);

AOI21xp5_ASAP7_75t_L g15263 ( 
.A1(n_14675),
.A2(n_5982),
.B(n_5981),
.Y(n_15263)
);

AND2x2_ASAP7_75t_L g15264 ( 
.A(n_14407),
.B(n_14289),
.Y(n_15264)
);

BUFx10_ASAP7_75t_L g15265 ( 
.A(n_14237),
.Y(n_15265)
);

NAND2xp5_ASAP7_75t_L g15266 ( 
.A(n_14294),
.B(n_1694),
.Y(n_15266)
);

AOI21xp5_ASAP7_75t_L g15267 ( 
.A1(n_14524),
.A2(n_5985),
.B(n_5983),
.Y(n_15267)
);

INVx2_ASAP7_75t_L g15268 ( 
.A(n_14114),
.Y(n_15268)
);

NAND2xp5_ASAP7_75t_L g15269 ( 
.A(n_14310),
.B(n_1695),
.Y(n_15269)
);

INVx1_ASAP7_75t_L g15270 ( 
.A(n_14117),
.Y(n_15270)
);

OAI21x1_ASAP7_75t_SL g15271 ( 
.A1(n_14488),
.A2(n_1695),
.B(n_1696),
.Y(n_15271)
);

AO31x2_ASAP7_75t_L g15272 ( 
.A1(n_14312),
.A2(n_1698),
.A3(n_1696),
.B(n_1697),
.Y(n_15272)
);

NAND2xp5_ASAP7_75t_L g15273 ( 
.A(n_14319),
.B(n_1697),
.Y(n_15273)
);

O2A1O1Ixp33_ASAP7_75t_L g15274 ( 
.A1(n_14707),
.A2(n_1701),
.B(n_1699),
.C(n_1700),
.Y(n_15274)
);

INVx1_ASAP7_75t_L g15275 ( 
.A(n_14330),
.Y(n_15275)
);

NOR2xp33_ASAP7_75t_L g15276 ( 
.A(n_14282),
.B(n_1699),
.Y(n_15276)
);

OAI21xp5_ASAP7_75t_L g15277 ( 
.A1(n_14189),
.A2(n_1700),
.B(n_1701),
.Y(n_15277)
);

AOI21xp5_ASAP7_75t_L g15278 ( 
.A1(n_14735),
.A2(n_5989),
.B(n_5987),
.Y(n_15278)
);

OAI21xp5_ASAP7_75t_L g15279 ( 
.A1(n_14678),
.A2(n_1702),
.B(n_1703),
.Y(n_15279)
);

OAI21xp5_ASAP7_75t_L g15280 ( 
.A1(n_14693),
.A2(n_1702),
.B(n_1703),
.Y(n_15280)
);

INVx1_ASAP7_75t_L g15281 ( 
.A(n_14344),
.Y(n_15281)
);

INVx2_ASAP7_75t_L g15282 ( 
.A(n_14228),
.Y(n_15282)
);

AOI21xp5_ASAP7_75t_L g15283 ( 
.A1(n_14754),
.A2(n_14807),
.B(n_14658),
.Y(n_15283)
);

OAI21x1_ASAP7_75t_L g15284 ( 
.A1(n_14702),
.A2(n_1704),
.B(n_1705),
.Y(n_15284)
);

AOI21xp5_ASAP7_75t_L g15285 ( 
.A1(n_14381),
.A2(n_5991),
.B(n_5990),
.Y(n_15285)
);

OAI22x1_ASAP7_75t_L g15286 ( 
.A1(n_14369),
.A2(n_1706),
.B1(n_1704),
.B2(n_1705),
.Y(n_15286)
);

AOI221x1_ASAP7_75t_L g15287 ( 
.A1(n_14345),
.A2(n_1708),
.B1(n_1706),
.B2(n_1707),
.C(n_1709),
.Y(n_15287)
);

INVx2_ASAP7_75t_L g15288 ( 
.A(n_14233),
.Y(n_15288)
);

AO31x2_ASAP7_75t_L g15289 ( 
.A1(n_14349),
.A2(n_1711),
.A3(n_1709),
.B(n_1710),
.Y(n_15289)
);

AOI21xp5_ASAP7_75t_L g15290 ( 
.A1(n_14708),
.A2(n_5993),
.B(n_5992),
.Y(n_15290)
);

AO31x2_ASAP7_75t_L g15291 ( 
.A1(n_14357),
.A2(n_14363),
.A3(n_14625),
.B(n_14618),
.Y(n_15291)
);

AOI21xp5_ASAP7_75t_L g15292 ( 
.A1(n_14783),
.A2(n_5995),
.B(n_5994),
.Y(n_15292)
);

INVx2_ASAP7_75t_L g15293 ( 
.A(n_14239),
.Y(n_15293)
);

OAI21x1_ASAP7_75t_L g15294 ( 
.A1(n_14685),
.A2(n_1711),
.B(n_1712),
.Y(n_15294)
);

INVx1_ASAP7_75t_L g15295 ( 
.A(n_14198),
.Y(n_15295)
);

AOI221xp5_ASAP7_75t_SL g15296 ( 
.A1(n_13952),
.A2(n_1714),
.B1(n_1712),
.B2(n_1713),
.C(n_1715),
.Y(n_15296)
);

AOI21xp5_ASAP7_75t_L g15297 ( 
.A1(n_14766),
.A2(n_5997),
.B(n_5996),
.Y(n_15297)
);

AO21x2_ASAP7_75t_L g15298 ( 
.A1(n_13918),
.A2(n_1713),
.B(n_1714),
.Y(n_15298)
);

BUFx2_ASAP7_75t_L g15299 ( 
.A(n_14262),
.Y(n_15299)
);

NAND2xp5_ASAP7_75t_L g15300 ( 
.A(n_14399),
.B(n_1715),
.Y(n_15300)
);

AOI21x1_ASAP7_75t_L g15301 ( 
.A1(n_13936),
.A2(n_1716),
.B(n_1717),
.Y(n_15301)
);

OAI22x1_ASAP7_75t_L g15302 ( 
.A1(n_14410),
.A2(n_1718),
.B1(n_1716),
.B2(n_1717),
.Y(n_15302)
);

A2O1A1Ixp33_ASAP7_75t_L g15303 ( 
.A1(n_14392),
.A2(n_1721),
.B(n_1719),
.C(n_1720),
.Y(n_15303)
);

A2O1A1Ixp33_ASAP7_75t_L g15304 ( 
.A1(n_14456),
.A2(n_1721),
.B(n_1719),
.C(n_1720),
.Y(n_15304)
);

OAI22xp5_ASAP7_75t_L g15305 ( 
.A1(n_14340),
.A2(n_1724),
.B1(n_1722),
.B2(n_1723),
.Y(n_15305)
);

INVx1_ASAP7_75t_L g15306 ( 
.A(n_14202),
.Y(n_15306)
);

AND2x4_ASAP7_75t_L g15307 ( 
.A(n_14267),
.B(n_1723),
.Y(n_15307)
);

A2O1A1Ixp33_ASAP7_75t_L g15308 ( 
.A1(n_14460),
.A2(n_1726),
.B(n_1724),
.C(n_1725),
.Y(n_15308)
);

CKINVDCx20_ASAP7_75t_R g15309 ( 
.A(n_14097),
.Y(n_15309)
);

AND2x2_ASAP7_75t_L g15310 ( 
.A(n_14352),
.B(n_1726),
.Y(n_15310)
);

OAI22x1_ASAP7_75t_L g15311 ( 
.A1(n_14212),
.A2(n_1729),
.B1(n_1727),
.B2(n_1728),
.Y(n_15311)
);

NAND2xp5_ASAP7_75t_L g15312 ( 
.A(n_14400),
.B(n_1728),
.Y(n_15312)
);

INVx1_ASAP7_75t_L g15313 ( 
.A(n_14213),
.Y(n_15313)
);

AO31x2_ASAP7_75t_L g15314 ( 
.A1(n_14275),
.A2(n_1731),
.A3(n_1729),
.B(n_1730),
.Y(n_15314)
);

AND2x2_ASAP7_75t_L g15315 ( 
.A(n_14216),
.B(n_1730),
.Y(n_15315)
);

AOI21xp5_ASAP7_75t_L g15316 ( 
.A1(n_13984),
.A2(n_14833),
.B(n_13998),
.Y(n_15316)
);

OAI21xp5_ASAP7_75t_L g15317 ( 
.A1(n_14176),
.A2(n_1732),
.B(n_1733),
.Y(n_15317)
);

OAI21x1_ASAP7_75t_L g15318 ( 
.A1(n_14687),
.A2(n_1732),
.B(n_1733),
.Y(n_15318)
);

OR2x6_ASAP7_75t_L g15319 ( 
.A(n_13905),
.B(n_1734),
.Y(n_15319)
);

OAI22xp5_ASAP7_75t_L g15320 ( 
.A1(n_14748),
.A2(n_1736),
.B1(n_1734),
.B2(n_1735),
.Y(n_15320)
);

INVx2_ASAP7_75t_L g15321 ( 
.A(n_14276),
.Y(n_15321)
);

AND2x4_ASAP7_75t_L g15322 ( 
.A(n_14285),
.B(n_1735),
.Y(n_15322)
);

AOI21xp5_ASAP7_75t_L g15323 ( 
.A1(n_13929),
.A2(n_14060),
.B(n_14009),
.Y(n_15323)
);

INVx3_ASAP7_75t_L g15324 ( 
.A(n_13974),
.Y(n_15324)
);

CKINVDCx11_ASAP7_75t_R g15325 ( 
.A(n_14241),
.Y(n_15325)
);

INVx2_ASAP7_75t_L g15326 ( 
.A(n_14287),
.Y(n_15326)
);

A2O1A1Ixp33_ASAP7_75t_L g15327 ( 
.A1(n_14468),
.A2(n_1738),
.B(n_1736),
.C(n_1737),
.Y(n_15327)
);

INVx2_ASAP7_75t_L g15328 ( 
.A(n_14288),
.Y(n_15328)
);

INVx1_ASAP7_75t_L g15329 ( 
.A(n_14007),
.Y(n_15329)
);

AOI21xp5_ASAP7_75t_L g15330 ( 
.A1(n_14712),
.A2(n_6000),
.B(n_5999),
.Y(n_15330)
);

OA21x2_ASAP7_75t_L g15331 ( 
.A1(n_14025),
.A2(n_1737),
.B(n_1738),
.Y(n_15331)
);

OR2x2_ASAP7_75t_L g15332 ( 
.A(n_14472),
.B(n_1739),
.Y(n_15332)
);

A2O1A1Ixp33_ASAP7_75t_L g15333 ( 
.A1(n_14537),
.A2(n_1741),
.B(n_1739),
.C(n_1740),
.Y(n_15333)
);

NAND2xp5_ASAP7_75t_L g15334 ( 
.A(n_14513),
.B(n_1740),
.Y(n_15334)
);

NAND2x1p5_ASAP7_75t_L g15335 ( 
.A(n_14434),
.B(n_6001),
.Y(n_15335)
);

AO32x2_ASAP7_75t_L g15336 ( 
.A1(n_14155),
.A2(n_14403),
.A3(n_14433),
.B1(n_14419),
.B2(n_14749),
.Y(n_15336)
);

O2A1O1Ixp33_ASAP7_75t_SL g15337 ( 
.A1(n_14370),
.A2(n_1743),
.B(n_1741),
.C(n_1742),
.Y(n_15337)
);

A2O1A1Ixp33_ASAP7_75t_L g15338 ( 
.A1(n_14801),
.A2(n_1745),
.B(n_1743),
.C(n_1744),
.Y(n_15338)
);

AO31x2_ASAP7_75t_L g15339 ( 
.A1(n_14296),
.A2(n_1746),
.A3(n_1744),
.B(n_1745),
.Y(n_15339)
);

INVx8_ASAP7_75t_L g15340 ( 
.A(n_13983),
.Y(n_15340)
);

A2O1A1Ixp33_ASAP7_75t_L g15341 ( 
.A1(n_14803),
.A2(n_1748),
.B(n_1746),
.C(n_1747),
.Y(n_15341)
);

NAND2xp5_ASAP7_75t_L g15342 ( 
.A(n_14579),
.B(n_14580),
.Y(n_15342)
);

AOI21xp5_ASAP7_75t_L g15343 ( 
.A1(n_14853),
.A2(n_14796),
.B(n_14639),
.Y(n_15343)
);

NAND2x1_ASAP7_75t_L g15344 ( 
.A(n_14299),
.B(n_1747),
.Y(n_15344)
);

OA21x2_ASAP7_75t_L g15345 ( 
.A1(n_14036),
.A2(n_1748),
.B(n_1749),
.Y(n_15345)
);

AO31x2_ASAP7_75t_L g15346 ( 
.A1(n_14314),
.A2(n_1751),
.A3(n_1749),
.B(n_1750),
.Y(n_15346)
);

OAI21x1_ASAP7_75t_L g15347 ( 
.A1(n_14692),
.A2(n_1750),
.B(n_1751),
.Y(n_15347)
);

AND2x2_ASAP7_75t_L g15348 ( 
.A(n_14447),
.B(n_1752),
.Y(n_15348)
);

INVx1_ASAP7_75t_L g15349 ( 
.A(n_14042),
.Y(n_15349)
);

O2A1O1Ixp33_ASAP7_75t_SL g15350 ( 
.A1(n_14372),
.A2(n_1754),
.B(n_1752),
.C(n_1753),
.Y(n_15350)
);

INVx2_ASAP7_75t_L g15351 ( 
.A(n_14317),
.Y(n_15351)
);

AOI22xp33_ASAP7_75t_L g15352 ( 
.A1(n_14453),
.A2(n_1755),
.B1(n_1753),
.B2(n_1754),
.Y(n_15352)
);

AOI21xp5_ASAP7_75t_L g15353 ( 
.A1(n_14724),
.A2(n_6003),
.B(n_6002),
.Y(n_15353)
);

OAI21x1_ASAP7_75t_L g15354 ( 
.A1(n_14695),
.A2(n_1755),
.B(n_1756),
.Y(n_15354)
);

OAI21x1_ASAP7_75t_L g15355 ( 
.A1(n_14703),
.A2(n_1757),
.B(n_1758),
.Y(n_15355)
);

AOI21xp5_ASAP7_75t_SL g15356 ( 
.A1(n_14218),
.A2(n_1757),
.B(n_1758),
.Y(n_15356)
);

NAND2xp5_ASAP7_75t_L g15357 ( 
.A(n_14582),
.B(n_1759),
.Y(n_15357)
);

NAND3xp33_ASAP7_75t_L g15358 ( 
.A(n_14088),
.B(n_1759),
.C(n_1760),
.Y(n_15358)
);

INVx3_ASAP7_75t_SL g15359 ( 
.A(n_14146),
.Y(n_15359)
);

NOR2xp67_ASAP7_75t_SL g15360 ( 
.A(n_14561),
.B(n_1760),
.Y(n_15360)
);

CKINVDCx9p33_ASAP7_75t_R g15361 ( 
.A(n_13990),
.Y(n_15361)
);

O2A1O1Ixp33_ASAP7_75t_L g15362 ( 
.A1(n_14812),
.A2(n_1763),
.B(n_1761),
.C(n_1762),
.Y(n_15362)
);

O2A1O1Ixp33_ASAP7_75t_L g15363 ( 
.A1(n_14816),
.A2(n_1763),
.B(n_1761),
.C(n_1762),
.Y(n_15363)
);

OAI22xp5_ASAP7_75t_L g15364 ( 
.A1(n_14621),
.A2(n_1766),
.B1(n_1764),
.B2(n_1765),
.Y(n_15364)
);

OAI21x1_ASAP7_75t_L g15365 ( 
.A1(n_14704),
.A2(n_1765),
.B(n_1766),
.Y(n_15365)
);

INVx1_ASAP7_75t_L g15366 ( 
.A(n_13985),
.Y(n_15366)
);

OAI21x1_ASAP7_75t_L g15367 ( 
.A1(n_14750),
.A2(n_1767),
.B(n_1768),
.Y(n_15367)
);

INVx1_ASAP7_75t_L g15368 ( 
.A(n_14054),
.Y(n_15368)
);

INVx2_ASAP7_75t_L g15369 ( 
.A(n_14481),
.Y(n_15369)
);

NAND2xp5_ASAP7_75t_L g15370 ( 
.A(n_14591),
.B(n_1768),
.Y(n_15370)
);

OAI21x1_ASAP7_75t_L g15371 ( 
.A1(n_14723),
.A2(n_1769),
.B(n_1770),
.Y(n_15371)
);

AOI21xp5_ASAP7_75t_L g15372 ( 
.A1(n_14725),
.A2(n_6005),
.B(n_6004),
.Y(n_15372)
);

A2O1A1Ixp33_ASAP7_75t_L g15373 ( 
.A1(n_14744),
.A2(n_1771),
.B(n_1769),
.C(n_1770),
.Y(n_15373)
);

INVx2_ASAP7_75t_SL g15374 ( 
.A(n_14377),
.Y(n_15374)
);

INVx1_ASAP7_75t_L g15375 ( 
.A(n_14061),
.Y(n_15375)
);

OA21x2_ASAP7_75t_L g15376 ( 
.A1(n_13920),
.A2(n_1771),
.B(n_1772),
.Y(n_15376)
);

AOI21xp5_ASAP7_75t_L g15377 ( 
.A1(n_14727),
.A2(n_6007),
.B(n_6006),
.Y(n_15377)
);

O2A1O1Ixp33_ASAP7_75t_L g15378 ( 
.A1(n_14728),
.A2(n_1774),
.B(n_1772),
.C(n_1773),
.Y(n_15378)
);

INVx1_ASAP7_75t_L g15379 ( 
.A(n_14068),
.Y(n_15379)
);

INVx2_ASAP7_75t_L g15380 ( 
.A(n_14486),
.Y(n_15380)
);

AOI21xp5_ASAP7_75t_L g15381 ( 
.A1(n_14742),
.A2(n_6010),
.B(n_6008),
.Y(n_15381)
);

O2A1O1Ixp33_ASAP7_75t_SL g15382 ( 
.A1(n_14374),
.A2(n_1775),
.B(n_1773),
.C(n_1774),
.Y(n_15382)
);

AOI21xp5_ASAP7_75t_L g15383 ( 
.A1(n_14083),
.A2(n_6012),
.B(n_6011),
.Y(n_15383)
);

AO32x2_ASAP7_75t_L g15384 ( 
.A1(n_14736),
.A2(n_1777),
.A3(n_1775),
.B1(n_1776),
.B2(n_1778),
.Y(n_15384)
);

INVx1_ASAP7_75t_L g15385 ( 
.A(n_14035),
.Y(n_15385)
);

A2O1A1Ixp33_ASAP7_75t_L g15386 ( 
.A1(n_14752),
.A2(n_1779),
.B(n_1776),
.C(n_1778),
.Y(n_15386)
);

A2O1A1Ixp33_ASAP7_75t_L g15387 ( 
.A1(n_14673),
.A2(n_1781),
.B(n_1779),
.C(n_1780),
.Y(n_15387)
);

OAI21x1_ASAP7_75t_L g15388 ( 
.A1(n_14730),
.A2(n_1781),
.B(n_1782),
.Y(n_15388)
);

OAI21x1_ASAP7_75t_L g15389 ( 
.A1(n_14731),
.A2(n_1782),
.B(n_1783),
.Y(n_15389)
);

AO31x2_ASAP7_75t_L g15390 ( 
.A1(n_14627),
.A2(n_14630),
.A3(n_14682),
.B(n_14755),
.Y(n_15390)
);

O2A1O1Ixp33_ASAP7_75t_SL g15391 ( 
.A1(n_14379),
.A2(n_1785),
.B(n_1783),
.C(n_1784),
.Y(n_15391)
);

AOI21xp5_ASAP7_75t_L g15392 ( 
.A1(n_14461),
.A2(n_6014),
.B(n_6013),
.Y(n_15392)
);

OAI22xp5_ASAP7_75t_L g15393 ( 
.A1(n_14631),
.A2(n_1786),
.B1(n_1784),
.B2(n_1785),
.Y(n_15393)
);

BUFx2_ASAP7_75t_L g15394 ( 
.A(n_14140),
.Y(n_15394)
);

NOR2xp67_ASAP7_75t_L g15395 ( 
.A(n_14592),
.B(n_1786),
.Y(n_15395)
);

BUFx10_ASAP7_75t_L g15396 ( 
.A(n_14327),
.Y(n_15396)
);

OAI21xp5_ASAP7_75t_L g15397 ( 
.A1(n_14475),
.A2(n_1787),
.B(n_1788),
.Y(n_15397)
);

AOI21xp5_ASAP7_75t_L g15398 ( 
.A1(n_14740),
.A2(n_6016),
.B(n_6015),
.Y(n_15398)
);

INVx2_ASAP7_75t_L g15399 ( 
.A(n_14500),
.Y(n_15399)
);

AO21x2_ASAP7_75t_L g15400 ( 
.A1(n_13922),
.A2(n_13924),
.B(n_13943),
.Y(n_15400)
);

AOI22xp5_ASAP7_75t_L g15401 ( 
.A1(n_14453),
.A2(n_1790),
.B1(n_1788),
.B2(n_1789),
.Y(n_15401)
);

AND2x2_ASAP7_75t_L g15402 ( 
.A(n_14501),
.B(n_1789),
.Y(n_15402)
);

INVx1_ASAP7_75t_L g15403 ( 
.A(n_14048),
.Y(n_15403)
);

AOI221x1_ASAP7_75t_L g15404 ( 
.A1(n_14594),
.A2(n_1792),
.B1(n_1790),
.B2(n_1791),
.C(n_1793),
.Y(n_15404)
);

AOI21xp5_ASAP7_75t_L g15405 ( 
.A1(n_14777),
.A2(n_6018),
.B(n_6017),
.Y(n_15405)
);

AOI21xp5_ASAP7_75t_L g15406 ( 
.A1(n_14457),
.A2(n_6020),
.B(n_6019),
.Y(n_15406)
);

INVx6_ASAP7_75t_L g15407 ( 
.A(n_13992),
.Y(n_15407)
);

OAI21x1_ASAP7_75t_L g15408 ( 
.A1(n_14733),
.A2(n_1791),
.B(n_1792),
.Y(n_15408)
);

O2A1O1Ixp33_ASAP7_75t_L g15409 ( 
.A1(n_14674),
.A2(n_1795),
.B(n_1793),
.C(n_1794),
.Y(n_15409)
);

OAI21x1_ASAP7_75t_L g15410 ( 
.A1(n_14743),
.A2(n_1794),
.B(n_1795),
.Y(n_15410)
);

BUFx6f_ASAP7_75t_L g15411 ( 
.A(n_13992),
.Y(n_15411)
);

AO32x2_ASAP7_75t_L g15412 ( 
.A1(n_14765),
.A2(n_14050),
.A3(n_14303),
.B1(n_14358),
.B2(n_14105),
.Y(n_15412)
);

NAND2xp5_ASAP7_75t_L g15413 ( 
.A(n_14509),
.B(n_1796),
.Y(n_15413)
);

AO31x2_ASAP7_75t_L g15414 ( 
.A1(n_14781),
.A2(n_1798),
.A3(n_1796),
.B(n_1797),
.Y(n_15414)
);

AO32x2_ASAP7_75t_L g15415 ( 
.A1(n_14613),
.A2(n_1799),
.A3(n_1797),
.B1(n_1798),
.B2(n_1800),
.Y(n_15415)
);

INVx8_ASAP7_75t_L g15416 ( 
.A(n_14037),
.Y(n_15416)
);

OAI21xp5_ASAP7_75t_L g15417 ( 
.A1(n_14637),
.A2(n_1799),
.B(n_1800),
.Y(n_15417)
);

INVxp33_ASAP7_75t_L g15418 ( 
.A(n_14291),
.Y(n_15418)
);

AND2x4_ASAP7_75t_L g15419 ( 
.A(n_14196),
.B(n_1801),
.Y(n_15419)
);

AOI21xp5_ASAP7_75t_L g15420 ( 
.A1(n_14827),
.A2(n_6022),
.B(n_6021),
.Y(n_15420)
);

OAI21x1_ASAP7_75t_L g15421 ( 
.A1(n_14758),
.A2(n_1802),
.B(n_1803),
.Y(n_15421)
);

O2A1O1Ixp33_ASAP7_75t_SL g15422 ( 
.A1(n_14383),
.A2(n_1806),
.B(n_1804),
.C(n_1805),
.Y(n_15422)
);

AO31x2_ASAP7_75t_L g15423 ( 
.A1(n_14799),
.A2(n_1806),
.A3(n_1804),
.B(n_1805),
.Y(n_15423)
);

INVx3_ASAP7_75t_L g15424 ( 
.A(n_14011),
.Y(n_15424)
);

AOI22xp33_ASAP7_75t_SL g15425 ( 
.A1(n_14757),
.A2(n_1809),
.B1(n_1807),
.B2(n_1808),
.Y(n_15425)
);

NAND2xp5_ASAP7_75t_L g15426 ( 
.A(n_14514),
.B(n_1807),
.Y(n_15426)
);

BUFx3_ASAP7_75t_L g15427 ( 
.A(n_14072),
.Y(n_15427)
);

OAI21xp5_ASAP7_75t_L g15428 ( 
.A1(n_14645),
.A2(n_1808),
.B(n_1809),
.Y(n_15428)
);

NOR2xp33_ASAP7_75t_L g15429 ( 
.A(n_14430),
.B(n_1810),
.Y(n_15429)
);

NOR2xp33_ASAP7_75t_SL g15430 ( 
.A(n_13935),
.B(n_1811),
.Y(n_15430)
);

AO31x2_ASAP7_75t_L g15431 ( 
.A1(n_14806),
.A2(n_1814),
.A3(n_1812),
.B(n_1813),
.Y(n_15431)
);

A2O1A1Ixp33_ASAP7_75t_L g15432 ( 
.A1(n_14696),
.A2(n_1815),
.B(n_1813),
.C(n_1814),
.Y(n_15432)
);

BUFx12f_ASAP7_75t_L g15433 ( 
.A(n_14037),
.Y(n_15433)
);

OAI21x1_ASAP7_75t_L g15434 ( 
.A1(n_14672),
.A2(n_1815),
.B(n_1816),
.Y(n_15434)
);

OR2x2_ASAP7_75t_L g15435 ( 
.A(n_14519),
.B(n_14270),
.Y(n_15435)
);

AOI22xp5_ASAP7_75t_L g15436 ( 
.A1(n_14860),
.A2(n_1818),
.B1(n_1816),
.B2(n_1817),
.Y(n_15436)
);

O2A1O1Ixp33_ASAP7_75t_L g15437 ( 
.A1(n_14663),
.A2(n_1819),
.B(n_1817),
.C(n_1818),
.Y(n_15437)
);

INVx2_ASAP7_75t_L g15438 ( 
.A(n_14096),
.Y(n_15438)
);

A2O1A1Ixp33_ASAP7_75t_L g15439 ( 
.A1(n_14722),
.A2(n_14588),
.B(n_14761),
.C(n_14738),
.Y(n_15439)
);

OR2x2_ASAP7_75t_L g15440 ( 
.A(n_14334),
.B(n_1819),
.Y(n_15440)
);

A2O1A1Ixp33_ASAP7_75t_L g15441 ( 
.A1(n_14190),
.A2(n_1822),
.B(n_1820),
.C(n_1821),
.Y(n_15441)
);

NOR2xp33_ASAP7_75t_L g15442 ( 
.A(n_14529),
.B(n_1820),
.Y(n_15442)
);

BUFx2_ASAP7_75t_L g15443 ( 
.A(n_14113),
.Y(n_15443)
);

NAND2xp5_ASAP7_75t_L g15444 ( 
.A(n_14049),
.B(n_1821),
.Y(n_15444)
);

NOR4xp25_ASAP7_75t_L g15445 ( 
.A(n_14638),
.B(n_1824),
.C(n_1822),
.D(n_1823),
.Y(n_15445)
);

INVx4_ASAP7_75t_L g15446 ( 
.A(n_14356),
.Y(n_15446)
);

INVx1_ASAP7_75t_L g15447 ( 
.A(n_13948),
.Y(n_15447)
);

NAND3xp33_ASAP7_75t_L g15448 ( 
.A(n_14689),
.B(n_1824),
.C(n_1825),
.Y(n_15448)
);

OAI21x1_ASAP7_75t_L g15449 ( 
.A1(n_14534),
.A2(n_1825),
.B(n_1826),
.Y(n_15449)
);

NAND2xp5_ASAP7_75t_L g15450 ( 
.A(n_14144),
.B(n_1826),
.Y(n_15450)
);

NAND2xp5_ASAP7_75t_L g15451 ( 
.A(n_13966),
.B(n_1827),
.Y(n_15451)
);

AOI21xp5_ASAP7_75t_L g15452 ( 
.A1(n_14711),
.A2(n_6024),
.B(n_6023),
.Y(n_15452)
);

NOR2xp33_ASAP7_75t_SL g15453 ( 
.A(n_14436),
.B(n_1827),
.Y(n_15453)
);

AO31x2_ASAP7_75t_L g15454 ( 
.A1(n_14770),
.A2(n_1830),
.A3(n_1828),
.B(n_1829),
.Y(n_15454)
);

AOI221x1_ASAP7_75t_L g15455 ( 
.A1(n_13979),
.A2(n_1830),
.B1(n_1828),
.B2(n_1829),
.C(n_1831),
.Y(n_15455)
);

AO31x2_ASAP7_75t_L g15456 ( 
.A1(n_14773),
.A2(n_1833),
.A3(n_1831),
.B(n_1832),
.Y(n_15456)
);

NAND2xp5_ASAP7_75t_L g15457 ( 
.A(n_14596),
.B(n_1833),
.Y(n_15457)
);

INVx2_ASAP7_75t_L g15458 ( 
.A(n_14252),
.Y(n_15458)
);

OR2x2_ASAP7_75t_L g15459 ( 
.A(n_13997),
.B(n_1834),
.Y(n_15459)
);

OAI21x1_ASAP7_75t_L g15460 ( 
.A1(n_13988),
.A2(n_1834),
.B(n_1835),
.Y(n_15460)
);

AOI221xp5_ASAP7_75t_L g15461 ( 
.A1(n_14238),
.A2(n_1838),
.B1(n_1836),
.B2(n_1837),
.C(n_1839),
.Y(n_15461)
);

NAND2xp5_ASAP7_75t_L g15462 ( 
.A(n_13981),
.B(n_13908),
.Y(n_15462)
);

INVx1_ASAP7_75t_L g15463 ( 
.A(n_13991),
.Y(n_15463)
);

AOI21xp5_ASAP7_75t_L g15464 ( 
.A1(n_14793),
.A2(n_14710),
.B(n_14476),
.Y(n_15464)
);

INVx1_ASAP7_75t_L g15465 ( 
.A(n_14080),
.Y(n_15465)
);

BUFx3_ASAP7_75t_L g15466 ( 
.A(n_14131),
.Y(n_15466)
);

AOI21xp5_ASAP7_75t_L g15467 ( 
.A1(n_14371),
.A2(n_6027),
.B(n_6026),
.Y(n_15467)
);

NOR2xp33_ASAP7_75t_L g15468 ( 
.A(n_14607),
.B(n_1836),
.Y(n_15468)
);

BUFx10_ASAP7_75t_L g15469 ( 
.A(n_14220),
.Y(n_15469)
);

OR2x2_ASAP7_75t_L g15470 ( 
.A(n_13926),
.B(n_1837),
.Y(n_15470)
);

OAI21xp5_ASAP7_75t_L g15471 ( 
.A1(n_14328),
.A2(n_1838),
.B(n_1839),
.Y(n_15471)
);

NOR2xp67_ASAP7_75t_L g15472 ( 
.A(n_14180),
.B(n_1840),
.Y(n_15472)
);

INVx1_ASAP7_75t_L g15473 ( 
.A(n_14081),
.Y(n_15473)
);

AOI211x1_ASAP7_75t_L g15474 ( 
.A1(n_14398),
.A2(n_1842),
.B(n_1840),
.C(n_1841),
.Y(n_15474)
);

NOR2xp33_ASAP7_75t_L g15475 ( 
.A(n_14496),
.B(n_1841),
.Y(n_15475)
);

OR2x6_ASAP7_75t_L g15476 ( 
.A(n_14561),
.B(n_1842),
.Y(n_15476)
);

INVx2_ASAP7_75t_L g15477 ( 
.A(n_14305),
.Y(n_15477)
);

INVx4_ASAP7_75t_L g15478 ( 
.A(n_14220),
.Y(n_15478)
);

OA21x2_ASAP7_75t_L g15479 ( 
.A1(n_13930),
.A2(n_1843),
.B(n_1844),
.Y(n_15479)
);

AOI21xp5_ASAP7_75t_L g15480 ( 
.A1(n_14655),
.A2(n_14825),
.B(n_14684),
.Y(n_15480)
);

OAI21x1_ASAP7_75t_L g15481 ( 
.A1(n_14652),
.A2(n_1843),
.B(n_1845),
.Y(n_15481)
);

AOI21xp5_ASAP7_75t_L g15482 ( 
.A1(n_14209),
.A2(n_6030),
.B(n_6028),
.Y(n_15482)
);

OAI21x1_ASAP7_75t_L g15483 ( 
.A1(n_14085),
.A2(n_1845),
.B(n_1846),
.Y(n_15483)
);

INVx2_ASAP7_75t_L g15484 ( 
.A(n_14318),
.Y(n_15484)
);

INVx2_ASAP7_75t_L g15485 ( 
.A(n_14116),
.Y(n_15485)
);

OAI21xp5_ASAP7_75t_L g15486 ( 
.A1(n_14668),
.A2(n_1846),
.B(n_1847),
.Y(n_15486)
);

AO31x2_ASAP7_75t_L g15487 ( 
.A1(n_14075),
.A2(n_1849),
.A3(n_1847),
.B(n_1848),
.Y(n_15487)
);

BUFx2_ASAP7_75t_SL g15488 ( 
.A(n_14053),
.Y(n_15488)
);

INVxp67_ASAP7_75t_SL g15489 ( 
.A(n_14086),
.Y(n_15489)
);

OAI21x1_ASAP7_75t_L g15490 ( 
.A1(n_14100),
.A2(n_14107),
.B(n_14103),
.Y(n_15490)
);

OAI21x1_ASAP7_75t_L g15491 ( 
.A1(n_14108),
.A2(n_1850),
.B(n_1851),
.Y(n_15491)
);

INVx5_ASAP7_75t_L g15492 ( 
.A(n_14201),
.Y(n_15492)
);

AOI221x1_ASAP7_75t_L g15493 ( 
.A1(n_14109),
.A2(n_1852),
.B1(n_1850),
.B2(n_1851),
.C(n_1853),
.Y(n_15493)
);

OR2x2_ASAP7_75t_L g15494 ( 
.A(n_14153),
.B(n_1852),
.Y(n_15494)
);

INVx1_ASAP7_75t_L g15495 ( 
.A(n_14112),
.Y(n_15495)
);

NAND2xp5_ASAP7_75t_L g15496 ( 
.A(n_13909),
.B(n_1854),
.Y(n_15496)
);

BUFx6f_ASAP7_75t_L g15497 ( 
.A(n_14026),
.Y(n_15497)
);

OA21x2_ASAP7_75t_L g15498 ( 
.A1(n_14148),
.A2(n_1854),
.B(n_1855),
.Y(n_15498)
);

OAI21x1_ASAP7_75t_L g15499 ( 
.A1(n_14124),
.A2(n_1855),
.B(n_1856),
.Y(n_15499)
);

CKINVDCx5p33_ASAP7_75t_R g15500 ( 
.A(n_14437),
.Y(n_15500)
);

INVx1_ASAP7_75t_L g15501 ( 
.A(n_14128),
.Y(n_15501)
);

BUFx3_ASAP7_75t_L g15502 ( 
.A(n_14193),
.Y(n_15502)
);

OAI21x1_ASAP7_75t_L g15503 ( 
.A1(n_14082),
.A2(n_1857),
.B(n_1858),
.Y(n_15503)
);

OR2x2_ASAP7_75t_L g15504 ( 
.A(n_14221),
.B(n_14454),
.Y(n_15504)
);

O2A1O1Ixp33_ASAP7_75t_L g15505 ( 
.A1(n_14787),
.A2(n_1860),
.B(n_1858),
.C(n_1859),
.Y(n_15505)
);

INVx2_ASAP7_75t_L g15506 ( 
.A(n_14451),
.Y(n_15506)
);

INVx1_ASAP7_75t_L g15507 ( 
.A(n_14151),
.Y(n_15507)
);

OAI21x1_ASAP7_75t_L g15508 ( 
.A1(n_14077),
.A2(n_1859),
.B(n_1860),
.Y(n_15508)
);

NAND2xp5_ASAP7_75t_L g15509 ( 
.A(n_13910),
.B(n_1861),
.Y(n_15509)
);

AOI21xp5_ASAP7_75t_L g15510 ( 
.A1(n_14709),
.A2(n_6032),
.B(n_6031),
.Y(n_15510)
);

AO21x2_ASAP7_75t_L g15511 ( 
.A1(n_13996),
.A2(n_1861),
.B(n_1862),
.Y(n_15511)
);

OAI22xp5_ASAP7_75t_L g15512 ( 
.A1(n_14662),
.A2(n_1864),
.B1(n_1862),
.B2(n_1863),
.Y(n_15512)
);

INVx1_ASAP7_75t_L g15513 ( 
.A(n_14152),
.Y(n_15513)
);

OAI21xp5_ASAP7_75t_L g15514 ( 
.A1(n_14688),
.A2(n_1863),
.B(n_1864),
.Y(n_15514)
);

INVx1_ASAP7_75t_L g15515 ( 
.A(n_14158),
.Y(n_15515)
);

NAND3xp33_ASAP7_75t_L g15516 ( 
.A(n_14789),
.B(n_1866),
.C(n_1867),
.Y(n_15516)
);

OAI21x1_ASAP7_75t_L g15517 ( 
.A1(n_14138),
.A2(n_1866),
.B(n_1867),
.Y(n_15517)
);

O2A1O1Ixp5_ASAP7_75t_L g15518 ( 
.A1(n_14694),
.A2(n_1870),
.B(n_1868),
.C(n_1869),
.Y(n_15518)
);

O2A1O1Ixp33_ASAP7_75t_SL g15519 ( 
.A1(n_14402),
.A2(n_1870),
.B(n_1868),
.C(n_1869),
.Y(n_15519)
);

NAND2xp5_ASAP7_75t_L g15520 ( 
.A(n_13932),
.B(n_1871),
.Y(n_15520)
);

INVx1_ASAP7_75t_L g15521 ( 
.A(n_14159),
.Y(n_15521)
);

OR2x6_ASAP7_75t_L g15522 ( 
.A(n_14612),
.B(n_1871),
.Y(n_15522)
);

OAI22xp5_ASAP7_75t_L g15523 ( 
.A1(n_14633),
.A2(n_1874),
.B1(n_1872),
.B2(n_1873),
.Y(n_15523)
);

OAI22xp5_ASAP7_75t_L g15524 ( 
.A1(n_14421),
.A2(n_1874),
.B1(n_1872),
.B2(n_1873),
.Y(n_15524)
);

INVx1_ASAP7_75t_L g15525 ( 
.A(n_14147),
.Y(n_15525)
);

HB1xp67_ASAP7_75t_L g15526 ( 
.A(n_13939),
.Y(n_15526)
);

INVx1_ASAP7_75t_L g15527 ( 
.A(n_14160),
.Y(n_15527)
);

AO32x2_ASAP7_75t_L g15528 ( 
.A1(n_14785),
.A2(n_1878),
.A3(n_1875),
.B1(n_1876),
.B2(n_1879),
.Y(n_15528)
);

AOI22xp33_ASAP7_75t_L g15529 ( 
.A1(n_14574),
.A2(n_1878),
.B1(n_1875),
.B2(n_1876),
.Y(n_15529)
);

NAND2xp5_ASAP7_75t_SL g15530 ( 
.A(n_14660),
.B(n_1879),
.Y(n_15530)
);

OAI21x1_ASAP7_75t_L g15531 ( 
.A1(n_14642),
.A2(n_14385),
.B(n_14376),
.Y(n_15531)
);

AND2x2_ASAP7_75t_L g15532 ( 
.A(n_14341),
.B(n_1880),
.Y(n_15532)
);

AND2x2_ASAP7_75t_L g15533 ( 
.A(n_14387),
.B(n_14470),
.Y(n_15533)
);

OR2x6_ASAP7_75t_L g15534 ( 
.A(n_14551),
.B(n_1880),
.Y(n_15534)
);

BUFx3_ASAP7_75t_L g15535 ( 
.A(n_14219),
.Y(n_15535)
);

NOR3xp33_ASAP7_75t_L g15536 ( 
.A(n_14590),
.B(n_1881),
.C(n_1882),
.Y(n_15536)
);

AO31x2_ASAP7_75t_L g15537 ( 
.A1(n_14000),
.A2(n_1884),
.A3(n_1882),
.B(n_1883),
.Y(n_15537)
);

INVx2_ASAP7_75t_L g15538 ( 
.A(n_14178),
.Y(n_15538)
);

OAI21x1_ASAP7_75t_L g15539 ( 
.A1(n_14477),
.A2(n_1883),
.B(n_1885),
.Y(n_15539)
);

NAND3xp33_ASAP7_75t_L g15540 ( 
.A(n_14834),
.B(n_1885),
.C(n_1886),
.Y(n_15540)
);

OAI21x1_ASAP7_75t_L g15541 ( 
.A1(n_14763),
.A2(n_1887),
.B(n_1888),
.Y(n_15541)
);

AOI221xp5_ASAP7_75t_SL g15542 ( 
.A1(n_14775),
.A2(n_1889),
.B1(n_1887),
.B2(n_1888),
.C(n_1890),
.Y(n_15542)
);

AOI21xp33_ASAP7_75t_L g15543 ( 
.A1(n_14640),
.A2(n_1889),
.B(n_1890),
.Y(n_15543)
);

BUFx4f_ASAP7_75t_L g15544 ( 
.A(n_14316),
.Y(n_15544)
);

AOI21xp5_ASAP7_75t_L g15545 ( 
.A1(n_14585),
.A2(n_6034),
.B(n_6033),
.Y(n_15545)
);

INVx2_ASAP7_75t_SL g15546 ( 
.A(n_14521),
.Y(n_15546)
);

CKINVDCx20_ASAP7_75t_R g15547 ( 
.A(n_14566),
.Y(n_15547)
);

BUFx3_ASAP7_75t_L g15548 ( 
.A(n_14474),
.Y(n_15548)
);

OAI21x1_ASAP7_75t_L g15549 ( 
.A1(n_14798),
.A2(n_14499),
.B(n_14482),
.Y(n_15549)
);

INVx1_ASAP7_75t_SL g15550 ( 
.A(n_14557),
.Y(n_15550)
);

BUFx3_ASAP7_75t_L g15551 ( 
.A(n_14028),
.Y(n_15551)
);

A2O1A1Ixp33_ASAP7_75t_L g15552 ( 
.A1(n_14715),
.A2(n_1893),
.B(n_1891),
.C(n_1892),
.Y(n_15552)
);

OAI22xp5_ASAP7_75t_L g15553 ( 
.A1(n_14653),
.A2(n_1895),
.B1(n_1891),
.B2(n_1894),
.Y(n_15553)
);

BUFx3_ASAP7_75t_L g15554 ( 
.A(n_14362),
.Y(n_15554)
);

INVx2_ASAP7_75t_SL g15555 ( 
.A(n_13941),
.Y(n_15555)
);

BUFx6f_ASAP7_75t_L g15556 ( 
.A(n_14490),
.Y(n_15556)
);

AOI211x1_ASAP7_75t_L g15557 ( 
.A1(n_14414),
.A2(n_14595),
.B(n_14599),
.C(n_14623),
.Y(n_15557)
);

INVx2_ASAP7_75t_L g15558 ( 
.A(n_13955),
.Y(n_15558)
);

AO31x2_ASAP7_75t_L g15559 ( 
.A1(n_14810),
.A2(n_1896),
.A3(n_1894),
.B(n_1895),
.Y(n_15559)
);

OAI21x1_ASAP7_75t_L g15560 ( 
.A1(n_14657),
.A2(n_1896),
.B(n_1897),
.Y(n_15560)
);

CKINVDCx5p33_ASAP7_75t_R g15561 ( 
.A(n_14463),
.Y(n_15561)
);

BUFx10_ASAP7_75t_L g15562 ( 
.A(n_14123),
.Y(n_15562)
);

AOI21xp33_ASAP7_75t_L g15563 ( 
.A1(n_14666),
.A2(n_1897),
.B(n_1898),
.Y(n_15563)
);

OAI21xp5_ASAP7_75t_L g15564 ( 
.A1(n_14201),
.A2(n_14718),
.B(n_14562),
.Y(n_15564)
);

AO21x2_ASAP7_75t_L g15565 ( 
.A1(n_14071),
.A2(n_1898),
.B(n_1899),
.Y(n_15565)
);

INVx1_ASAP7_75t_L g15566 ( 
.A(n_14034),
.Y(n_15566)
);

A2O1A1Ixp33_ASAP7_75t_L g15567 ( 
.A1(n_14811),
.A2(n_1901),
.B(n_1899),
.C(n_1900),
.Y(n_15567)
);

NOR2xp67_ASAP7_75t_L g15568 ( 
.A(n_14191),
.B(n_1900),
.Y(n_15568)
);

INVx3_ASAP7_75t_L g15569 ( 
.A(n_15446),
.Y(n_15569)
);

INVx6_ASAP7_75t_L g15570 ( 
.A(n_15090),
.Y(n_15570)
);

AND2x6_ASAP7_75t_L g15571 ( 
.A(n_15239),
.B(n_14542),
.Y(n_15571)
);

OA21x2_ASAP7_75t_L g15572 ( 
.A1(n_15031),
.A2(n_14184),
.B(n_14166),
.Y(n_15572)
);

HB1xp67_ASAP7_75t_L g15573 ( 
.A(n_15291),
.Y(n_15573)
);

INVx1_ASAP7_75t_L g15574 ( 
.A(n_14901),
.Y(n_15574)
);

BUFx3_ASAP7_75t_L g15575 ( 
.A(n_15021),
.Y(n_15575)
);

OAI21x1_ASAP7_75t_L g15576 ( 
.A1(n_15174),
.A2(n_14224),
.B(n_14207),
.Y(n_15576)
);

BUFx2_ASAP7_75t_L g15577 ( 
.A(n_14936),
.Y(n_15577)
);

AOI22xp33_ASAP7_75t_L g15578 ( 
.A1(n_14923),
.A2(n_14741),
.B1(n_14794),
.B2(n_14643),
.Y(n_15578)
);

OA21x2_ASAP7_75t_L g15579 ( 
.A1(n_14992),
.A2(n_14164),
.B(n_14226),
.Y(n_15579)
);

HB1xp67_ASAP7_75t_L g15580 ( 
.A(n_15291),
.Y(n_15580)
);

OAI21x1_ASAP7_75t_L g15581 ( 
.A1(n_14963),
.A2(n_14230),
.B(n_14229),
.Y(n_15581)
);

OAI22xp5_ASAP7_75t_L g15582 ( 
.A1(n_15222),
.A2(n_14654),
.B1(n_14683),
.B2(n_14667),
.Y(n_15582)
);

AND2x2_ASAP7_75t_L g15583 ( 
.A(n_15119),
.B(n_14015),
.Y(n_15583)
);

INVx2_ASAP7_75t_L g15584 ( 
.A(n_14882),
.Y(n_15584)
);

NOR2xp33_ASAP7_75t_L g15585 ( 
.A(n_15097),
.B(n_14493),
.Y(n_15585)
);

OR3x4_ASAP7_75t_SL g15586 ( 
.A(n_15024),
.B(n_13947),
.C(n_14644),
.Y(n_15586)
);

INVx1_ASAP7_75t_L g15587 ( 
.A(n_14998),
.Y(n_15587)
);

INVx2_ASAP7_75t_SL g15588 ( 
.A(n_14885),
.Y(n_15588)
);

AND2x2_ASAP7_75t_L g15589 ( 
.A(n_14941),
.B(n_14498),
.Y(n_15589)
);

OAI21x1_ASAP7_75t_L g15590 ( 
.A1(n_14881),
.A2(n_14234),
.B(n_14231),
.Y(n_15590)
);

HB1xp67_ASAP7_75t_L g15591 ( 
.A(n_14872),
.Y(n_15591)
);

NAND2xp5_ASAP7_75t_L g15592 ( 
.A(n_15489),
.B(n_13989),
.Y(n_15592)
);

OAI22xp5_ASAP7_75t_L g15593 ( 
.A1(n_15492),
.A2(n_14760),
.B1(n_14771),
.B2(n_14404),
.Y(n_15593)
);

AOI21xp5_ASAP7_75t_L g15594 ( 
.A1(n_14867),
.A2(n_14895),
.B(n_14878),
.Y(n_15594)
);

OAI21x1_ASAP7_75t_L g15595 ( 
.A1(n_15343),
.A2(n_14248),
.B(n_14243),
.Y(n_15595)
);

BUFx3_ASAP7_75t_L g15596 ( 
.A(n_15044),
.Y(n_15596)
);

CKINVDCx5p33_ASAP7_75t_R g15597 ( 
.A(n_14884),
.Y(n_15597)
);

INVx2_ASAP7_75t_L g15598 ( 
.A(n_14906),
.Y(n_15598)
);

NAND2xp33_ASAP7_75t_L g15599 ( 
.A(n_15124),
.B(n_14201),
.Y(n_15599)
);

OAI21x1_ASAP7_75t_L g15600 ( 
.A1(n_15072),
.A2(n_14870),
.B(n_14868),
.Y(n_15600)
);

NOR2xp33_ASAP7_75t_L g15601 ( 
.A(n_15359),
.B(n_14559),
.Y(n_15601)
);

OAI21x1_ASAP7_75t_L g15602 ( 
.A1(n_15137),
.A2(n_14254),
.B(n_14253),
.Y(n_15602)
);

AO21x2_ASAP7_75t_L g15603 ( 
.A1(n_14932),
.A2(n_14976),
.B(n_14969),
.Y(n_15603)
);

INVx2_ASAP7_75t_L g15604 ( 
.A(n_14999),
.Y(n_15604)
);

OA21x2_ASAP7_75t_L g15605 ( 
.A1(n_14863),
.A2(n_15132),
.B(n_15490),
.Y(n_15605)
);

OAI22x1_ASAP7_75t_L g15606 ( 
.A1(n_14929),
.A2(n_14583),
.B1(n_14602),
.B2(n_14598),
.Y(n_15606)
);

AOI22xp33_ASAP7_75t_L g15607 ( 
.A1(n_14921),
.A2(n_15129),
.B1(n_14910),
.B2(n_14879),
.Y(n_15607)
);

OAI21xp33_ASAP7_75t_L g15608 ( 
.A1(n_14937),
.A2(n_13982),
.B(n_14817),
.Y(n_15608)
);

OAI21x1_ASAP7_75t_L g15609 ( 
.A1(n_14924),
.A2(n_14259),
.B(n_14258),
.Y(n_15609)
);

OA21x2_ASAP7_75t_L g15610 ( 
.A1(n_15342),
.A2(n_14261),
.B(n_14260),
.Y(n_15610)
);

OAI21x1_ASAP7_75t_L g15611 ( 
.A1(n_14913),
.A2(n_14293),
.B(n_14280),
.Y(n_15611)
);

INVx1_ASAP7_75t_L g15612 ( 
.A(n_15008),
.Y(n_15612)
);

INVx1_ASAP7_75t_SL g15613 ( 
.A(n_15023),
.Y(n_15613)
);

INVx1_ASAP7_75t_L g15614 ( 
.A(n_14902),
.Y(n_15614)
);

OAI22xp5_ASAP7_75t_L g15615 ( 
.A1(n_15492),
.A2(n_14697),
.B1(n_14659),
.B2(n_14541),
.Y(n_15615)
);

BUFx2_ASAP7_75t_L g15616 ( 
.A(n_15013),
.Y(n_15616)
);

AND2x2_ASAP7_75t_L g15617 ( 
.A(n_15076),
.B(n_14390),
.Y(n_15617)
);

AO31x2_ASAP7_75t_L g15618 ( 
.A1(n_15211),
.A2(n_14295),
.A3(n_14298),
.B(n_14297),
.Y(n_15618)
);

NAND2x1p5_ASAP7_75t_L g15619 ( 
.A(n_15124),
.B(n_14426),
.Y(n_15619)
);

OAI21x1_ASAP7_75t_L g15620 ( 
.A1(n_15283),
.A2(n_14304),
.B(n_14301),
.Y(n_15620)
);

NAND2x1_ASAP7_75t_L g15621 ( 
.A(n_15126),
.B(n_14091),
.Y(n_15621)
);

INVx1_ASAP7_75t_L g15622 ( 
.A(n_14905),
.Y(n_15622)
);

INVx3_ASAP7_75t_L g15623 ( 
.A(n_15469),
.Y(n_15623)
);

INVx2_ASAP7_75t_L g15624 ( 
.A(n_14959),
.Y(n_15624)
);

INVx5_ASAP7_75t_L g15625 ( 
.A(n_15476),
.Y(n_15625)
);

OR2x2_ASAP7_75t_L g15626 ( 
.A(n_15030),
.B(n_14443),
.Y(n_15626)
);

AOI221xp5_ASAP7_75t_L g15627 ( 
.A1(n_15148),
.A2(n_14611),
.B1(n_14192),
.B2(n_14204),
.C(n_14203),
.Y(n_15627)
);

BUFx3_ASAP7_75t_L g15628 ( 
.A(n_15309),
.Y(n_15628)
);

NOR2xp67_ASAP7_75t_L g15629 ( 
.A(n_15256),
.B(n_14553),
.Y(n_15629)
);

NAND2xp5_ASAP7_75t_L g15630 ( 
.A(n_15153),
.B(n_14333),
.Y(n_15630)
);

AOI21xp5_ASAP7_75t_SL g15631 ( 
.A1(n_14956),
.A2(n_14555),
.B(n_14660),
.Y(n_15631)
);

AOI222xp33_ASAP7_75t_L g15632 ( 
.A1(n_15176),
.A2(n_14706),
.B1(n_14786),
.B2(n_14823),
.C1(n_14185),
.C2(n_14478),
.Y(n_15632)
);

INVx1_ASAP7_75t_L g15633 ( 
.A(n_14916),
.Y(n_15633)
);

INVx3_ASAP7_75t_L g15634 ( 
.A(n_15478),
.Y(n_15634)
);

AO21x2_ASAP7_75t_L g15635 ( 
.A1(n_14954),
.A2(n_14321),
.B(n_14313),
.Y(n_15635)
);

OAI21x1_ASAP7_75t_L g15636 ( 
.A1(n_14874),
.A2(n_14329),
.B(n_14322),
.Y(n_15636)
);

INVx1_ASAP7_75t_L g15637 ( 
.A(n_14939),
.Y(n_15637)
);

OAI21x1_ASAP7_75t_L g15638 ( 
.A1(n_14927),
.A2(n_14331),
.B(n_14206),
.Y(n_15638)
);

AOI22xp33_ASAP7_75t_L g15639 ( 
.A1(n_14889),
.A2(n_14734),
.B1(n_14622),
.B2(n_14584),
.Y(n_15639)
);

NAND2xp5_ASAP7_75t_L g15640 ( 
.A(n_15463),
.B(n_14346),
.Y(n_15640)
);

AND2x2_ASAP7_75t_L g15641 ( 
.A(n_15061),
.B(n_14617),
.Y(n_15641)
);

INVx1_ASAP7_75t_SL g15642 ( 
.A(n_15118),
.Y(n_15642)
);

BUFx6f_ASAP7_75t_L g15643 ( 
.A(n_15497),
.Y(n_15643)
);

OAI21xp5_ASAP7_75t_L g15644 ( 
.A1(n_14940),
.A2(n_14197),
.B(n_14448),
.Y(n_15644)
);

OAI21x1_ASAP7_75t_L g15645 ( 
.A1(n_14919),
.A2(n_14635),
.B(n_14629),
.Y(n_15645)
);

INVx3_ASAP7_75t_L g15646 ( 
.A(n_15548),
.Y(n_15646)
);

NAND2x1p5_ASAP7_75t_L g15647 ( 
.A(n_15256),
.B(n_14471),
.Y(n_15647)
);

NOR2xp33_ASAP7_75t_SL g15648 ( 
.A(n_15141),
.B(n_14523),
.Y(n_15648)
);

OAI21x1_ASAP7_75t_SL g15649 ( 
.A1(n_15243),
.A2(n_14480),
.B(n_14450),
.Y(n_15649)
);

INVx1_ASAP7_75t_L g15650 ( 
.A(n_14946),
.Y(n_15650)
);

OAI21x1_ASAP7_75t_L g15651 ( 
.A1(n_14918),
.A2(n_14746),
.B(n_14489),
.Y(n_15651)
);

INVx2_ASAP7_75t_L g15652 ( 
.A(n_14996),
.Y(n_15652)
);

OAI21xp5_ASAP7_75t_L g15653 ( 
.A1(n_14893),
.A2(n_14504),
.B(n_14484),
.Y(n_15653)
);

INVx1_ASAP7_75t_L g15654 ( 
.A(n_14960),
.Y(n_15654)
);

OAI22xp33_ASAP7_75t_L g15655 ( 
.A1(n_15100),
.A2(n_14734),
.B1(n_14516),
.B2(n_14471),
.Y(n_15655)
);

BUFx2_ASAP7_75t_L g15656 ( 
.A(n_14917),
.Y(n_15656)
);

NAND2x1p5_ASAP7_75t_L g15657 ( 
.A(n_14983),
.B(n_14516),
.Y(n_15657)
);

OAI21x1_ASAP7_75t_L g15658 ( 
.A1(n_14886),
.A2(n_14510),
.B(n_14507),
.Y(n_15658)
);

NAND2xp5_ASAP7_75t_SL g15659 ( 
.A(n_15058),
.B(n_14490),
.Y(n_15659)
);

AND2x2_ASAP7_75t_L g15660 ( 
.A(n_15394),
.B(n_14029),
.Y(n_15660)
);

NOR2xp33_ASAP7_75t_L g15661 ( 
.A(n_15125),
.B(n_14512),
.Y(n_15661)
);

O2A1O1Ixp33_ASAP7_75t_SL g15662 ( 
.A1(n_15439),
.A2(n_14518),
.B(n_14530),
.C(n_14525),
.Y(n_15662)
);

OR2x6_ASAP7_75t_L g15663 ( 
.A(n_15231),
.B(n_14110),
.Y(n_15663)
);

CKINVDCx8_ASAP7_75t_R g15664 ( 
.A(n_15147),
.Y(n_15664)
);

AOI211xp5_ASAP7_75t_L g15665 ( 
.A1(n_15356),
.A2(n_14569),
.B(n_14536),
.C(n_14546),
.Y(n_15665)
);

INVx1_ASAP7_75t_L g15666 ( 
.A(n_14961),
.Y(n_15666)
);

BUFx6f_ASAP7_75t_L g15667 ( 
.A(n_15497),
.Y(n_15667)
);

INVx2_ASAP7_75t_L g15668 ( 
.A(n_15241),
.Y(n_15668)
);

BUFx2_ASAP7_75t_L g15669 ( 
.A(n_14978),
.Y(n_15669)
);

A2O1A1Ixp33_ASAP7_75t_L g15670 ( 
.A1(n_15437),
.A2(n_14587),
.B(n_14605),
.C(n_14576),
.Y(n_15670)
);

INVx1_ASAP7_75t_L g15671 ( 
.A(n_14989),
.Y(n_15671)
);

NOR2x1_ASAP7_75t_SL g15672 ( 
.A(n_15488),
.B(n_14062),
.Y(n_15672)
);

NAND2x1p5_ASAP7_75t_L g15673 ( 
.A(n_15531),
.B(n_14515),
.Y(n_15673)
);

OAI22xp5_ASAP7_75t_L g15674 ( 
.A1(n_15103),
.A2(n_14547),
.B1(n_14567),
.B2(n_14531),
.Y(n_15674)
);

OAI21x1_ASAP7_75t_L g15675 ( 
.A1(n_14942),
.A2(n_14578),
.B(n_14577),
.Y(n_15675)
);

OR2x2_ASAP7_75t_L g15676 ( 
.A(n_15030),
.B(n_14896),
.Y(n_15676)
);

OAI21xp5_ASAP7_75t_L g15677 ( 
.A1(n_14903),
.A2(n_14354),
.B(n_14351),
.Y(n_15677)
);

HB1xp67_ASAP7_75t_L g15678 ( 
.A(n_15390),
.Y(n_15678)
);

AND2x4_ASAP7_75t_L g15679 ( 
.A(n_14966),
.B(n_14332),
.Y(n_15679)
);

OA21x2_ASAP7_75t_L g15680 ( 
.A1(n_15009),
.A2(n_14355),
.B(n_14089),
.Y(n_15680)
);

OA21x2_ASAP7_75t_L g15681 ( 
.A1(n_15027),
.A2(n_15071),
.B(n_15029),
.Y(n_15681)
);

INVx1_ASAP7_75t_L g15682 ( 
.A(n_14993),
.Y(n_15682)
);

BUFx4_ASAP7_75t_R g15683 ( 
.A(n_15058),
.Y(n_15683)
);

BUFx12f_ASAP7_75t_L g15684 ( 
.A(n_15325),
.Y(n_15684)
);

AND2x2_ASAP7_75t_L g15685 ( 
.A(n_15443),
.B(n_14876),
.Y(n_15685)
);

OAI22xp5_ASAP7_75t_L g15686 ( 
.A1(n_15401),
.A2(n_14589),
.B1(n_14751),
.B2(n_14719),
.Y(n_15686)
);

INVx2_ASAP7_75t_L g15687 ( 
.A(n_15268),
.Y(n_15687)
);

INVx3_ASAP7_75t_SL g15688 ( 
.A(n_15561),
.Y(n_15688)
);

AOI21xp5_ASAP7_75t_L g15689 ( 
.A1(n_14911),
.A2(n_14624),
.B(n_14699),
.Y(n_15689)
);

AND2x2_ASAP7_75t_SL g15690 ( 
.A(n_15210),
.B(n_14161),
.Y(n_15690)
);

OAI21x1_ASAP7_75t_L g15691 ( 
.A1(n_15113),
.A2(n_14172),
.B(n_14125),
.Y(n_15691)
);

INVx2_ASAP7_75t_L g15692 ( 
.A(n_15218),
.Y(n_15692)
);

INVx2_ASAP7_75t_L g15693 ( 
.A(n_15032),
.Y(n_15693)
);

CKINVDCx20_ASAP7_75t_R g15694 ( 
.A(n_14875),
.Y(n_15694)
);

AND2x2_ASAP7_75t_L g15695 ( 
.A(n_15112),
.B(n_14183),
.Y(n_15695)
);

NAND2xp5_ASAP7_75t_L g15696 ( 
.A(n_15465),
.B(n_14526),
.Y(n_15696)
);

NAND2xp5_ASAP7_75t_L g15697 ( 
.A(n_15473),
.B(n_14532),
.Y(n_15697)
);

OAI21x1_ASAP7_75t_L g15698 ( 
.A1(n_15056),
.A2(n_14648),
.B(n_14173),
.Y(n_15698)
);

OA21x2_ASAP7_75t_L g15699 ( 
.A1(n_15220),
.A2(n_14375),
.B(n_14364),
.Y(n_15699)
);

O2A1O1Ixp33_ASAP7_75t_L g15700 ( 
.A1(n_15155),
.A2(n_14615),
.B(n_14549),
.C(n_14497),
.Y(n_15700)
);

OAI22xp5_ASAP7_75t_L g15701 ( 
.A1(n_15130),
.A2(n_14628),
.B1(n_14269),
.B2(n_14016),
.Y(n_15701)
);

INVx2_ASAP7_75t_L g15702 ( 
.A(n_15034),
.Y(n_15702)
);

INVx1_ASAP7_75t_L g15703 ( 
.A(n_15232),
.Y(n_15703)
);

NAND2xp5_ASAP7_75t_L g15704 ( 
.A(n_15495),
.B(n_14167),
.Y(n_15704)
);

INVx2_ASAP7_75t_L g15705 ( 
.A(n_14883),
.Y(n_15705)
);

INVx3_ASAP7_75t_L g15706 ( 
.A(n_14930),
.Y(n_15706)
);

BUFx3_ASAP7_75t_L g15707 ( 
.A(n_14984),
.Y(n_15707)
);

INVx1_ASAP7_75t_L g15708 ( 
.A(n_15270),
.Y(n_15708)
);

INVx1_ASAP7_75t_L g15709 ( 
.A(n_15275),
.Y(n_15709)
);

AOI22xp33_ASAP7_75t_SL g15710 ( 
.A1(n_14971),
.A2(n_14520),
.B1(n_14505),
.B2(n_14664),
.Y(n_15710)
);

BUFx12f_ASAP7_75t_L g15711 ( 
.A(n_15265),
.Y(n_15711)
);

AND2x4_ASAP7_75t_L g15712 ( 
.A(n_15204),
.B(n_14290),
.Y(n_15712)
);

OAI21x1_ASAP7_75t_L g15713 ( 
.A1(n_14907),
.A2(n_14119),
.B(n_14320),
.Y(n_15713)
);

OAI21x1_ASAP7_75t_L g15714 ( 
.A1(n_15198),
.A2(n_14306),
.B(n_14386),
.Y(n_15714)
);

NAND3xp33_ASAP7_75t_L g15715 ( 
.A(n_15114),
.B(n_15461),
.C(n_15081),
.Y(n_15715)
);

INVx2_ASAP7_75t_L g15716 ( 
.A(n_14898),
.Y(n_15716)
);

HB1xp67_ASAP7_75t_L g15717 ( 
.A(n_15390),
.Y(n_15717)
);

INVx1_ASAP7_75t_L g15718 ( 
.A(n_15281),
.Y(n_15718)
);

NOR2xp33_ASAP7_75t_SL g15719 ( 
.A(n_15216),
.B(n_14494),
.Y(n_15719)
);

INVx2_ASAP7_75t_L g15720 ( 
.A(n_14944),
.Y(n_15720)
);

AND2x2_ASAP7_75t_L g15721 ( 
.A(n_15264),
.B(n_14222),
.Y(n_15721)
);

OAI22xp33_ASAP7_75t_L g15722 ( 
.A1(n_15022),
.A2(n_14732),
.B1(n_14177),
.B2(n_14211),
.Y(n_15722)
);

NOR2xp33_ASAP7_75t_L g15723 ( 
.A(n_15197),
.B(n_14101),
.Y(n_15723)
);

OAI21x1_ASAP7_75t_L g15724 ( 
.A1(n_15549),
.A2(n_14265),
.B(n_14245),
.Y(n_15724)
);

NAND2xp5_ASAP7_75t_L g15725 ( 
.A(n_15501),
.B(n_15368),
.Y(n_15725)
);

OR2x6_ASAP7_75t_L g15726 ( 
.A(n_14948),
.B(n_14271),
.Y(n_15726)
);

INVx2_ASAP7_75t_L g15727 ( 
.A(n_15246),
.Y(n_15727)
);

AND2x4_ASAP7_75t_L g15728 ( 
.A(n_15438),
.B(n_14273),
.Y(n_15728)
);

AOI21xp5_ASAP7_75t_L g15729 ( 
.A1(n_14912),
.A2(n_14396),
.B(n_14393),
.Y(n_15729)
);

NOR2xp33_ASAP7_75t_L g15730 ( 
.A(n_14988),
.B(n_14413),
.Y(n_15730)
);

INVx3_ASAP7_75t_L g15731 ( 
.A(n_15108),
.Y(n_15731)
);

OAI21xp5_ASAP7_75t_L g15732 ( 
.A1(n_15156),
.A2(n_14432),
.B(n_14431),
.Y(n_15732)
);

INVx1_ASAP7_75t_L g15733 ( 
.A(n_15073),
.Y(n_15733)
);

O2A1O1Ixp33_ASAP7_75t_SL g15734 ( 
.A1(n_15217),
.A2(n_14573),
.B(n_14610),
.C(n_14277),
.Y(n_15734)
);

OA21x2_ASAP7_75t_L g15735 ( 
.A1(n_15078),
.A2(n_14439),
.B(n_14435),
.Y(n_15735)
);

AO21x2_ASAP7_75t_L g15736 ( 
.A1(n_14964),
.A2(n_14483),
.B(n_14466),
.Y(n_15736)
);

INVx1_ASAP7_75t_L g15737 ( 
.A(n_15086),
.Y(n_15737)
);

NAND2xp5_ASAP7_75t_L g15738 ( 
.A(n_15375),
.B(n_14502),
.Y(n_15738)
);

HB1xp67_ASAP7_75t_L g15739 ( 
.A(n_15203),
.Y(n_15739)
);

AO31x2_ASAP7_75t_L g15740 ( 
.A1(n_14922),
.A2(n_14780),
.A3(n_1903),
.B(n_1901),
.Y(n_15740)
);

NAND2xp5_ASAP7_75t_L g15741 ( 
.A(n_15379),
.B(n_1902),
.Y(n_15741)
);

BUFx10_ASAP7_75t_L g15742 ( 
.A(n_14864),
.Y(n_15742)
);

INVx2_ASAP7_75t_L g15743 ( 
.A(n_15299),
.Y(n_15743)
);

NAND2xp5_ASAP7_75t_L g15744 ( 
.A(n_15447),
.B(n_1902),
.Y(n_15744)
);

OAI22xp33_ASAP7_75t_L g15745 ( 
.A1(n_15128),
.A2(n_1905),
.B1(n_1903),
.B2(n_1904),
.Y(n_15745)
);

BUFx3_ASAP7_75t_L g15746 ( 
.A(n_15433),
.Y(n_15746)
);

AO21x2_ASAP7_75t_L g15747 ( 
.A1(n_15172),
.A2(n_1904),
.B(n_1906),
.Y(n_15747)
);

OAI21x1_ASAP7_75t_L g15748 ( 
.A1(n_15069),
.A2(n_1906),
.B(n_1907),
.Y(n_15748)
);

CKINVDCx14_ASAP7_75t_R g15749 ( 
.A(n_15544),
.Y(n_15749)
);

OAI21x1_ASAP7_75t_L g15750 ( 
.A1(n_15088),
.A2(n_1907),
.B(n_1908),
.Y(n_15750)
);

CKINVDCx5p33_ASAP7_75t_R g15751 ( 
.A(n_14951),
.Y(n_15751)
);

OAI22xp33_ASAP7_75t_L g15752 ( 
.A1(n_14871),
.A2(n_1910),
.B1(n_1908),
.B2(n_1909),
.Y(n_15752)
);

AOI22xp33_ASAP7_75t_SL g15753 ( 
.A1(n_15194),
.A2(n_1911),
.B1(n_1909),
.B2(n_1910),
.Y(n_15753)
);

AO21x2_ASAP7_75t_L g15754 ( 
.A1(n_15395),
.A2(n_15017),
.B(n_15033),
.Y(n_15754)
);

INVx1_ASAP7_75t_L g15755 ( 
.A(n_15120),
.Y(n_15755)
);

NAND2xp33_ASAP7_75t_L g15756 ( 
.A(n_15058),
.B(n_1911),
.Y(n_15756)
);

NAND2xp5_ASAP7_75t_L g15757 ( 
.A(n_15507),
.B(n_15513),
.Y(n_15757)
);

OAI21xp33_ASAP7_75t_SL g15758 ( 
.A1(n_15169),
.A2(n_1912),
.B(n_1914),
.Y(n_15758)
);

INVx1_ASAP7_75t_L g15759 ( 
.A(n_15134),
.Y(n_15759)
);

OAI21x1_ASAP7_75t_L g15760 ( 
.A1(n_15157),
.A2(n_1912),
.B(n_1914),
.Y(n_15760)
);

AND2x4_ASAP7_75t_L g15761 ( 
.A(n_15458),
.B(n_1915),
.Y(n_15761)
);

OAI22xp5_ASAP7_75t_L g15762 ( 
.A1(n_15352),
.A2(n_1918),
.B1(n_1916),
.B2(n_1917),
.Y(n_15762)
);

OAI21x1_ASAP7_75t_L g15763 ( 
.A1(n_15163),
.A2(n_1917),
.B(n_1918),
.Y(n_15763)
);

NAND2xp5_ASAP7_75t_L g15764 ( 
.A(n_15515),
.B(n_1919),
.Y(n_15764)
);

OA21x2_ASAP7_75t_L g15765 ( 
.A1(n_15144),
.A2(n_1919),
.B(n_1920),
.Y(n_15765)
);

INVx1_ASAP7_75t_L g15766 ( 
.A(n_15146),
.Y(n_15766)
);

AOI21xp33_ASAP7_75t_SL g15767 ( 
.A1(n_14948),
.A2(n_1920),
.B(n_1921),
.Y(n_15767)
);

AND2x4_ASAP7_75t_L g15768 ( 
.A(n_15477),
.B(n_1922),
.Y(n_15768)
);

OA21x2_ASAP7_75t_L g15769 ( 
.A1(n_15164),
.A2(n_1922),
.B(n_1923),
.Y(n_15769)
);

OAI21x1_ASAP7_75t_L g15770 ( 
.A1(n_15178),
.A2(n_1924),
.B(n_1925),
.Y(n_15770)
);

OAI21x1_ASAP7_75t_L g15771 ( 
.A1(n_14943),
.A2(n_1924),
.B(n_1925),
.Y(n_15771)
);

NOR2xp67_ASAP7_75t_SL g15772 ( 
.A(n_15051),
.B(n_1926),
.Y(n_15772)
);

INVx2_ASAP7_75t_L g15773 ( 
.A(n_15080),
.Y(n_15773)
);

INVx2_ASAP7_75t_L g15774 ( 
.A(n_15082),
.Y(n_15774)
);

AO21x2_ASAP7_75t_L g15775 ( 
.A1(n_15004),
.A2(n_1927),
.B(n_1928),
.Y(n_15775)
);

OR2x6_ASAP7_75t_L g15776 ( 
.A(n_15316),
.B(n_1928),
.Y(n_15776)
);

AOI21xp5_ASAP7_75t_L g15777 ( 
.A1(n_14891),
.A2(n_14915),
.B(n_14866),
.Y(n_15777)
);

OR2x2_ASAP7_75t_L g15778 ( 
.A(n_15435),
.B(n_1929),
.Y(n_15778)
);

INVx1_ASAP7_75t_L g15779 ( 
.A(n_15369),
.Y(n_15779)
);

CKINVDCx20_ASAP7_75t_R g15780 ( 
.A(n_15059),
.Y(n_15780)
);

NOR2xp33_ASAP7_75t_SL g15781 ( 
.A(n_15255),
.B(n_1929),
.Y(n_15781)
);

INVx1_ASAP7_75t_L g15782 ( 
.A(n_15380),
.Y(n_15782)
);

INVx2_ASAP7_75t_L g15783 ( 
.A(n_15091),
.Y(n_15783)
);

AOI21xp5_ASAP7_75t_L g15784 ( 
.A1(n_14934),
.A2(n_14928),
.B(n_14931),
.Y(n_15784)
);

OAI21x1_ASAP7_75t_L g15785 ( 
.A1(n_15133),
.A2(n_1930),
.B(n_1931),
.Y(n_15785)
);

OAI22xp5_ASAP7_75t_SL g15786 ( 
.A1(n_15425),
.A2(n_15557),
.B1(n_15474),
.B2(n_15445),
.Y(n_15786)
);

AO21x2_ASAP7_75t_L g15787 ( 
.A1(n_15300),
.A2(n_1930),
.B(n_1931),
.Y(n_15787)
);

INVx2_ASAP7_75t_L g15788 ( 
.A(n_15092),
.Y(n_15788)
);

OAI21x1_ASAP7_75t_L g15789 ( 
.A1(n_14897),
.A2(n_1932),
.B(n_1933),
.Y(n_15789)
);

NOR2xp67_ASAP7_75t_L g15790 ( 
.A(n_15374),
.B(n_1932),
.Y(n_15790)
);

NAND2xp5_ASAP7_75t_L g15791 ( 
.A(n_15521),
.B(n_1933),
.Y(n_15791)
);

BUFx3_ASAP7_75t_L g15792 ( 
.A(n_14880),
.Y(n_15792)
);

AOI22xp33_ASAP7_75t_L g15793 ( 
.A1(n_14914),
.A2(n_1936),
.B1(n_1934),
.B2(n_1935),
.Y(n_15793)
);

INVx6_ASAP7_75t_L g15794 ( 
.A(n_15396),
.Y(n_15794)
);

OAI22xp5_ASAP7_75t_L g15795 ( 
.A1(n_15358),
.A2(n_1936),
.B1(n_1934),
.B2(n_1935),
.Y(n_15795)
);

OA21x2_ASAP7_75t_L g15796 ( 
.A1(n_15116),
.A2(n_1937),
.B(n_1938),
.Y(n_15796)
);

NAND2x1p5_ASAP7_75t_L g15797 ( 
.A(n_15139),
.B(n_14887),
.Y(n_15797)
);

INVx1_ASAP7_75t_L g15798 ( 
.A(n_15399),
.Y(n_15798)
);

INVx1_ASAP7_75t_L g15799 ( 
.A(n_15295),
.Y(n_15799)
);

NAND2xp5_ASAP7_75t_L g15800 ( 
.A(n_15400),
.B(n_15329),
.Y(n_15800)
);

AOI22xp33_ASAP7_75t_L g15801 ( 
.A1(n_15043),
.A2(n_1939),
.B1(n_1937),
.B2(n_1938),
.Y(n_15801)
);

INVx1_ASAP7_75t_L g15802 ( 
.A(n_15306),
.Y(n_15802)
);

OAI21xp5_ASAP7_75t_L g15803 ( 
.A1(n_14899),
.A2(n_1939),
.B(n_1940),
.Y(n_15803)
);

AOI21xp33_ASAP7_75t_L g15804 ( 
.A1(n_15362),
.A2(n_15363),
.B(n_15409),
.Y(n_15804)
);

CKINVDCx5p33_ASAP7_75t_R g15805 ( 
.A(n_15060),
.Y(n_15805)
);

INVx2_ASAP7_75t_L g15806 ( 
.A(n_15173),
.Y(n_15806)
);

OAI21xp5_ASAP7_75t_L g15807 ( 
.A1(n_15564),
.A2(n_1940),
.B(n_1941),
.Y(n_15807)
);

AOI21x1_ASAP7_75t_L g15808 ( 
.A1(n_15096),
.A2(n_1941),
.B(n_1942),
.Y(n_15808)
);

OAI21x1_ASAP7_75t_L g15809 ( 
.A1(n_15066),
.A2(n_1942),
.B(n_1943),
.Y(n_15809)
);

OAI21x1_ASAP7_75t_L g15810 ( 
.A1(n_15068),
.A2(n_1944),
.B(n_1945),
.Y(n_15810)
);

INVx2_ASAP7_75t_L g15811 ( 
.A(n_15185),
.Y(n_15811)
);

INVxp67_ASAP7_75t_L g15812 ( 
.A(n_15050),
.Y(n_15812)
);

BUFx12f_ASAP7_75t_L g15813 ( 
.A(n_15149),
.Y(n_15813)
);

OAI22xp5_ASAP7_75t_L g15814 ( 
.A1(n_14894),
.A2(n_1946),
.B1(n_1944),
.B2(n_1945),
.Y(n_15814)
);

INVx1_ASAP7_75t_L g15815 ( 
.A(n_15313),
.Y(n_15815)
);

OAI21x1_ASAP7_75t_L g15816 ( 
.A1(n_15223),
.A2(n_1946),
.B(n_1947),
.Y(n_15816)
);

OA21x2_ASAP7_75t_L g15817 ( 
.A1(n_15233),
.A2(n_1948),
.B(n_1949),
.Y(n_15817)
);

OAI21x1_ASAP7_75t_L g15818 ( 
.A1(n_15235),
.A2(n_15324),
.B(n_15251),
.Y(n_15818)
);

OA21x2_ASAP7_75t_L g15819 ( 
.A1(n_15349),
.A2(n_1949),
.B(n_1950),
.Y(n_15819)
);

OAI21xp5_ASAP7_75t_L g15820 ( 
.A1(n_15182),
.A2(n_1950),
.B(n_1951),
.Y(n_15820)
);

NAND2x1p5_ASAP7_75t_L g15821 ( 
.A(n_15236),
.B(n_1952),
.Y(n_15821)
);

AO21x2_ASAP7_75t_L g15822 ( 
.A1(n_15312),
.A2(n_1952),
.B(n_1953),
.Y(n_15822)
);

NAND2xp5_ASAP7_75t_SL g15823 ( 
.A(n_14892),
.B(n_1953),
.Y(n_15823)
);

INVx2_ASAP7_75t_L g15824 ( 
.A(n_15238),
.Y(n_15824)
);

OAI21x1_ASAP7_75t_L g15825 ( 
.A1(n_15424),
.A2(n_15150),
.B(n_15110),
.Y(n_15825)
);

OAI21x1_ASAP7_75t_L g15826 ( 
.A1(n_15179),
.A2(n_1954),
.B(n_1955),
.Y(n_15826)
);

O2A1O1Ixp33_ASAP7_75t_L g15827 ( 
.A1(n_14975),
.A2(n_1956),
.B(n_1954),
.C(n_1955),
.Y(n_15827)
);

AOI22xp33_ASAP7_75t_L g15828 ( 
.A1(n_14920),
.A2(n_1958),
.B1(n_1956),
.B2(n_1957),
.Y(n_15828)
);

AOI22xp5_ASAP7_75t_L g15829 ( 
.A1(n_15542),
.A2(n_1959),
.B1(n_1957),
.B2(n_1958),
.Y(n_15829)
);

NAND2xp5_ASAP7_75t_L g15830 ( 
.A(n_15248),
.B(n_14995),
.Y(n_15830)
);

BUFx4_ASAP7_75t_SL g15831 ( 
.A(n_14900),
.Y(n_15831)
);

AND2x2_ASAP7_75t_L g15832 ( 
.A(n_15533),
.B(n_15526),
.Y(n_15832)
);

BUFx3_ASAP7_75t_L g15833 ( 
.A(n_15427),
.Y(n_15833)
);

AND2x4_ASAP7_75t_L g15834 ( 
.A(n_15484),
.B(n_1959),
.Y(n_15834)
);

OAI21x1_ASAP7_75t_L g15835 ( 
.A1(n_15190),
.A2(n_1960),
.B(n_1961),
.Y(n_15835)
);

INVx5_ASAP7_75t_L g15836 ( 
.A(n_15476),
.Y(n_15836)
);

OAI21x1_ASAP7_75t_L g15837 ( 
.A1(n_15206),
.A2(n_1960),
.B(n_1961),
.Y(n_15837)
);

INVx2_ASAP7_75t_SL g15838 ( 
.A(n_15089),
.Y(n_15838)
);

AND2x2_ASAP7_75t_L g15839 ( 
.A(n_15485),
.B(n_1962),
.Y(n_15839)
);

AO21x2_ASAP7_75t_L g15840 ( 
.A1(n_15334),
.A2(n_1962),
.B(n_1963),
.Y(n_15840)
);

OR2x2_ASAP7_75t_L g15841 ( 
.A(n_15366),
.B(n_1963),
.Y(n_15841)
);

BUFx6f_ASAP7_75t_L g15842 ( 
.A(n_15143),
.Y(n_15842)
);

INVx2_ASAP7_75t_L g15843 ( 
.A(n_15282),
.Y(n_15843)
);

NOR2xp33_ASAP7_75t_L g15844 ( 
.A(n_15209),
.B(n_1964),
.Y(n_15844)
);

OAI21x1_ASAP7_75t_L g15845 ( 
.A1(n_15288),
.A2(n_15321),
.B(n_15293),
.Y(n_15845)
);

OAI21x1_ASAP7_75t_L g15846 ( 
.A1(n_15326),
.A2(n_1964),
.B(n_1965),
.Y(n_15846)
);

INVx1_ASAP7_75t_L g15847 ( 
.A(n_15328),
.Y(n_15847)
);

AOI22xp33_ASAP7_75t_L g15848 ( 
.A1(n_15536),
.A2(n_1967),
.B1(n_1965),
.B2(n_1966),
.Y(n_15848)
);

BUFx12f_ASAP7_75t_L g15849 ( 
.A(n_15500),
.Y(n_15849)
);

OAI21x1_ASAP7_75t_L g15850 ( 
.A1(n_15003),
.A2(n_1966),
.B(n_1967),
.Y(n_15850)
);

INVx2_ASAP7_75t_SL g15851 ( 
.A(n_15340),
.Y(n_15851)
);

AOI21x1_ASAP7_75t_L g15852 ( 
.A1(n_15117),
.A2(n_1968),
.B(n_1969),
.Y(n_15852)
);

AND2x4_ASAP7_75t_L g15853 ( 
.A(n_15107),
.B(n_1968),
.Y(n_15853)
);

OAI21xp5_ASAP7_75t_L g15854 ( 
.A1(n_15448),
.A2(n_1969),
.B(n_1970),
.Y(n_15854)
);

BUFx3_ASAP7_75t_L g15855 ( 
.A(n_15466),
.Y(n_15855)
);

AO21x2_ASAP7_75t_L g15856 ( 
.A1(n_15357),
.A2(n_1970),
.B(n_1971),
.Y(n_15856)
);

AOI21xp5_ASAP7_75t_L g15857 ( 
.A1(n_14935),
.A2(n_1972),
.B(n_1973),
.Y(n_15857)
);

OAI21x1_ASAP7_75t_L g15858 ( 
.A1(n_15006),
.A2(n_1972),
.B(n_1973),
.Y(n_15858)
);

NAND2xp5_ASAP7_75t_L g15859 ( 
.A(n_15351),
.B(n_1974),
.Y(n_15859)
);

AOI211xp5_ASAP7_75t_L g15860 ( 
.A1(n_14986),
.A2(n_1976),
.B(n_1974),
.C(n_1975),
.Y(n_15860)
);

AOI22x1_ASAP7_75t_L g15861 ( 
.A1(n_15302),
.A2(n_1977),
.B1(n_1975),
.B2(n_1976),
.Y(n_15861)
);

INVx2_ASAP7_75t_L g15862 ( 
.A(n_15506),
.Y(n_15862)
);

O2A1O1Ixp33_ASAP7_75t_SL g15863 ( 
.A1(n_15432),
.A2(n_1979),
.B(n_1977),
.C(n_1978),
.Y(n_15863)
);

OAI21x1_ASAP7_75t_L g15864 ( 
.A1(n_15028),
.A2(n_1978),
.B(n_1980),
.Y(n_15864)
);

INVx1_ASAP7_75t_L g15865 ( 
.A(n_15525),
.Y(n_15865)
);

AND2x4_ASAP7_75t_L g15866 ( 
.A(n_15196),
.B(n_1981),
.Y(n_15866)
);

INVx2_ASAP7_75t_L g15867 ( 
.A(n_15504),
.Y(n_15867)
);

OAI21x1_ASAP7_75t_L g15868 ( 
.A1(n_15062),
.A2(n_1981),
.B(n_1982),
.Y(n_15868)
);

NAND2xp5_ASAP7_75t_L g15869 ( 
.A(n_15527),
.B(n_1982),
.Y(n_15869)
);

INVx2_ASAP7_75t_L g15870 ( 
.A(n_15538),
.Y(n_15870)
);

INVx2_ASAP7_75t_L g15871 ( 
.A(n_15041),
.Y(n_15871)
);

OAI21x1_ASAP7_75t_L g15872 ( 
.A1(n_15131),
.A2(n_1983),
.B(n_1984),
.Y(n_15872)
);

OAI21x1_ASAP7_75t_L g15873 ( 
.A1(n_14957),
.A2(n_1983),
.B(n_1984),
.Y(n_15873)
);

NAND2xp5_ASAP7_75t_L g15874 ( 
.A(n_15385),
.B(n_1985),
.Y(n_15874)
);

INVx1_ASAP7_75t_L g15875 ( 
.A(n_15403),
.Y(n_15875)
);

INVx5_ASAP7_75t_L g15876 ( 
.A(n_15534),
.Y(n_15876)
);

OAI21x1_ASAP7_75t_L g15877 ( 
.A1(n_15253),
.A2(n_1986),
.B(n_1987),
.Y(n_15877)
);

HB1xp67_ASAP7_75t_L g15878 ( 
.A(n_15084),
.Y(n_15878)
);

OAI21x1_ASAP7_75t_L g15879 ( 
.A1(n_14967),
.A2(n_1986),
.B(n_1987),
.Y(n_15879)
);

CKINVDCx5p33_ASAP7_75t_R g15880 ( 
.A(n_15547),
.Y(n_15880)
);

AND2x4_ASAP7_75t_L g15881 ( 
.A(n_15055),
.B(n_1988),
.Y(n_15881)
);

INVx1_ASAP7_75t_L g15882 ( 
.A(n_15566),
.Y(n_15882)
);

OAI211xp5_ASAP7_75t_L g15883 ( 
.A1(n_14955),
.A2(n_1991),
.B(n_1989),
.C(n_1990),
.Y(n_15883)
);

OAI22xp5_ASAP7_75t_L g15884 ( 
.A1(n_15516),
.A2(n_1991),
.B1(n_1989),
.B2(n_1990),
.Y(n_15884)
);

OAI21x1_ASAP7_75t_L g15885 ( 
.A1(n_14974),
.A2(n_1992),
.B(n_1993),
.Y(n_15885)
);

OAI21x1_ASAP7_75t_L g15886 ( 
.A1(n_14977),
.A2(n_1992),
.B(n_1994),
.Y(n_15886)
);

AOI21xp5_ASAP7_75t_L g15887 ( 
.A1(n_14938),
.A2(n_14945),
.B(n_14947),
.Y(n_15887)
);

BUFx6f_ASAP7_75t_L g15888 ( 
.A(n_15143),
.Y(n_15888)
);

OAI22xp5_ASAP7_75t_L g15889 ( 
.A1(n_15540),
.A2(n_15529),
.B1(n_15177),
.B2(n_15436),
.Y(n_15889)
);

AOI21xp5_ASAP7_75t_L g15890 ( 
.A1(n_14904),
.A2(n_1994),
.B(n_1995),
.Y(n_15890)
);

OAI21x1_ASAP7_75t_L g15891 ( 
.A1(n_14991),
.A2(n_1995),
.B(n_1996),
.Y(n_15891)
);

INVx2_ASAP7_75t_L g15892 ( 
.A(n_15332),
.Y(n_15892)
);

OAI21x1_ASAP7_75t_L g15893 ( 
.A1(n_15294),
.A2(n_1996),
.B(n_1997),
.Y(n_15893)
);

AND2x4_ASAP7_75t_L g15894 ( 
.A(n_15546),
.B(n_1997),
.Y(n_15894)
);

OAI22xp5_ASAP7_75t_L g15895 ( 
.A1(n_15170),
.A2(n_2000),
.B1(n_1998),
.B2(n_1999),
.Y(n_15895)
);

OR2x2_ASAP7_75t_L g15896 ( 
.A(n_15558),
.B(n_1998),
.Y(n_15896)
);

OAI21x1_ASAP7_75t_L g15897 ( 
.A1(n_15318),
.A2(n_1999),
.B(n_2000),
.Y(n_15897)
);

OA21x2_ASAP7_75t_L g15898 ( 
.A1(n_15462),
.A2(n_2001),
.B(n_2002),
.Y(n_15898)
);

INVx2_ASAP7_75t_L g15899 ( 
.A(n_15551),
.Y(n_15899)
);

AND2x4_ASAP7_75t_L g15900 ( 
.A(n_15045),
.B(n_2001),
.Y(n_15900)
);

AOI22x1_ASAP7_75t_L g15901 ( 
.A1(n_14865),
.A2(n_2004),
.B1(n_2002),
.B2(n_2003),
.Y(n_15901)
);

INVx3_ASAP7_75t_L g15902 ( 
.A(n_15159),
.Y(n_15902)
);

AOI21xp33_ASAP7_75t_L g15903 ( 
.A1(n_15187),
.A2(n_2003),
.B(n_2004),
.Y(n_15903)
);

INVx1_ASAP7_75t_L g15904 ( 
.A(n_14958),
.Y(n_15904)
);

OAI21x1_ASAP7_75t_L g15905 ( 
.A1(n_15347),
.A2(n_2005),
.B(n_2007),
.Y(n_15905)
);

OAI21x1_ASAP7_75t_L g15906 ( 
.A1(n_15354),
.A2(n_2005),
.B(n_2007),
.Y(n_15906)
);

HB1xp67_ASAP7_75t_L g15907 ( 
.A(n_15376),
.Y(n_15907)
);

AOI21xp5_ASAP7_75t_L g15908 ( 
.A1(n_14908),
.A2(n_15000),
.B(n_14980),
.Y(n_15908)
);

NOR2xp33_ASAP7_75t_SL g15909 ( 
.A(n_15550),
.B(n_2008),
.Y(n_15909)
);

INVx2_ASAP7_75t_L g15910 ( 
.A(n_15554),
.Y(n_15910)
);

BUFx12f_ASAP7_75t_L g15911 ( 
.A(n_15470),
.Y(n_15911)
);

INVx2_ASAP7_75t_L g15912 ( 
.A(n_15158),
.Y(n_15912)
);

OAI21xp5_ASAP7_75t_L g15913 ( 
.A1(n_15480),
.A2(n_15274),
.B(n_15237),
.Y(n_15913)
);

INVx2_ASAP7_75t_L g15914 ( 
.A(n_15555),
.Y(n_15914)
);

NAND2xp5_ASAP7_75t_L g15915 ( 
.A(n_15442),
.B(n_2008),
.Y(n_15915)
);

NAND2xp5_ASAP7_75t_L g15916 ( 
.A(n_15025),
.B(n_2009),
.Y(n_15916)
);

AOI22xp33_ASAP7_75t_L g15917 ( 
.A1(n_15226),
.A2(n_2011),
.B1(n_2009),
.B2(n_2010),
.Y(n_15917)
);

INVx2_ASAP7_75t_L g15918 ( 
.A(n_14973),
.Y(n_15918)
);

INVx1_ASAP7_75t_L g15919 ( 
.A(n_15074),
.Y(n_15919)
);

BUFx2_ASAP7_75t_L g15920 ( 
.A(n_15502),
.Y(n_15920)
);

NOR2xp67_ASAP7_75t_L g15921 ( 
.A(n_15229),
.B(n_2010),
.Y(n_15921)
);

INVx1_ASAP7_75t_L g15922 ( 
.A(n_15098),
.Y(n_15922)
);

AOI21x1_ASAP7_75t_L g15923 ( 
.A1(n_15167),
.A2(n_2011),
.B(n_2012),
.Y(n_15923)
);

OR2x6_ASAP7_75t_L g15924 ( 
.A(n_15319),
.B(n_2012),
.Y(n_15924)
);

OAI21x1_ASAP7_75t_L g15925 ( 
.A1(n_15355),
.A2(n_2013),
.B(n_2014),
.Y(n_15925)
);

OAI21x1_ASAP7_75t_L g15926 ( 
.A1(n_15365),
.A2(n_2013),
.B(n_2014),
.Y(n_15926)
);

INVx1_ASAP7_75t_L g15927 ( 
.A(n_15142),
.Y(n_15927)
);

OAI21x1_ASAP7_75t_L g15928 ( 
.A1(n_15371),
.A2(n_2015),
.B(n_2016),
.Y(n_15928)
);

OAI21x1_ASAP7_75t_L g15929 ( 
.A1(n_15388),
.A2(n_2015),
.B(n_2016),
.Y(n_15929)
);

INVx3_ASAP7_75t_L g15930 ( 
.A(n_15180),
.Y(n_15930)
);

BUFx3_ASAP7_75t_L g15931 ( 
.A(n_15535),
.Y(n_15931)
);

BUFx3_ASAP7_75t_L g15932 ( 
.A(n_15340),
.Y(n_15932)
);

INVx2_ASAP7_75t_L g15933 ( 
.A(n_15201),
.Y(n_15933)
);

AOI21xp5_ASAP7_75t_L g15934 ( 
.A1(n_15010),
.A2(n_2017),
.B(n_2018),
.Y(n_15934)
);

NOR2xp33_ASAP7_75t_L g15935 ( 
.A(n_15418),
.B(n_2017),
.Y(n_15935)
);

AO31x2_ASAP7_75t_L g15936 ( 
.A1(n_14982),
.A2(n_2020),
.A3(n_2018),
.B(n_2019),
.Y(n_15936)
);

OAI21x1_ASAP7_75t_L g15937 ( 
.A1(n_15389),
.A2(n_2019),
.B(n_2020),
.Y(n_15937)
);

OAI21x1_ASAP7_75t_L g15938 ( 
.A1(n_15408),
.A2(n_2021),
.B(n_2022),
.Y(n_15938)
);

INVx1_ASAP7_75t_L g15939 ( 
.A(n_15087),
.Y(n_15939)
);

AO21x2_ASAP7_75t_L g15940 ( 
.A1(n_15370),
.A2(n_15154),
.B(n_15127),
.Y(n_15940)
);

OAI21x1_ASAP7_75t_L g15941 ( 
.A1(n_15410),
.A2(n_2021),
.B(n_2022),
.Y(n_15941)
);

OAI21x1_ASAP7_75t_L g15942 ( 
.A1(n_15421),
.A2(n_2023),
.B(n_2024),
.Y(n_15942)
);

NAND2xp5_ASAP7_75t_L g15943 ( 
.A(n_15440),
.B(n_2023),
.Y(n_15943)
);

OA21x2_ASAP7_75t_L g15944 ( 
.A1(n_15184),
.A2(n_15192),
.B(n_15188),
.Y(n_15944)
);

INVx1_ASAP7_75t_L g15945 ( 
.A(n_15087),
.Y(n_15945)
);

NAND2xp5_ASAP7_75t_L g15946 ( 
.A(n_14890),
.B(n_15479),
.Y(n_15946)
);

A2O1A1Ixp33_ASAP7_75t_L g15947 ( 
.A1(n_15378),
.A2(n_2027),
.B(n_2025),
.C(n_2026),
.Y(n_15947)
);

INVx4_ASAP7_75t_L g15948 ( 
.A(n_15416),
.Y(n_15948)
);

AOI22xp33_ASAP7_75t_L g15949 ( 
.A1(n_15297),
.A2(n_2027),
.B1(n_2025),
.B2(n_2026),
.Y(n_15949)
);

A2O1A1Ixp33_ASAP7_75t_L g15950 ( 
.A1(n_15505),
.A2(n_2030),
.B(n_2028),
.C(n_2029),
.Y(n_15950)
);

OAI21x1_ASAP7_75t_L g15951 ( 
.A1(n_15367),
.A2(n_15284),
.B(n_15434),
.Y(n_15951)
);

INVx1_ASAP7_75t_L g15952 ( 
.A(n_15095),
.Y(n_15952)
);

AND2x2_ASAP7_75t_L g15953 ( 
.A(n_15556),
.B(n_2028),
.Y(n_15953)
);

OAI22xp5_ASAP7_75t_L g15954 ( 
.A1(n_15303),
.A2(n_2032),
.B1(n_2030),
.B2(n_2031),
.Y(n_15954)
);

AO31x2_ASAP7_75t_L g15955 ( 
.A1(n_14968),
.A2(n_2033),
.A3(n_2031),
.B(n_2032),
.Y(n_15955)
);

INVx2_ASAP7_75t_L g15956 ( 
.A(n_14949),
.Y(n_15956)
);

OAI211xp5_ASAP7_75t_L g15957 ( 
.A1(n_15166),
.A2(n_2035),
.B(n_2033),
.C(n_2034),
.Y(n_15957)
);

OAI21x1_ASAP7_75t_L g15958 ( 
.A1(n_15481),
.A2(n_2034),
.B(n_2035),
.Y(n_15958)
);

AND2x2_ASAP7_75t_L g15959 ( 
.A(n_15556),
.B(n_2036),
.Y(n_15959)
);

BUFx3_ASAP7_75t_L g15960 ( 
.A(n_15416),
.Y(n_15960)
);

OAI21x1_ASAP7_75t_L g15961 ( 
.A1(n_15460),
.A2(n_2036),
.B(n_2037),
.Y(n_15961)
);

INVx1_ASAP7_75t_L g15962 ( 
.A(n_15095),
.Y(n_15962)
);

OAI21x1_ASAP7_75t_L g15963 ( 
.A1(n_15483),
.A2(n_15499),
.B(n_15491),
.Y(n_15963)
);

OA21x2_ASAP7_75t_L g15964 ( 
.A1(n_15199),
.A2(n_2038),
.B(n_2039),
.Y(n_15964)
);

OAI21x1_ASAP7_75t_L g15965 ( 
.A1(n_15541),
.A2(n_2038),
.B(n_2039),
.Y(n_15965)
);

OR2x6_ASAP7_75t_L g15966 ( 
.A(n_15319),
.B(n_2040),
.Y(n_15966)
);

NAND2x1p5_ASAP7_75t_L g15967 ( 
.A(n_15109),
.B(n_2040),
.Y(n_15967)
);

OAI22xp5_ASAP7_75t_L g15968 ( 
.A1(n_15304),
.A2(n_2043),
.B1(n_2041),
.B2(n_2042),
.Y(n_15968)
);

INVx1_ASAP7_75t_L g15969 ( 
.A(n_15136),
.Y(n_15969)
);

NAND2xp5_ASAP7_75t_L g15970 ( 
.A(n_15205),
.B(n_2042),
.Y(n_15970)
);

NAND3xp33_ASAP7_75t_L g15971 ( 
.A(n_15441),
.B(n_2043),
.C(n_2044),
.Y(n_15971)
);

AND2x2_ASAP7_75t_L g15972 ( 
.A(n_14953),
.B(n_2044),
.Y(n_15972)
);

AOI21x1_ASAP7_75t_L g15973 ( 
.A1(n_15214),
.A2(n_2045),
.B(n_2046),
.Y(n_15973)
);

INVx1_ASAP7_75t_L g15974 ( 
.A(n_15136),
.Y(n_15974)
);

INVxp67_ASAP7_75t_L g15975 ( 
.A(n_15298),
.Y(n_15975)
);

BUFx3_ASAP7_75t_L g15976 ( 
.A(n_15407),
.Y(n_15976)
);

AOI21x1_ASAP7_75t_L g15977 ( 
.A1(n_15225),
.A2(n_2045),
.B(n_2046),
.Y(n_15977)
);

NAND2xp5_ASAP7_75t_L g15978 ( 
.A(n_15331),
.B(n_2047),
.Y(n_15978)
);

OAI21x1_ASAP7_75t_L g15979 ( 
.A1(n_15323),
.A2(n_2047),
.B(n_2048),
.Y(n_15979)
);

INVx1_ASAP7_75t_L g15980 ( 
.A(n_15040),
.Y(n_15980)
);

CKINVDCx9p33_ASAP7_75t_R g15981 ( 
.A(n_15361),
.Y(n_15981)
);

OAI21x1_ASAP7_75t_L g15982 ( 
.A1(n_15245),
.A2(n_2048),
.B(n_2049),
.Y(n_15982)
);

OA21x2_ASAP7_75t_L g15983 ( 
.A1(n_15247),
.A2(n_2049),
.B(n_2050),
.Y(n_15983)
);

AOI21xp5_ASAP7_75t_L g15984 ( 
.A1(n_15039),
.A2(n_2050),
.B(n_2051),
.Y(n_15984)
);

INVx1_ASAP7_75t_L g15985 ( 
.A(n_15047),
.Y(n_15985)
);

AOI21xp5_ASAP7_75t_L g15986 ( 
.A1(n_15101),
.A2(n_2051),
.B(n_2052),
.Y(n_15986)
);

INVx1_ASAP7_75t_L g15987 ( 
.A(n_15106),
.Y(n_15987)
);

OR2x2_ASAP7_75t_L g15988 ( 
.A(n_15459),
.B(n_2052),
.Y(n_15988)
);

AND2x4_ASAP7_75t_L g15989 ( 
.A(n_14981),
.B(n_2053),
.Y(n_15989)
);

BUFx4_ASAP7_75t_SL g15990 ( 
.A(n_15534),
.Y(n_15990)
);

INVx2_ASAP7_75t_L g15991 ( 
.A(n_15122),
.Y(n_15991)
);

OA21x2_ASAP7_75t_L g15992 ( 
.A1(n_15257),
.A2(n_2053),
.B(n_2054),
.Y(n_15992)
);

NOR2xp33_ASAP7_75t_SL g15993 ( 
.A(n_15430),
.B(n_2054),
.Y(n_15993)
);

AND2x2_ASAP7_75t_L g15994 ( 
.A(n_15015),
.B(n_2055),
.Y(n_15994)
);

INVx2_ASAP7_75t_L g15995 ( 
.A(n_15345),
.Y(n_15995)
);

INVx1_ASAP7_75t_L g15996 ( 
.A(n_15046),
.Y(n_15996)
);

INVx2_ASAP7_75t_L g15997 ( 
.A(n_14981),
.Y(n_15997)
);

INVx1_ASAP7_75t_L g15998 ( 
.A(n_15046),
.Y(n_15998)
);

O2A1O1Ixp33_ASAP7_75t_SL g15999 ( 
.A1(n_15494),
.A2(n_2057),
.B(n_2055),
.C(n_2056),
.Y(n_15999)
);

NAND2xp5_ASAP7_75t_L g16000 ( 
.A(n_15498),
.B(n_15262),
.Y(n_16000)
);

NAND2xp5_ASAP7_75t_L g16001 ( 
.A(n_15276),
.B(n_2056),
.Y(n_16001)
);

OAI21x1_ASAP7_75t_L g16002 ( 
.A1(n_15301),
.A2(n_2057),
.B(n_2058),
.Y(n_16002)
);

OAI21xp5_ASAP7_75t_L g16003 ( 
.A1(n_15518),
.A2(n_2058),
.B(n_2059),
.Y(n_16003)
);

NAND2x1p5_ASAP7_75t_L g16004 ( 
.A(n_15360),
.B(n_2059),
.Y(n_16004)
);

INVx1_ASAP7_75t_L g16005 ( 
.A(n_15413),
.Y(n_16005)
);

OAI21x1_ASAP7_75t_L g16006 ( 
.A1(n_15037),
.A2(n_2060),
.B(n_2061),
.Y(n_16006)
);

NAND2xp5_ASAP7_75t_L g16007 ( 
.A(n_14997),
.B(n_2060),
.Y(n_16007)
);

AOI22xp5_ASAP7_75t_L g16008 ( 
.A1(n_15296),
.A2(n_2064),
.B1(n_2061),
.B2(n_2063),
.Y(n_16008)
);

BUFx6f_ASAP7_75t_L g16009 ( 
.A(n_15145),
.Y(n_16009)
);

AOI221xp5_ASAP7_75t_SL g16010 ( 
.A1(n_14985),
.A2(n_15259),
.B1(n_14962),
.B2(n_15260),
.C(n_15213),
.Y(n_16010)
);

INVx1_ASAP7_75t_L g16011 ( 
.A(n_15426),
.Y(n_16011)
);

CKINVDCx16_ASAP7_75t_R g16012 ( 
.A(n_15036),
.Y(n_16012)
);

OAI21xp5_ASAP7_75t_L g16013 ( 
.A1(n_15093),
.A2(n_2063),
.B(n_2064),
.Y(n_16013)
);

A2O1A1Ixp33_ASAP7_75t_L g16014 ( 
.A1(n_15181),
.A2(n_2068),
.B(n_2065),
.C(n_2066),
.Y(n_16014)
);

OAI22xp5_ASAP7_75t_L g16015 ( 
.A1(n_15308),
.A2(n_2069),
.B1(n_2065),
.B2(n_2068),
.Y(n_16015)
);

INVx1_ASAP7_75t_L g16016 ( 
.A(n_15160),
.Y(n_16016)
);

OAI21xp5_ASAP7_75t_L g16017 ( 
.A1(n_15261),
.A2(n_2069),
.B(n_2070),
.Y(n_16017)
);

BUFx6f_ASAP7_75t_L g16018 ( 
.A(n_15145),
.Y(n_16018)
);

OAI21x1_ASAP7_75t_L g16019 ( 
.A1(n_15449),
.A2(n_2070),
.B(n_2071),
.Y(n_16019)
);

INVx2_ASAP7_75t_L g16020 ( 
.A(n_15005),
.Y(n_16020)
);

INVx1_ASAP7_75t_L g16021 ( 
.A(n_15160),
.Y(n_16021)
);

INVx1_ASAP7_75t_L g16022 ( 
.A(n_15161),
.Y(n_16022)
);

AOI221xp5_ASAP7_75t_L g16023 ( 
.A1(n_15337),
.A2(n_2073),
.B1(n_2071),
.B2(n_2072),
.C(n_2074),
.Y(n_16023)
);

AOI22xp33_ASAP7_75t_L g16024 ( 
.A1(n_15277),
.A2(n_2074),
.B1(n_2072),
.B2(n_2073),
.Y(n_16024)
);

AOI22xp5_ASAP7_75t_L g16025 ( 
.A1(n_14926),
.A2(n_2077),
.B1(n_2075),
.B2(n_2076),
.Y(n_16025)
);

AOI22xp33_ASAP7_75t_L g16026 ( 
.A1(n_15317),
.A2(n_15471),
.B1(n_15397),
.B2(n_15240),
.Y(n_16026)
);

OAI22xp5_ASAP7_75t_L g16027 ( 
.A1(n_15327),
.A2(n_2077),
.B1(n_2075),
.B2(n_2076),
.Y(n_16027)
);

AO21x2_ASAP7_75t_L g16028 ( 
.A1(n_15266),
.A2(n_2078),
.B(n_2080),
.Y(n_16028)
);

INVx2_ASAP7_75t_SL g16029 ( 
.A(n_14972),
.Y(n_16029)
);

OAI22xp33_ASAP7_75t_L g16030 ( 
.A1(n_15162),
.A2(n_2081),
.B1(n_2078),
.B2(n_2080),
.Y(n_16030)
);

INVx2_ASAP7_75t_L g16031 ( 
.A(n_15005),
.Y(n_16031)
);

NOR2xp33_ASAP7_75t_L g16032 ( 
.A(n_15429),
.B(n_2081),
.Y(n_16032)
);

AND2x4_ASAP7_75t_L g16033 ( 
.A(n_15011),
.B(n_2082),
.Y(n_16033)
);

BUFx2_ASAP7_75t_L g16034 ( 
.A(n_15011),
.Y(n_16034)
);

AND2x4_ASAP7_75t_L g16035 ( 
.A(n_15075),
.B(n_2082),
.Y(n_16035)
);

BUFx12f_ASAP7_75t_L g16036 ( 
.A(n_15532),
.Y(n_16036)
);

OAI21x1_ASAP7_75t_L g16037 ( 
.A1(n_15464),
.A2(n_2083),
.B(n_2084),
.Y(n_16037)
);

NAND2x1_ASAP7_75t_L g16038 ( 
.A(n_15522),
.B(n_2083),
.Y(n_16038)
);

INVx3_ASAP7_75t_L g16039 ( 
.A(n_15186),
.Y(n_16039)
);

OAI21x1_ASAP7_75t_L g16040 ( 
.A1(n_15344),
.A2(n_2084),
.B(n_2085),
.Y(n_16040)
);

AND2x4_ASAP7_75t_L g16041 ( 
.A(n_15075),
.B(n_2085),
.Y(n_16041)
);

AOI22xp33_ASAP7_75t_L g16042 ( 
.A1(n_15053),
.A2(n_2088),
.B1(n_2086),
.B2(n_2087),
.Y(n_16042)
);

BUFx6f_ASAP7_75t_L g16043 ( 
.A(n_15186),
.Y(n_16043)
);

OAI21x1_ASAP7_75t_L g16044 ( 
.A1(n_15026),
.A2(n_2086),
.B(n_2087),
.Y(n_16044)
);

NAND2x1p5_ASAP7_75t_L g16045 ( 
.A(n_15530),
.B(n_2088),
.Y(n_16045)
);

AOI22xp33_ASAP7_75t_L g16046 ( 
.A1(n_14994),
.A2(n_2091),
.B1(n_2089),
.B2(n_2090),
.Y(n_16046)
);

INVx1_ASAP7_75t_L g16047 ( 
.A(n_15161),
.Y(n_16047)
);

INVx2_ASAP7_75t_L g16048 ( 
.A(n_15234),
.Y(n_16048)
);

INVx1_ASAP7_75t_L g16049 ( 
.A(n_14970),
.Y(n_16049)
);

A2O1A1Ixp33_ASAP7_75t_L g16050 ( 
.A1(n_15067),
.A2(n_2091),
.B(n_2089),
.C(n_2090),
.Y(n_16050)
);

AO31x2_ASAP7_75t_L g16051 ( 
.A1(n_15152),
.A2(n_15219),
.A3(n_15287),
.B(n_15168),
.Y(n_16051)
);

INVx2_ASAP7_75t_L g16052 ( 
.A(n_15315),
.Y(n_16052)
);

AOI22xp33_ASAP7_75t_L g16053 ( 
.A1(n_15001),
.A2(n_2094),
.B1(n_2092),
.B2(n_2093),
.Y(n_16053)
);

AO31x2_ASAP7_75t_L g16054 ( 
.A1(n_15404),
.A2(n_2094),
.A3(n_2092),
.B(n_2093),
.Y(n_16054)
);

INVx2_ASAP7_75t_L g16055 ( 
.A(n_15307),
.Y(n_16055)
);

OAI22xp5_ASAP7_75t_L g16056 ( 
.A1(n_15333),
.A2(n_2097),
.B1(n_2095),
.B2(n_2096),
.Y(n_16056)
);

OAI21x1_ASAP7_75t_L g16057 ( 
.A1(n_15269),
.A2(n_2095),
.B(n_2097),
.Y(n_16057)
);

NAND2x1p5_ASAP7_75t_L g16058 ( 
.A(n_15171),
.B(n_2098),
.Y(n_16058)
);

NOR2xp33_ASAP7_75t_L g16059 ( 
.A(n_15444),
.B(n_2098),
.Y(n_16059)
);

INVx1_ASAP7_75t_L g16060 ( 
.A(n_14970),
.Y(n_16060)
);

OA21x2_ASAP7_75t_L g16061 ( 
.A1(n_15273),
.A2(n_2099),
.B(n_2100),
.Y(n_16061)
);

NOR2xp67_ASAP7_75t_L g16062 ( 
.A(n_15472),
.B(n_15568),
.Y(n_16062)
);

HB1xp67_ASAP7_75t_L g16063 ( 
.A(n_15487),
.Y(n_16063)
);

INVx1_ASAP7_75t_L g16064 ( 
.A(n_15230),
.Y(n_16064)
);

NAND2xp5_ASAP7_75t_L g16065 ( 
.A(n_15402),
.B(n_2099),
.Y(n_16065)
);

INVx2_ASAP7_75t_L g16066 ( 
.A(n_15322),
.Y(n_16066)
);

INVx1_ASAP7_75t_L g16067 ( 
.A(n_15230),
.Y(n_16067)
);

INVx2_ASAP7_75t_SL g16068 ( 
.A(n_15200),
.Y(n_16068)
);

CKINVDCx6p67_ASAP7_75t_R g16069 ( 
.A(n_15522),
.Y(n_16069)
);

INVx3_ASAP7_75t_SL g16070 ( 
.A(n_15200),
.Y(n_16070)
);

OAI21x1_ASAP7_75t_SL g16071 ( 
.A1(n_15271),
.A2(n_15514),
.B(n_15486),
.Y(n_16071)
);

AOI21xp5_ASAP7_75t_L g16072 ( 
.A1(n_15290),
.A2(n_2100),
.B(n_2101),
.Y(n_16072)
);

INVx1_ASAP7_75t_L g16073 ( 
.A(n_15252),
.Y(n_16073)
);

INVx1_ASAP7_75t_L g16074 ( 
.A(n_15252),
.Y(n_16074)
);

INVx1_ASAP7_75t_L g16075 ( 
.A(n_15272),
.Y(n_16075)
);

OAI21xp5_ASAP7_75t_L g16076 ( 
.A1(n_15115),
.A2(n_15065),
.B(n_15121),
.Y(n_16076)
);

NAND2xp5_ASAP7_75t_L g16077 ( 
.A(n_15310),
.B(n_2101),
.Y(n_16077)
);

OAI21x1_ASAP7_75t_L g16078 ( 
.A1(n_15539),
.A2(n_2102),
.B(n_2103),
.Y(n_16078)
);

AOI21xp5_ASAP7_75t_L g16079 ( 
.A1(n_15002),
.A2(n_2102),
.B(n_2103),
.Y(n_16079)
);

OA21x2_ASAP7_75t_L g16080 ( 
.A1(n_15457),
.A2(n_2104),
.B(n_2105),
.Y(n_16080)
);

NAND2xp5_ASAP7_75t_L g16081 ( 
.A(n_15468),
.B(n_2104),
.Y(n_16081)
);

NAND3x1_ASAP7_75t_L g16082 ( 
.A(n_15348),
.B(n_15020),
.C(n_15279),
.Y(n_16082)
);

AOI21x1_ASAP7_75t_L g16083 ( 
.A1(n_14869),
.A2(n_2105),
.B(n_2106),
.Y(n_16083)
);

OAI22xp5_ASAP7_75t_L g16084 ( 
.A1(n_15552),
.A2(n_2109),
.B1(n_2106),
.B2(n_2107),
.Y(n_16084)
);

INVx3_ASAP7_75t_L g16085 ( 
.A(n_15742),
.Y(n_16085)
);

INVx3_ASAP7_75t_L g16086 ( 
.A(n_15684),
.Y(n_16086)
);

OA21x2_ASAP7_75t_L g16087 ( 
.A1(n_15577),
.A2(n_15455),
.B(n_14877),
.Y(n_16087)
);

AND2x2_ASAP7_75t_L g16088 ( 
.A(n_15616),
.B(n_15336),
.Y(n_16088)
);

NAND2xp5_ASAP7_75t_L g16089 ( 
.A(n_15610),
.B(n_15487),
.Y(n_16089)
);

NOR2xp67_ASAP7_75t_L g16090 ( 
.A(n_15625),
.B(n_15207),
.Y(n_16090)
);

INVx1_ASAP7_75t_L g16091 ( 
.A(n_15703),
.Y(n_16091)
);

AND2x4_ASAP7_75t_L g16092 ( 
.A(n_15569),
.B(n_15411),
.Y(n_16092)
);

AND2x2_ASAP7_75t_L g16093 ( 
.A(n_15735),
.B(n_15598),
.Y(n_16093)
);

AND2x2_ASAP7_75t_L g16094 ( 
.A(n_15724),
.B(n_15336),
.Y(n_16094)
);

OR2x2_ASAP7_75t_L g16095 ( 
.A(n_15626),
.B(n_15451),
.Y(n_16095)
);

INVx2_ASAP7_75t_L g16096 ( 
.A(n_15681),
.Y(n_16096)
);

A2O1A1Ixp33_ASAP7_75t_L g16097 ( 
.A1(n_15887),
.A2(n_15280),
.B(n_15428),
.C(n_15417),
.Y(n_16097)
);

AOI211xp5_ASAP7_75t_L g16098 ( 
.A1(n_15777),
.A2(n_15563),
.B(n_15543),
.C(n_15102),
.Y(n_16098)
);

NOR2xp67_ASAP7_75t_L g16099 ( 
.A(n_15625),
.B(n_15286),
.Y(n_16099)
);

OR2x2_ASAP7_75t_L g16100 ( 
.A(n_15692),
.B(n_15496),
.Y(n_16100)
);

INVx1_ASAP7_75t_L g16101 ( 
.A(n_15708),
.Y(n_16101)
);

OR2x2_ASAP7_75t_L g16102 ( 
.A(n_15867),
.B(n_15509),
.Y(n_16102)
);

NOR2xp67_ASAP7_75t_L g16103 ( 
.A(n_15836),
.B(n_15812),
.Y(n_16103)
);

AND2x4_ASAP7_75t_L g16104 ( 
.A(n_15672),
.B(n_15411),
.Y(n_16104)
);

AOI21xp5_ASAP7_75t_L g16105 ( 
.A1(n_15594),
.A2(n_15202),
.B(n_15350),
.Y(n_16105)
);

CKINVDCx5p33_ASAP7_75t_R g16106 ( 
.A(n_15880),
.Y(n_16106)
);

INVx3_ASAP7_75t_L g16107 ( 
.A(n_15575),
.Y(n_16107)
);

OR2x2_ASAP7_75t_L g16108 ( 
.A(n_15800),
.B(n_15520),
.Y(n_16108)
);

AOI21xp5_ASAP7_75t_L g16109 ( 
.A1(n_15784),
.A2(n_15908),
.B(n_15913),
.Y(n_16109)
);

AND2x2_ASAP7_75t_L g16110 ( 
.A(n_15619),
.B(n_15007),
.Y(n_16110)
);

INVx1_ASAP7_75t_L g16111 ( 
.A(n_15574),
.Y(n_16111)
);

NAND2xp5_ASAP7_75t_L g16112 ( 
.A(n_15946),
.B(n_15537),
.Y(n_16112)
);

OAI22xp5_ASAP7_75t_L g16113 ( 
.A1(n_15607),
.A2(n_15567),
.B1(n_15012),
.B2(n_15052),
.Y(n_16113)
);

INVx1_ASAP7_75t_L g16114 ( 
.A(n_15587),
.Y(n_16114)
);

AOI21x1_ASAP7_75t_SL g16115 ( 
.A1(n_16000),
.A2(n_15450),
.B(n_15419),
.Y(n_16115)
);

NOR2xp33_ASAP7_75t_L g16116 ( 
.A(n_15642),
.B(n_15079),
.Y(n_16116)
);

NAND2xp5_ASAP7_75t_L g16117 ( 
.A(n_15940),
.B(n_15537),
.Y(n_16117)
);

INVxp67_ASAP7_75t_SL g16118 ( 
.A(n_15629),
.Y(n_16118)
);

NAND2xp5_ASAP7_75t_L g16119 ( 
.A(n_15944),
.B(n_15221),
.Y(n_16119)
);

A2O1A1Ixp33_ASAP7_75t_L g16120 ( 
.A1(n_15890),
.A2(n_15373),
.B(n_15341),
.C(n_15338),
.Y(n_16120)
);

NAND2xp5_ASAP7_75t_L g16121 ( 
.A(n_15636),
.B(n_15221),
.Y(n_16121)
);

NOR2xp67_ASAP7_75t_L g16122 ( 
.A(n_15836),
.B(n_15311),
.Y(n_16122)
);

INVx1_ASAP7_75t_L g16123 ( 
.A(n_15612),
.Y(n_16123)
);

O2A1O1Ixp33_ASAP7_75t_L g16124 ( 
.A1(n_15804),
.A2(n_15018),
.B(n_15064),
.C(n_15054),
.Y(n_16124)
);

CKINVDCx5p33_ASAP7_75t_R g16125 ( 
.A(n_15694),
.Y(n_16125)
);

AND2x4_ASAP7_75t_L g16126 ( 
.A(n_15634),
.B(n_15314),
.Y(n_16126)
);

AND2x2_ASAP7_75t_L g16127 ( 
.A(n_15685),
.B(n_15412),
.Y(n_16127)
);

INVx1_ASAP7_75t_L g16128 ( 
.A(n_15614),
.Y(n_16128)
);

CKINVDCx20_ASAP7_75t_R g16129 ( 
.A(n_15780),
.Y(n_16129)
);

AOI21xp5_ASAP7_75t_L g16130 ( 
.A1(n_15803),
.A2(n_15391),
.B(n_15382),
.Y(n_16130)
);

AND2x2_ASAP7_75t_L g16131 ( 
.A(n_15727),
.B(n_15412),
.Y(n_16131)
);

INVx1_ASAP7_75t_L g16132 ( 
.A(n_15622),
.Y(n_16132)
);

INVxp67_ASAP7_75t_L g16133 ( 
.A(n_15907),
.Y(n_16133)
);

INVx2_ASAP7_75t_L g16134 ( 
.A(n_15845),
.Y(n_16134)
);

A2O1A1Ixp33_ASAP7_75t_L g16135 ( 
.A1(n_15715),
.A2(n_15475),
.B(n_15085),
.C(n_15224),
.Y(n_16135)
);

HB1xp67_ASAP7_75t_L g16136 ( 
.A(n_15591),
.Y(n_16136)
);

NAND2xp5_ASAP7_75t_L g16137 ( 
.A(n_15579),
.B(n_15611),
.Y(n_16137)
);

NAND2x1p5_ASAP7_75t_L g16138 ( 
.A(n_15656),
.B(n_15669),
.Y(n_16138)
);

NOR2x2_ASAP7_75t_L g16139 ( 
.A(n_15663),
.B(n_15105),
.Y(n_16139)
);

INVx1_ASAP7_75t_SL g16140 ( 
.A(n_15981),
.Y(n_16140)
);

AND2x4_ASAP7_75t_L g16141 ( 
.A(n_15623),
.B(n_15314),
.Y(n_16141)
);

AOI21xp5_ASAP7_75t_L g16142 ( 
.A1(n_15599),
.A2(n_15519),
.B(n_15422),
.Y(n_16142)
);

INVx2_ASAP7_75t_L g16143 ( 
.A(n_15818),
.Y(n_16143)
);

OAI22xp5_ASAP7_75t_L g16144 ( 
.A1(n_16026),
.A2(n_15387),
.B1(n_15386),
.B2(n_15212),
.Y(n_16144)
);

INVx2_ASAP7_75t_L g16145 ( 
.A(n_15743),
.Y(n_16145)
);

INVx1_ASAP7_75t_L g16146 ( 
.A(n_15633),
.Y(n_16146)
);

AOI21x1_ASAP7_75t_SL g16147 ( 
.A1(n_15970),
.A2(n_15105),
.B(n_14987),
.Y(n_16147)
);

INVx1_ASAP7_75t_L g16148 ( 
.A(n_15637),
.Y(n_16148)
);

NAND2xp5_ASAP7_75t_L g16149 ( 
.A(n_15609),
.B(n_15019),
.Y(n_16149)
);

OR2x2_ASAP7_75t_L g16150 ( 
.A(n_15680),
.B(n_15339),
.Y(n_16150)
);

BUFx6f_ASAP7_75t_L g16151 ( 
.A(n_15643),
.Y(n_16151)
);

OAI22xp5_ASAP7_75t_L g16152 ( 
.A1(n_15829),
.A2(n_15175),
.B1(n_15208),
.B2(n_15320),
.Y(n_16152)
);

OAI22xp5_ASAP7_75t_L g16153 ( 
.A1(n_16082),
.A2(n_15393),
.B1(n_15512),
.B2(n_15364),
.Y(n_16153)
);

AND2x2_ASAP7_75t_L g16154 ( 
.A(n_15824),
.B(n_15335),
.Y(n_16154)
);

AOI21xp5_ASAP7_75t_L g16155 ( 
.A1(n_15857),
.A2(n_15140),
.B(n_15138),
.Y(n_16155)
);

OR2x6_ASAP7_75t_L g16156 ( 
.A(n_15621),
.B(n_15094),
.Y(n_16156)
);

NAND2xp5_ASAP7_75t_L g16157 ( 
.A(n_15689),
.B(n_15339),
.Y(n_16157)
);

AND2x4_ASAP7_75t_L g16158 ( 
.A(n_15646),
.B(n_15346),
.Y(n_16158)
);

A2O1A1Ixp33_ASAP7_75t_L g16159 ( 
.A1(n_15820),
.A2(n_15038),
.B(n_15545),
.C(n_15392),
.Y(n_16159)
);

AND2x2_ASAP7_75t_L g16160 ( 
.A(n_15699),
.B(n_15562),
.Y(n_16160)
);

CKINVDCx20_ASAP7_75t_R g16161 ( 
.A(n_15628),
.Y(n_16161)
);

NAND2xp5_ASAP7_75t_L g16162 ( 
.A(n_15638),
.B(n_15346),
.Y(n_16162)
);

A2O1A1Ixp33_ASAP7_75t_L g16163 ( 
.A1(n_16076),
.A2(n_15049),
.B(n_15372),
.C(n_15353),
.Y(n_16163)
);

AND2x2_ASAP7_75t_L g16164 ( 
.A(n_15645),
.B(n_14888),
.Y(n_16164)
);

AND2x2_ASAP7_75t_L g16165 ( 
.A(n_15832),
.B(n_16034),
.Y(n_16165)
);

AOI21xp5_ASAP7_75t_SL g16166 ( 
.A1(n_15797),
.A2(n_15493),
.B(n_15511),
.Y(n_16166)
);

AND2x2_ASAP7_75t_L g16167 ( 
.A(n_15660),
.B(n_14888),
.Y(n_16167)
);

AOI21xp5_ASAP7_75t_L g16168 ( 
.A1(n_15903),
.A2(n_15195),
.B(n_15193),
.Y(n_16168)
);

INVx2_ASAP7_75t_SL g16169 ( 
.A(n_15831),
.Y(n_16169)
);

OR2x2_ASAP7_75t_L g16170 ( 
.A(n_15871),
.B(n_15559),
.Y(n_16170)
);

AND2x4_ASAP7_75t_L g16171 ( 
.A(n_15920),
.B(n_15454),
.Y(n_16171)
);

BUFx10_ASAP7_75t_L g16172 ( 
.A(n_15935),
.Y(n_16172)
);

INVx2_ASAP7_75t_L g16173 ( 
.A(n_15843),
.Y(n_16173)
);

NOR2xp67_ASAP7_75t_L g16174 ( 
.A(n_15876),
.B(n_15099),
.Y(n_16174)
);

AND2x2_ASAP7_75t_L g16175 ( 
.A(n_15892),
.B(n_15454),
.Y(n_16175)
);

INVx3_ASAP7_75t_L g16176 ( 
.A(n_15711),
.Y(n_16176)
);

AOI21xp5_ASAP7_75t_L g16177 ( 
.A1(n_15662),
.A2(n_15381),
.B(n_15377),
.Y(n_16177)
);

INVx1_ASAP7_75t_L g16178 ( 
.A(n_15650),
.Y(n_16178)
);

NAND2xp5_ASAP7_75t_L g16179 ( 
.A(n_15602),
.B(n_15559),
.Y(n_16179)
);

INVx2_ASAP7_75t_L g16180 ( 
.A(n_15862),
.Y(n_16180)
);

AOI21xp5_ASAP7_75t_SL g16181 ( 
.A1(n_15827),
.A2(n_15565),
.B(n_14990),
.Y(n_16181)
);

AND2x2_ASAP7_75t_L g16182 ( 
.A(n_15714),
.B(n_15691),
.Y(n_16182)
);

NAND2xp5_ASAP7_75t_L g16183 ( 
.A(n_15603),
.B(n_15272),
.Y(n_16183)
);

AND2x4_ASAP7_75t_L g16184 ( 
.A(n_15902),
.B(n_15456),
.Y(n_16184)
);

AOI21xp5_ASAP7_75t_L g16185 ( 
.A1(n_15889),
.A2(n_15042),
.B(n_15191),
.Y(n_16185)
);

NAND2xp5_ASAP7_75t_L g16186 ( 
.A(n_15754),
.B(n_15289),
.Y(n_16186)
);

O2A1O1Ixp5_ASAP7_75t_L g16187 ( 
.A1(n_15957),
.A2(n_15933),
.B(n_15995),
.C(n_15919),
.Y(n_16187)
);

INVx2_ASAP7_75t_SL g16188 ( 
.A(n_15570),
.Y(n_16188)
);

AND2x4_ASAP7_75t_L g16189 ( 
.A(n_15930),
.B(n_15456),
.Y(n_16189)
);

INVx1_ASAP7_75t_L g16190 ( 
.A(n_15654),
.Y(n_16190)
);

HB1xp67_ASAP7_75t_L g16191 ( 
.A(n_15739),
.Y(n_16191)
);

NAND2xp5_ASAP7_75t_L g16192 ( 
.A(n_15618),
.B(n_15289),
.Y(n_16192)
);

NOR2xp33_ASAP7_75t_L g16193 ( 
.A(n_15664),
.B(n_15453),
.Y(n_16193)
);

INVx2_ASAP7_75t_L g16194 ( 
.A(n_15773),
.Y(n_16194)
);

BUFx8_ASAP7_75t_SL g16195 ( 
.A(n_15643),
.Y(n_16195)
);

AND2x2_ASAP7_75t_L g16196 ( 
.A(n_15713),
.B(n_15414),
.Y(n_16196)
);

AND2x4_ASAP7_75t_L g16197 ( 
.A(n_15706),
.B(n_15659),
.Y(n_16197)
);

INVx2_ASAP7_75t_L g16198 ( 
.A(n_15774),
.Y(n_16198)
);

INVx1_ASAP7_75t_L g16199 ( 
.A(n_15666),
.Y(n_16199)
);

CKINVDCx20_ASAP7_75t_R g16200 ( 
.A(n_15749),
.Y(n_16200)
);

INVxp67_ASAP7_75t_L g16201 ( 
.A(n_15635),
.Y(n_16201)
);

HB1xp67_ASAP7_75t_L g16202 ( 
.A(n_15676),
.Y(n_16202)
);

AND2x2_ASAP7_75t_L g16203 ( 
.A(n_15641),
.B(n_15414),
.Y(n_16203)
);

AND2x4_ASAP7_75t_L g16204 ( 
.A(n_15663),
.B(n_15731),
.Y(n_16204)
);

NAND2xp5_ASAP7_75t_L g16205 ( 
.A(n_15618),
.B(n_15423),
.Y(n_16205)
);

AOI21xp5_ASAP7_75t_L g16206 ( 
.A1(n_15752),
.A2(n_15405),
.B(n_15452),
.Y(n_16206)
);

O2A1O1Ixp33_ASAP7_75t_SL g16207 ( 
.A1(n_16038),
.A2(n_15523),
.B(n_15553),
.C(n_14987),
.Y(n_16207)
);

INVx1_ASAP7_75t_L g16208 ( 
.A(n_15671),
.Y(n_16208)
);

AND2x4_ASAP7_75t_L g16209 ( 
.A(n_15833),
.B(n_15423),
.Y(n_16209)
);

INVx2_ASAP7_75t_L g16210 ( 
.A(n_15783),
.Y(n_16210)
);

BUFx3_ASAP7_75t_L g16211 ( 
.A(n_15849),
.Y(n_16211)
);

A2O1A1Ixp33_ASAP7_75t_L g16212 ( 
.A1(n_15860),
.A2(n_15292),
.B(n_14965),
.C(n_15135),
.Y(n_16212)
);

AND2x2_ASAP7_75t_L g16213 ( 
.A(n_15698),
.B(n_15431),
.Y(n_16213)
);

NAND2xp5_ASAP7_75t_L g16214 ( 
.A(n_15980),
.B(n_15431),
.Y(n_16214)
);

AND2x4_ASAP7_75t_L g16215 ( 
.A(n_15855),
.B(n_15931),
.Y(n_16215)
);

INVx3_ASAP7_75t_L g16216 ( 
.A(n_15813),
.Y(n_16216)
);

INVx1_ASAP7_75t_SL g16217 ( 
.A(n_15613),
.Y(n_16217)
);

NAND2xp5_ASAP7_75t_L g16218 ( 
.A(n_15985),
.B(n_15151),
.Y(n_16218)
);

NOR2xp33_ASAP7_75t_L g16219 ( 
.A(n_15794),
.B(n_15035),
.Y(n_16219)
);

AND2x2_ASAP7_75t_L g16220 ( 
.A(n_15583),
.B(n_15589),
.Y(n_16220)
);

AND2x2_ASAP7_75t_L g16221 ( 
.A(n_15590),
.B(n_14909),
.Y(n_16221)
);

AO22x2_ASAP7_75t_L g16222 ( 
.A1(n_15975),
.A2(n_15524),
.B1(n_15258),
.B2(n_15305),
.Y(n_16222)
);

INVx1_ASAP7_75t_L g16223 ( 
.A(n_15682),
.Y(n_16223)
);

AND2x2_ASAP7_75t_L g16224 ( 
.A(n_15617),
.B(n_14909),
.Y(n_16224)
);

A2O1A1Ixp33_ASAP7_75t_SL g16225 ( 
.A1(n_15854),
.A2(n_15406),
.B(n_15057),
.C(n_15014),
.Y(n_16225)
);

INVx2_ASAP7_75t_L g16226 ( 
.A(n_15788),
.Y(n_16226)
);

OR2x2_ASAP7_75t_L g16227 ( 
.A(n_15904),
.B(n_15151),
.Y(n_16227)
);

NOR2xp33_ASAP7_75t_L g16228 ( 
.A(n_15596),
.B(n_15648),
.Y(n_16228)
);

NOR2x2_ASAP7_75t_L g16229 ( 
.A(n_15776),
.B(n_15415),
.Y(n_16229)
);

INVxp67_ASAP7_75t_L g16230 ( 
.A(n_15898),
.Y(n_16230)
);

AND2x2_ASAP7_75t_L g16231 ( 
.A(n_15914),
.B(n_14873),
.Y(n_16231)
);

INVx1_ASAP7_75t_SL g16232 ( 
.A(n_15990),
.Y(n_16232)
);

NAND2xp5_ASAP7_75t_L g16233 ( 
.A(n_15987),
.B(n_16005),
.Y(n_16233)
);

INVx2_ASAP7_75t_L g16234 ( 
.A(n_15806),
.Y(n_16234)
);

AND2x2_ASAP7_75t_L g16235 ( 
.A(n_15878),
.B(n_14873),
.Y(n_16235)
);

AOI21xp5_ASAP7_75t_L g16236 ( 
.A1(n_15756),
.A2(n_15934),
.B(n_15807),
.Y(n_16236)
);

INVx1_ASAP7_75t_L g16237 ( 
.A(n_15604),
.Y(n_16237)
);

INVx1_ASAP7_75t_L g16238 ( 
.A(n_15709),
.Y(n_16238)
);

INVx1_ASAP7_75t_L g16239 ( 
.A(n_15718),
.Y(n_16239)
);

AND2x2_ASAP7_75t_L g16240 ( 
.A(n_15657),
.B(n_15183),
.Y(n_16240)
);

INVx1_ASAP7_75t_L g16241 ( 
.A(n_15799),
.Y(n_16241)
);

NAND2xp5_ASAP7_75t_L g16242 ( 
.A(n_16011),
.B(n_15228),
.Y(n_16242)
);

AOI21xp5_ASAP7_75t_L g16243 ( 
.A1(n_15734),
.A2(n_15250),
.B(n_15263),
.Y(n_16243)
);

NAND2xp5_ASAP7_75t_L g16244 ( 
.A(n_15572),
.B(n_15560),
.Y(n_16244)
);

AND2x2_ASAP7_75t_L g16245 ( 
.A(n_15595),
.B(n_15508),
.Y(n_16245)
);

NAND2xp5_ASAP7_75t_L g16246 ( 
.A(n_15576),
.B(n_15503),
.Y(n_16246)
);

OA21x2_ASAP7_75t_L g16247 ( 
.A1(n_15584),
.A2(n_15517),
.B(n_15077),
.Y(n_16247)
);

INVx2_ASAP7_75t_L g16248 ( 
.A(n_15811),
.Y(n_16248)
);

NOR2xp67_ASAP7_75t_L g16249 ( 
.A(n_15876),
.B(n_15267),
.Y(n_16249)
);

AND2x4_ASAP7_75t_L g16250 ( 
.A(n_15588),
.B(n_15398),
.Y(n_16250)
);

NAND2xp5_ASAP7_75t_L g16251 ( 
.A(n_15581),
.B(n_15725),
.Y(n_16251)
);

INVx1_ASAP7_75t_L g16252 ( 
.A(n_15802),
.Y(n_16252)
);

BUFx6f_ASAP7_75t_L g16253 ( 
.A(n_15667),
.Y(n_16253)
);

INVx1_ASAP7_75t_L g16254 ( 
.A(n_15815),
.Y(n_16254)
);

INVx3_ASAP7_75t_SL g16255 ( 
.A(n_15924),
.Y(n_16255)
);

INVx2_ASAP7_75t_L g16256 ( 
.A(n_15693),
.Y(n_16256)
);

NOR2xp33_ASAP7_75t_L g16257 ( 
.A(n_15688),
.B(n_15330),
.Y(n_16257)
);

AOI21xp5_ASAP7_75t_L g16258 ( 
.A1(n_15947),
.A2(n_15070),
.B(n_15063),
.Y(n_16258)
);

INVx2_ASAP7_75t_L g16259 ( 
.A(n_15702),
.Y(n_16259)
);

AND2x2_ASAP7_75t_L g16260 ( 
.A(n_15997),
.B(n_15189),
.Y(n_16260)
);

INVx1_ASAP7_75t_L g16261 ( 
.A(n_15733),
.Y(n_16261)
);

INVx1_ASAP7_75t_L g16262 ( 
.A(n_15737),
.Y(n_16262)
);

NAND2xp5_ASAP7_75t_L g16263 ( 
.A(n_16063),
.B(n_15510),
.Y(n_16263)
);

AND2x2_ASAP7_75t_L g16264 ( 
.A(n_16020),
.B(n_15189),
.Y(n_16264)
);

NAND2xp5_ASAP7_75t_L g16265 ( 
.A(n_15757),
.B(n_15104),
.Y(n_16265)
);

INVxp67_ASAP7_75t_L g16266 ( 
.A(n_16080),
.Y(n_16266)
);

NAND2xp5_ASAP7_75t_L g16267 ( 
.A(n_15922),
.B(n_15165),
.Y(n_16267)
);

O2A1O1Ixp33_ASAP7_75t_L g16268 ( 
.A1(n_15999),
.A2(n_15420),
.B(n_14950),
.C(n_14952),
.Y(n_16268)
);

NOR2xp33_ASAP7_75t_L g16269 ( 
.A(n_15948),
.B(n_15278),
.Y(n_16269)
);

NAND2xp5_ASAP7_75t_L g16270 ( 
.A(n_15927),
.B(n_15285),
.Y(n_16270)
);

INVxp67_ASAP7_75t_L g16271 ( 
.A(n_15964),
.Y(n_16271)
);

BUFx6f_ASAP7_75t_L g16272 ( 
.A(n_15667),
.Y(n_16272)
);

INVx1_ASAP7_75t_SL g16273 ( 
.A(n_15683),
.Y(n_16273)
);

AOI21xp5_ASAP7_75t_L g16274 ( 
.A1(n_15786),
.A2(n_15244),
.B(n_15242),
.Y(n_16274)
);

AND2x4_ASAP7_75t_L g16275 ( 
.A(n_15838),
.B(n_15467),
.Y(n_16275)
);

OR2x6_ASAP7_75t_L g16276 ( 
.A(n_15631),
.B(n_15083),
.Y(n_16276)
);

INVx3_ASAP7_75t_L g16277 ( 
.A(n_15746),
.Y(n_16277)
);

CKINVDCx12_ASAP7_75t_R g16278 ( 
.A(n_15924),
.Y(n_16278)
);

BUFx6f_ASAP7_75t_L g16279 ( 
.A(n_15932),
.Y(n_16279)
);

NOR2xp33_ASAP7_75t_L g16280 ( 
.A(n_16012),
.B(n_15383),
.Y(n_16280)
);

A2O1A1Ixp33_ASAP7_75t_L g16281 ( 
.A1(n_16025),
.A2(n_15016),
.B(n_14979),
.C(n_15215),
.Y(n_16281)
);

NAND2xp5_ASAP7_75t_L g16282 ( 
.A(n_15620),
.B(n_15111),
.Y(n_16282)
);

OAI22xp5_ASAP7_75t_L g16283 ( 
.A1(n_16008),
.A2(n_15528),
.B1(n_15048),
.B2(n_15249),
.Y(n_16283)
);

AOI21xp5_ASAP7_75t_L g16284 ( 
.A1(n_16072),
.A2(n_15123),
.B(n_15227),
.Y(n_16284)
);

INVx1_ASAP7_75t_L g16285 ( 
.A(n_15755),
.Y(n_16285)
);

AND2x2_ASAP7_75t_L g16286 ( 
.A(n_16031),
.B(n_15415),
.Y(n_16286)
);

NOR2xp33_ASAP7_75t_SL g16287 ( 
.A(n_15690),
.B(n_15482),
.Y(n_16287)
);

OAI22xp5_ASAP7_75t_L g16288 ( 
.A1(n_15578),
.A2(n_15528),
.B1(n_15048),
.B2(n_15249),
.Y(n_16288)
);

AOI221x1_ASAP7_75t_SL g16289 ( 
.A1(n_15722),
.A2(n_16062),
.B1(n_15665),
.B2(n_15608),
.C(n_15745),
.Y(n_16289)
);

INVx1_ASAP7_75t_L g16290 ( 
.A(n_15759),
.Y(n_16290)
);

A2O1A1Ixp33_ASAP7_75t_SL g16291 ( 
.A1(n_15772),
.A2(n_15254),
.B(n_14925),
.C(n_15384),
.Y(n_16291)
);

NAND2xp5_ASAP7_75t_L g16292 ( 
.A(n_15630),
.B(n_2109),
.Y(n_16292)
);

OR2x2_ASAP7_75t_L g16293 ( 
.A(n_15592),
.B(n_2110),
.Y(n_16293)
);

AND2x2_ASAP7_75t_L g16294 ( 
.A(n_15600),
.B(n_14933),
.Y(n_16294)
);

A2O1A1Ixp33_ASAP7_75t_L g16295 ( 
.A1(n_15700),
.A2(n_15384),
.B(n_14933),
.C(n_2113),
.Y(n_16295)
);

NAND2xp5_ASAP7_75t_L g16296 ( 
.A(n_15729),
.B(n_2111),
.Y(n_16296)
);

INVxp67_ASAP7_75t_SL g16297 ( 
.A(n_15678),
.Y(n_16297)
);

INVx2_ASAP7_75t_SL g16298 ( 
.A(n_15960),
.Y(n_16298)
);

A2O1A1Ixp33_ASAP7_75t_L g16299 ( 
.A1(n_15971),
.A2(n_2114),
.B(n_2111),
.C(n_2112),
.Y(n_16299)
);

AND2x2_ASAP7_75t_L g16300 ( 
.A(n_15899),
.B(n_2112),
.Y(n_16300)
);

CKINVDCx16_ASAP7_75t_R g16301 ( 
.A(n_15719),
.Y(n_16301)
);

NAND3xp33_ASAP7_75t_L g16302 ( 
.A(n_15901),
.B(n_2114),
.C(n_2115),
.Y(n_16302)
);

OR2x2_ASAP7_75t_L g16303 ( 
.A(n_15870),
.B(n_2115),
.Y(n_16303)
);

INVx1_ASAP7_75t_L g16304 ( 
.A(n_15766),
.Y(n_16304)
);

AND2x2_ASAP7_75t_L g16305 ( 
.A(n_15910),
.B(n_2116),
.Y(n_16305)
);

AOI21xp5_ASAP7_75t_L g16306 ( 
.A1(n_16030),
.A2(n_2116),
.B(n_2117),
.Y(n_16306)
);

OR2x2_ASAP7_75t_L g16307 ( 
.A(n_15696),
.B(n_2117),
.Y(n_16307)
);

NAND2xp5_ASAP7_75t_L g16308 ( 
.A(n_15830),
.B(n_2118),
.Y(n_16308)
);

HB1xp67_ASAP7_75t_L g16309 ( 
.A(n_15996),
.Y(n_16309)
);

AND2x2_ASAP7_75t_L g16310 ( 
.A(n_15912),
.B(n_2118),
.Y(n_16310)
);

INVx1_ASAP7_75t_L g16311 ( 
.A(n_15865),
.Y(n_16311)
);

NAND2xp5_ASAP7_75t_L g16312 ( 
.A(n_15882),
.B(n_2119),
.Y(n_16312)
);

NOR2xp67_ASAP7_75t_L g16313 ( 
.A(n_15606),
.B(n_2119),
.Y(n_16313)
);

BUFx4_ASAP7_75t_R g16314 ( 
.A(n_15792),
.Y(n_16314)
);

A2O1A1Ixp33_ASAP7_75t_L g16315 ( 
.A1(n_15758),
.A2(n_16010),
.B(n_15670),
.C(n_16023),
.Y(n_16315)
);

INVx1_ASAP7_75t_L g16316 ( 
.A(n_15875),
.Y(n_16316)
);

A2O1A1Ixp33_ASAP7_75t_L g16317 ( 
.A1(n_16017),
.A2(n_2122),
.B(n_2120),
.C(n_2121),
.Y(n_16317)
);

HB1xp67_ASAP7_75t_L g16318 ( 
.A(n_15998),
.Y(n_16318)
);

A2O1A1Ixp33_ASAP7_75t_L g16319 ( 
.A1(n_16003),
.A2(n_2122),
.B(n_2120),
.C(n_2121),
.Y(n_16319)
);

OR2x2_ASAP7_75t_L g16320 ( 
.A(n_15697),
.B(n_15640),
.Y(n_16320)
);

NAND2xp5_ASAP7_75t_L g16321 ( 
.A(n_15658),
.B(n_15675),
.Y(n_16321)
);

NOR2xp67_ASAP7_75t_L g16322 ( 
.A(n_15717),
.B(n_2123),
.Y(n_16322)
);

BUFx3_ASAP7_75t_L g16323 ( 
.A(n_16036),
.Y(n_16323)
);

O2A1O1Ixp5_ASAP7_75t_L g16324 ( 
.A1(n_15653),
.A2(n_2125),
.B(n_2123),
.C(n_2124),
.Y(n_16324)
);

O2A1O1Ixp5_ASAP7_75t_L g16325 ( 
.A1(n_15978),
.A2(n_2127),
.B(n_2125),
.C(n_2126),
.Y(n_16325)
);

INVx2_ASAP7_75t_L g16326 ( 
.A(n_15705),
.Y(n_16326)
);

NAND2xp5_ASAP7_75t_L g16327 ( 
.A(n_15963),
.B(n_2126),
.Y(n_16327)
);

INVx1_ASAP7_75t_L g16328 ( 
.A(n_16049),
.Y(n_16328)
);

CKINVDCx5p33_ASAP7_75t_R g16329 ( 
.A(n_15597),
.Y(n_16329)
);

BUFx4f_ASAP7_75t_SL g16330 ( 
.A(n_16069),
.Y(n_16330)
);

NAND2xp5_ASAP7_75t_L g16331 ( 
.A(n_15605),
.B(n_2127),
.Y(n_16331)
);

AND2x4_ASAP7_75t_SL g16332 ( 
.A(n_15726),
.B(n_2128),
.Y(n_16332)
);

AND2x4_ASAP7_75t_L g16333 ( 
.A(n_16068),
.B(n_2129),
.Y(n_16333)
);

AND2x2_ASAP7_75t_L g16334 ( 
.A(n_15918),
.B(n_2129),
.Y(n_16334)
);

AND2x2_ASAP7_75t_L g16335 ( 
.A(n_15721),
.B(n_2130),
.Y(n_16335)
);

INVx1_ASAP7_75t_L g16336 ( 
.A(n_16060),
.Y(n_16336)
);

INVx1_ASAP7_75t_L g16337 ( 
.A(n_16064),
.Y(n_16337)
);

A2O1A1Ixp33_ASAP7_75t_L g16338 ( 
.A1(n_15950),
.A2(n_2132),
.B(n_2130),
.C(n_2131),
.Y(n_16338)
);

O2A1O1Ixp5_ASAP7_75t_L g16339 ( 
.A1(n_15823),
.A2(n_2133),
.B(n_2131),
.C(n_2132),
.Y(n_16339)
);

CKINVDCx20_ASAP7_75t_R g16340 ( 
.A(n_15707),
.Y(n_16340)
);

NAND2xp5_ASAP7_75t_L g16341 ( 
.A(n_15651),
.B(n_2133),
.Y(n_16341)
);

AND2x2_ASAP7_75t_L g16342 ( 
.A(n_15712),
.B(n_2134),
.Y(n_16342)
);

INVx2_ASAP7_75t_L g16343 ( 
.A(n_15716),
.Y(n_16343)
);

AND2x2_ASAP7_75t_L g16344 ( 
.A(n_16052),
.B(n_2134),
.Y(n_16344)
);

INVxp67_ASAP7_75t_L g16345 ( 
.A(n_15983),
.Y(n_16345)
);

INVx1_ASAP7_75t_L g16346 ( 
.A(n_16067),
.Y(n_16346)
);

NAND2xp5_ASAP7_75t_L g16347 ( 
.A(n_16073),
.B(n_2135),
.Y(n_16347)
);

AND2x2_ASAP7_75t_L g16348 ( 
.A(n_16048),
.B(n_2135),
.Y(n_16348)
);

OAI22xp5_ASAP7_75t_L g16349 ( 
.A1(n_15710),
.A2(n_2138),
.B1(n_2136),
.B2(n_2137),
.Y(n_16349)
);

A2O1A1Ixp33_ASAP7_75t_L g16350 ( 
.A1(n_16013),
.A2(n_2138),
.B(n_2136),
.C(n_2137),
.Y(n_16350)
);

AND2x4_ASAP7_75t_L g16351 ( 
.A(n_15976),
.B(n_2139),
.Y(n_16351)
);

A2O1A1Ixp33_ASAP7_75t_L g16352 ( 
.A1(n_16050),
.A2(n_2141),
.B(n_2139),
.C(n_2140),
.Y(n_16352)
);

O2A1O1Ixp33_ASAP7_75t_L g16353 ( 
.A1(n_16071),
.A2(n_2142),
.B(n_2140),
.C(n_2141),
.Y(n_16353)
);

A2O1A1Ixp33_ASAP7_75t_L g16354 ( 
.A1(n_15883),
.A2(n_16014),
.B(n_16032),
.C(n_15984),
.Y(n_16354)
);

HB1xp67_ASAP7_75t_L g16355 ( 
.A(n_15939),
.Y(n_16355)
);

HB1xp67_ASAP7_75t_L g16356 ( 
.A(n_15945),
.Y(n_16356)
);

INVx1_ASAP7_75t_L g16357 ( 
.A(n_16074),
.Y(n_16357)
);

INVxp67_ASAP7_75t_L g16358 ( 
.A(n_15992),
.Y(n_16358)
);

AOI21xp5_ASAP7_75t_L g16359 ( 
.A1(n_15986),
.A2(n_16079),
.B(n_15863),
.Y(n_16359)
);

INVx2_ASAP7_75t_L g16360 ( 
.A(n_15720),
.Y(n_16360)
);

NAND2xp5_ASAP7_75t_L g16361 ( 
.A(n_16075),
.B(n_2142),
.Y(n_16361)
);

OR2x2_ASAP7_75t_L g16362 ( 
.A(n_15704),
.B(n_15738),
.Y(n_16362)
);

AOI21xp5_ASAP7_75t_L g16363 ( 
.A1(n_15776),
.A2(n_2143),
.B(n_2144),
.Y(n_16363)
);

BUFx4_ASAP7_75t_R g16364 ( 
.A(n_15586),
.Y(n_16364)
);

NAND2xp5_ASAP7_75t_L g16365 ( 
.A(n_15952),
.B(n_2145),
.Y(n_16365)
);

CKINVDCx6p67_ASAP7_75t_R g16366 ( 
.A(n_15966),
.Y(n_16366)
);

AOI21xp5_ASAP7_75t_L g16367 ( 
.A1(n_15884),
.A2(n_2145),
.B(n_2146),
.Y(n_16367)
);

AND2x4_ASAP7_75t_L g16368 ( 
.A(n_16039),
.B(n_2146),
.Y(n_16368)
);

AND2x2_ASAP7_75t_L g16369 ( 
.A(n_15991),
.B(n_2147),
.Y(n_16369)
);

BUFx6f_ASAP7_75t_L g16370 ( 
.A(n_15842),
.Y(n_16370)
);

INVx1_ASAP7_75t_L g16371 ( 
.A(n_15962),
.Y(n_16371)
);

INVx1_ASAP7_75t_L g16372 ( 
.A(n_15969),
.Y(n_16372)
);

INVx1_ASAP7_75t_L g16373 ( 
.A(n_15974),
.Y(n_16373)
);

INVx2_ASAP7_75t_L g16374 ( 
.A(n_15624),
.Y(n_16374)
);

A2O1A1Ixp33_ASAP7_75t_SL g16375 ( 
.A1(n_15793),
.A2(n_2149),
.B(n_2147),
.C(n_2148),
.Y(n_16375)
);

AND2x4_ASAP7_75t_L g16376 ( 
.A(n_15679),
.B(n_2148),
.Y(n_16376)
);

AOI221x1_ASAP7_75t_L g16377 ( 
.A1(n_15767),
.A2(n_2152),
.B1(n_2150),
.B2(n_2151),
.C(n_2153),
.Y(n_16377)
);

AND2x2_ASAP7_75t_L g16378 ( 
.A(n_15695),
.B(n_2150),
.Y(n_16378)
);

NAND2xp5_ASAP7_75t_L g16379 ( 
.A(n_16016),
.B(n_2151),
.Y(n_16379)
);

NAND2xp5_ASAP7_75t_L g16380 ( 
.A(n_16021),
.B(n_2152),
.Y(n_16380)
);

AND2x2_ASAP7_75t_L g16381 ( 
.A(n_15673),
.B(n_2153),
.Y(n_16381)
);

INVx8_ASAP7_75t_L g16382 ( 
.A(n_15966),
.Y(n_16382)
);

OAI22xp5_ASAP7_75t_SL g16383 ( 
.A1(n_15732),
.A2(n_2157),
.B1(n_2155),
.B2(n_2156),
.Y(n_16383)
);

AND2x2_ASAP7_75t_L g16384 ( 
.A(n_15728),
.B(n_2155),
.Y(n_16384)
);

NAND2xp5_ASAP7_75t_L g16385 ( 
.A(n_16022),
.B(n_2156),
.Y(n_16385)
);

NOR2xp33_ASAP7_75t_L g16386 ( 
.A(n_15644),
.B(n_2157),
.Y(n_16386)
);

INVx2_ASAP7_75t_L g16387 ( 
.A(n_15652),
.Y(n_16387)
);

BUFx12f_ASAP7_75t_L g16388 ( 
.A(n_15988),
.Y(n_16388)
);

NAND2xp5_ASAP7_75t_L g16389 ( 
.A(n_16047),
.B(n_2158),
.Y(n_16389)
);

AND2x4_ASAP7_75t_L g16390 ( 
.A(n_16055),
.B(n_2159),
.Y(n_16390)
);

AND2x2_ASAP7_75t_L g16391 ( 
.A(n_15956),
.B(n_16066),
.Y(n_16391)
);

INVx3_ASAP7_75t_L g16392 ( 
.A(n_15842),
.Y(n_16392)
);

AND2x2_ASAP7_75t_L g16393 ( 
.A(n_15647),
.B(n_2159),
.Y(n_16393)
);

AOI21xp5_ASAP7_75t_L g16394 ( 
.A1(n_15814),
.A2(n_2160),
.B(n_2161),
.Y(n_16394)
);

OAI22xp5_ASAP7_75t_L g16395 ( 
.A1(n_15801),
.A2(n_2164),
.B1(n_2161),
.B2(n_2163),
.Y(n_16395)
);

AND2x2_ASAP7_75t_L g16396 ( 
.A(n_15668),
.B(n_2163),
.Y(n_16396)
);

AND2x2_ASAP7_75t_L g16397 ( 
.A(n_15687),
.B(n_2164),
.Y(n_16397)
);

A2O1A1Ixp33_ASAP7_75t_L g16398 ( 
.A1(n_15781),
.A2(n_16037),
.B(n_15993),
.C(n_15979),
.Y(n_16398)
);

A2O1A1Ixp33_ASAP7_75t_L g16399 ( 
.A1(n_15909),
.A2(n_2167),
.B(n_2165),
.C(n_2166),
.Y(n_16399)
);

NAND2xp5_ASAP7_75t_L g16400 ( 
.A(n_15778),
.B(n_2165),
.Y(n_16400)
);

INVx1_ASAP7_75t_L g16401 ( 
.A(n_15779),
.Y(n_16401)
);

INVx2_ASAP7_75t_L g16402 ( 
.A(n_15847),
.Y(n_16402)
);

INVx1_ASAP7_75t_L g16403 ( 
.A(n_15782),
.Y(n_16403)
);

BUFx3_ASAP7_75t_L g16404 ( 
.A(n_16070),
.Y(n_16404)
);

A2O1A1Ixp33_ASAP7_75t_L g16405 ( 
.A1(n_15677),
.A2(n_2168),
.B(n_2166),
.C(n_2167),
.Y(n_16405)
);

OR2x2_ASAP7_75t_L g16406 ( 
.A(n_15798),
.B(n_2168),
.Y(n_16406)
);

AOI21xp5_ASAP7_75t_SL g16407 ( 
.A1(n_15819),
.A2(n_2169),
.B(n_2170),
.Y(n_16407)
);

NAND2xp5_ASAP7_75t_SL g16408 ( 
.A(n_15655),
.B(n_2169),
.Y(n_16408)
);

NOR2xp33_ASAP7_75t_L g16409 ( 
.A(n_15723),
.B(n_2171),
.Y(n_16409)
);

AOI21x1_ASAP7_75t_SL g16410 ( 
.A1(n_15741),
.A2(n_2171),
.B(n_2172),
.Y(n_16410)
);

AOI21xp5_ASAP7_75t_L g16411 ( 
.A1(n_15593),
.A2(n_2172),
.B(n_2173),
.Y(n_16411)
);

NOR2xp33_ASAP7_75t_L g16412 ( 
.A(n_15736),
.B(n_2174),
.Y(n_16412)
);

INVx2_ASAP7_75t_L g16413 ( 
.A(n_15825),
.Y(n_16413)
);

INVx2_ASAP7_75t_L g16414 ( 
.A(n_15573),
.Y(n_16414)
);

INVx1_ASAP7_75t_L g16415 ( 
.A(n_15765),
.Y(n_16415)
);

NAND2xp5_ASAP7_75t_SL g16416 ( 
.A(n_15615),
.B(n_2175),
.Y(n_16416)
);

HB1xp67_ASAP7_75t_L g16417 ( 
.A(n_15769),
.Y(n_16417)
);

NAND2xp5_ASAP7_75t_L g16418 ( 
.A(n_15744),
.B(n_2175),
.Y(n_16418)
);

AOI22xp5_ASAP7_75t_L g16419 ( 
.A1(n_15954),
.A2(n_2178),
.B1(n_2176),
.B2(n_2177),
.Y(n_16419)
);

INVx1_ASAP7_75t_L g16420 ( 
.A(n_15580),
.Y(n_16420)
);

CKINVDCx5p33_ASAP7_75t_R g16421 ( 
.A(n_15751),
.Y(n_16421)
);

INVx1_ASAP7_75t_L g16422 ( 
.A(n_15859),
.Y(n_16422)
);

O2A1O1Ixp33_ASAP7_75t_L g16423 ( 
.A1(n_15968),
.A2(n_2178),
.B(n_2176),
.C(n_2177),
.Y(n_16423)
);

INVx2_ASAP7_75t_L g16424 ( 
.A(n_15649),
.Y(n_16424)
);

OA21x2_ASAP7_75t_L g16425 ( 
.A1(n_15951),
.A2(n_2179),
.B(n_2180),
.Y(n_16425)
);

AND2x2_ASAP7_75t_L g16426 ( 
.A(n_15639),
.B(n_2179),
.Y(n_16426)
);

AND2x2_ASAP7_75t_L g16427 ( 
.A(n_15851),
.B(n_2180),
.Y(n_16427)
);

INVx1_ASAP7_75t_L g16428 ( 
.A(n_15841),
.Y(n_16428)
);

NAND2xp5_ASAP7_75t_L g16429 ( 
.A(n_15764),
.B(n_2181),
.Y(n_16429)
);

INVx2_ASAP7_75t_SL g16430 ( 
.A(n_15726),
.Y(n_16430)
);

OA21x2_ASAP7_75t_L g16431 ( 
.A1(n_15791),
.A2(n_2181),
.B(n_2182),
.Y(n_16431)
);

INVx2_ASAP7_75t_L g16432 ( 
.A(n_16061),
.Y(n_16432)
);

AND2x2_ASAP7_75t_L g16433 ( 
.A(n_15888),
.B(n_2182),
.Y(n_16433)
);

BUFx3_ASAP7_75t_L g16434 ( 
.A(n_15888),
.Y(n_16434)
);

INVxp33_ASAP7_75t_L g16435 ( 
.A(n_15601),
.Y(n_16435)
);

OR2x2_ASAP7_75t_L g16436 ( 
.A(n_15896),
.B(n_2183),
.Y(n_16436)
);

NOR2x1_ASAP7_75t_SL g16437 ( 
.A(n_15747),
.B(n_2184),
.Y(n_16437)
);

BUFx2_ASAP7_75t_L g16438 ( 
.A(n_15911),
.Y(n_16438)
);

AND2x2_ASAP7_75t_L g16439 ( 
.A(n_16009),
.B(n_2184),
.Y(n_16439)
);

NOR2xp33_ASAP7_75t_L g16440 ( 
.A(n_15674),
.B(n_2185),
.Y(n_16440)
);

O2A1O1Ixp33_ASAP7_75t_L g16441 ( 
.A1(n_16015),
.A2(n_2187),
.B(n_2185),
.C(n_2186),
.Y(n_16441)
);

NAND2xp5_ASAP7_75t_L g16442 ( 
.A(n_15869),
.B(n_2186),
.Y(n_16442)
);

NAND2xp5_ASAP7_75t_L g16443 ( 
.A(n_15874),
.B(n_2187),
.Y(n_16443)
);

A2O1A1Ixp33_ASAP7_75t_L g16444 ( 
.A1(n_16059),
.A2(n_15921),
.B(n_16056),
.C(n_16027),
.Y(n_16444)
);

NOR2xp67_ASAP7_75t_L g16445 ( 
.A(n_15790),
.B(n_2188),
.Y(n_16445)
);

CKINVDCx5p33_ASAP7_75t_R g16446 ( 
.A(n_15805),
.Y(n_16446)
);

INVx1_ASAP7_75t_SL g16447 ( 
.A(n_15900),
.Y(n_16447)
);

INVx1_ASAP7_75t_L g16448 ( 
.A(n_15817),
.Y(n_16448)
);

INVx2_ASAP7_75t_L g16449 ( 
.A(n_16009),
.Y(n_16449)
);

NAND2xp5_ASAP7_75t_L g16450 ( 
.A(n_15787),
.B(n_2188),
.Y(n_16450)
);

AND2x2_ASAP7_75t_L g16451 ( 
.A(n_16018),
.B(n_2189),
.Y(n_16451)
);

INVx2_ASAP7_75t_L g16452 ( 
.A(n_16018),
.Y(n_16452)
);

NOR2xp33_ASAP7_75t_R g16453 ( 
.A(n_16029),
.B(n_2189),
.Y(n_16453)
);

INVx1_ASAP7_75t_L g16454 ( 
.A(n_15796),
.Y(n_16454)
);

INVx2_ASAP7_75t_L g16455 ( 
.A(n_16043),
.Y(n_16455)
);

AND2x2_ASAP7_75t_L g16456 ( 
.A(n_16043),
.B(n_2190),
.Y(n_16456)
);

INVx2_ASAP7_75t_L g16457 ( 
.A(n_15771),
.Y(n_16457)
);

OR2x2_ASAP7_75t_L g16458 ( 
.A(n_15943),
.B(n_2190),
.Y(n_16458)
);

AND2x4_ASAP7_75t_SL g16459 ( 
.A(n_15853),
.B(n_15866),
.Y(n_16459)
);

CKINVDCx6p67_ASAP7_75t_R g16460 ( 
.A(n_15989),
.Y(n_16460)
);

INVx2_ASAP7_75t_L g16461 ( 
.A(n_16083),
.Y(n_16461)
);

NAND2xp5_ASAP7_75t_L g16462 ( 
.A(n_15822),
.B(n_2191),
.Y(n_16462)
);

NAND2x1p5_ASAP7_75t_L g16463 ( 
.A(n_15881),
.B(n_2191),
.Y(n_16463)
);

AOI21x1_ASAP7_75t_SL g16464 ( 
.A1(n_15761),
.A2(n_2192),
.B(n_2193),
.Y(n_16464)
);

NAND2xp5_ASAP7_75t_L g16465 ( 
.A(n_15840),
.B(n_15856),
.Y(n_16465)
);

BUFx12f_ASAP7_75t_L g16466 ( 
.A(n_16033),
.Y(n_16466)
);

OR2x6_ASAP7_75t_L g16467 ( 
.A(n_15821),
.B(n_2192),
.Y(n_16467)
);

NOR2xp33_ASAP7_75t_L g16468 ( 
.A(n_16081),
.B(n_2193),
.Y(n_16468)
);

OA21x2_ASAP7_75t_L g16469 ( 
.A1(n_15789),
.A2(n_2194),
.B(n_2195),
.Y(n_16469)
);

OR2x2_ASAP7_75t_L g16470 ( 
.A(n_16028),
.B(n_2194),
.Y(n_16470)
);

A2O1A1Ixp33_ASAP7_75t_L g16471 ( 
.A1(n_15895),
.A2(n_2197),
.B(n_2195),
.C(n_2196),
.Y(n_16471)
);

AOI21xp5_ASAP7_75t_L g16472 ( 
.A1(n_15795),
.A2(n_2196),
.B(n_2197),
.Y(n_16472)
);

INVx2_ASAP7_75t_L g16473 ( 
.A(n_15768),
.Y(n_16473)
);

INVx1_ASAP7_75t_L g16474 ( 
.A(n_15839),
.Y(n_16474)
);

HB1xp67_ASAP7_75t_L g16475 ( 
.A(n_15982),
.Y(n_16475)
);

OR2x2_ASAP7_75t_L g16476 ( 
.A(n_15916),
.B(n_2198),
.Y(n_16476)
);

AND2x2_ASAP7_75t_L g16477 ( 
.A(n_15661),
.B(n_2198),
.Y(n_16477)
);

BUFx3_ASAP7_75t_L g16478 ( 
.A(n_15894),
.Y(n_16478)
);

INVx2_ASAP7_75t_L g16479 ( 
.A(n_15834),
.Y(n_16479)
);

HB1xp67_ASAP7_75t_L g16480 ( 
.A(n_16002),
.Y(n_16480)
);

OAI22xp5_ASAP7_75t_L g16481 ( 
.A1(n_16046),
.A2(n_2201),
.B1(n_2199),
.B2(n_2200),
.Y(n_16481)
);

A2O1A1Ixp33_ASAP7_75t_SL g16482 ( 
.A1(n_15828),
.A2(n_2201),
.B(n_2199),
.C(n_2200),
.Y(n_16482)
);

INVx1_ASAP7_75t_L g16483 ( 
.A(n_15852),
.Y(n_16483)
);

AND2x2_ASAP7_75t_L g16484 ( 
.A(n_15730),
.B(n_2202),
.Y(n_16484)
);

INVx2_ASAP7_75t_L g16485 ( 
.A(n_15953),
.Y(n_16485)
);

HB1xp67_ASAP7_75t_L g16486 ( 
.A(n_15846),
.Y(n_16486)
);

NOR2xp33_ASAP7_75t_R g16487 ( 
.A(n_15571),
.B(n_2202),
.Y(n_16487)
);

INVx1_ASAP7_75t_L g16488 ( 
.A(n_15923),
.Y(n_16488)
);

AND2x2_ASAP7_75t_L g16489 ( 
.A(n_15994),
.B(n_2203),
.Y(n_16489)
);

OR2x6_ASAP7_75t_SL g16490 ( 
.A(n_15582),
.B(n_2203),
.Y(n_16490)
);

OAI22xp5_ASAP7_75t_L g16491 ( 
.A1(n_16053),
.A2(n_2206),
.B1(n_2204),
.B2(n_2205),
.Y(n_16491)
);

INVx1_ASAP7_75t_L g16492 ( 
.A(n_15973),
.Y(n_16492)
);

HB1xp67_ASAP7_75t_L g16493 ( 
.A(n_15977),
.Y(n_16493)
);

INVx1_ASAP7_75t_L g16494 ( 
.A(n_15808),
.Y(n_16494)
);

NOR2xp33_ASAP7_75t_L g16495 ( 
.A(n_15915),
.B(n_15585),
.Y(n_16495)
);

NAND2xp5_ASAP7_75t_L g16496 ( 
.A(n_15627),
.B(n_2204),
.Y(n_16496)
);

AOI21xp5_ASAP7_75t_L g16497 ( 
.A1(n_16084),
.A2(n_2205),
.B(n_2206),
.Y(n_16497)
);

INVx1_ASAP7_75t_L g16498 ( 
.A(n_15816),
.Y(n_16498)
);

NAND2xp5_ASAP7_75t_L g16499 ( 
.A(n_16057),
.B(n_2207),
.Y(n_16499)
);

AOI21xp5_ASAP7_75t_L g16500 ( 
.A1(n_15701),
.A2(n_2208),
.B(n_2209),
.Y(n_16500)
);

NAND2xp5_ASAP7_75t_L g16501 ( 
.A(n_15571),
.B(n_2208),
.Y(n_16501)
);

AND2x2_ASAP7_75t_L g16502 ( 
.A(n_15972),
.B(n_2209),
.Y(n_16502)
);

OR2x2_ASAP7_75t_L g16503 ( 
.A(n_16065),
.B(n_2210),
.Y(n_16503)
);

A2O1A1Ixp33_ASAP7_75t_L g16504 ( 
.A1(n_15753),
.A2(n_2213),
.B(n_2211),
.C(n_2212),
.Y(n_16504)
);

NAND2xp5_ASAP7_75t_L g16505 ( 
.A(n_15571),
.B(n_2211),
.Y(n_16505)
);

AND2x2_ASAP7_75t_L g16506 ( 
.A(n_15959),
.B(n_2212),
.Y(n_16506)
);

AND2x4_ASAP7_75t_L g16507 ( 
.A(n_16078),
.B(n_2213),
.Y(n_16507)
);

AOI21xp5_ASAP7_75t_SL g16508 ( 
.A1(n_16045),
.A2(n_2214),
.B(n_2215),
.Y(n_16508)
);

AND2x2_ASAP7_75t_L g16509 ( 
.A(n_15844),
.B(n_15967),
.Y(n_16509)
);

OR2x2_ASAP7_75t_L g16510 ( 
.A(n_16077),
.B(n_2214),
.Y(n_16510)
);

BUFx4_ASAP7_75t_R g16511 ( 
.A(n_16004),
.Y(n_16511)
);

OAI22xp5_ASAP7_75t_L g16512 ( 
.A1(n_15917),
.A2(n_2219),
.B1(n_2216),
.B2(n_2218),
.Y(n_16512)
);

AND2x2_ASAP7_75t_L g16513 ( 
.A(n_16058),
.B(n_15961),
.Y(n_16513)
);

HB1xp67_ASAP7_75t_L g16514 ( 
.A(n_15965),
.Y(n_16514)
);

INVx1_ASAP7_75t_L g16515 ( 
.A(n_15879),
.Y(n_16515)
);

A2O1A1Ixp33_ASAP7_75t_SL g16516 ( 
.A1(n_15848),
.A2(n_2219),
.B(n_2216),
.C(n_2218),
.Y(n_16516)
);

OAI22xp5_ASAP7_75t_L g16517 ( 
.A1(n_16042),
.A2(n_2222),
.B1(n_2220),
.B2(n_2221),
.Y(n_16517)
);

O2A1O1Ixp33_ASAP7_75t_L g16518 ( 
.A1(n_15775),
.A2(n_2223),
.B(n_2220),
.C(n_2222),
.Y(n_16518)
);

INVx2_ASAP7_75t_L g16519 ( 
.A(n_15872),
.Y(n_16519)
);

AOI21xp5_ASAP7_75t_L g16520 ( 
.A1(n_16024),
.A2(n_2223),
.B(n_2224),
.Y(n_16520)
);

HB1xp67_ASAP7_75t_L g16521 ( 
.A(n_15748),
.Y(n_16521)
);

INVx2_ASAP7_75t_L g16522 ( 
.A(n_16314),
.Y(n_16522)
);

OAI21x1_ASAP7_75t_L g16523 ( 
.A1(n_16138),
.A2(n_15810),
.B(n_15760),
.Y(n_16523)
);

INVx1_ASAP7_75t_L g16524 ( 
.A(n_16355),
.Y(n_16524)
);

AND2x2_ASAP7_75t_L g16525 ( 
.A(n_16301),
.B(n_15686),
.Y(n_16525)
);

INVx2_ASAP7_75t_L g16526 ( 
.A(n_16404),
.Y(n_16526)
);

HB1xp67_ASAP7_75t_L g16527 ( 
.A(n_16136),
.Y(n_16527)
);

BUFx3_ASAP7_75t_L g16528 ( 
.A(n_16195),
.Y(n_16528)
);

BUFx3_ASAP7_75t_L g16529 ( 
.A(n_16200),
.Y(n_16529)
);

CKINVDCx6p67_ASAP7_75t_R g16530 ( 
.A(n_16278),
.Y(n_16530)
);

OA21x2_ASAP7_75t_L g16531 ( 
.A1(n_16109),
.A2(n_15886),
.B(n_15885),
.Y(n_16531)
);

INVx1_ASAP7_75t_L g16532 ( 
.A(n_16356),
.Y(n_16532)
);

OAI21x1_ASAP7_75t_L g16533 ( 
.A1(n_16096),
.A2(n_15763),
.B(n_15750),
.Y(n_16533)
);

OAI21x1_ASAP7_75t_L g16534 ( 
.A1(n_16160),
.A2(n_15770),
.B(n_15891),
.Y(n_16534)
);

INVx2_ASAP7_75t_L g16535 ( 
.A(n_16438),
.Y(n_16535)
);

INVx1_ASAP7_75t_L g16536 ( 
.A(n_16309),
.Y(n_16536)
);

CKINVDCx11_ASAP7_75t_R g16537 ( 
.A(n_16232),
.Y(n_16537)
);

NAND2xp5_ASAP7_75t_L g16538 ( 
.A(n_16412),
.B(n_16001),
.Y(n_16538)
);

INVx1_ASAP7_75t_L g16539 ( 
.A(n_16318),
.Y(n_16539)
);

INVx1_ASAP7_75t_L g16540 ( 
.A(n_16328),
.Y(n_16540)
);

INVx2_ASAP7_75t_L g16541 ( 
.A(n_16165),
.Y(n_16541)
);

AO21x2_ASAP7_75t_L g16542 ( 
.A1(n_16331),
.A2(n_16007),
.B(n_15958),
.Y(n_16542)
);

AND2x2_ASAP7_75t_L g16543 ( 
.A(n_16273),
.B(n_16035),
.Y(n_16543)
);

OR2x2_ASAP7_75t_L g16544 ( 
.A(n_16095),
.B(n_16108),
.Y(n_16544)
);

INVx1_ASAP7_75t_L g16545 ( 
.A(n_16336),
.Y(n_16545)
);

AND2x2_ASAP7_75t_L g16546 ( 
.A(n_16140),
.B(n_16041),
.Y(n_16546)
);

INVx2_ASAP7_75t_L g16547 ( 
.A(n_16197),
.Y(n_16547)
);

INVx1_ASAP7_75t_L g16548 ( 
.A(n_16337),
.Y(n_16548)
);

HB1xp67_ASAP7_75t_L g16549 ( 
.A(n_16191),
.Y(n_16549)
);

BUFx12f_ASAP7_75t_L g16550 ( 
.A(n_16169),
.Y(n_16550)
);

HB1xp67_ASAP7_75t_L g16551 ( 
.A(n_16103),
.Y(n_16551)
);

INVx3_ASAP7_75t_L g16552 ( 
.A(n_16086),
.Y(n_16552)
);

INVx1_ASAP7_75t_L g16553 ( 
.A(n_16346),
.Y(n_16553)
);

INVx2_ASAP7_75t_L g16554 ( 
.A(n_16430),
.Y(n_16554)
);

NAND2x1p5_ASAP7_75t_L g16555 ( 
.A(n_16174),
.B(n_16006),
.Y(n_16555)
);

NAND2xp5_ASAP7_75t_L g16556 ( 
.A(n_16230),
.B(n_15632),
.Y(n_16556)
);

INVx1_ASAP7_75t_L g16557 ( 
.A(n_16357),
.Y(n_16557)
);

INVx2_ASAP7_75t_L g16558 ( 
.A(n_16220),
.Y(n_16558)
);

CKINVDCx6p67_ASAP7_75t_R g16559 ( 
.A(n_16255),
.Y(n_16559)
);

INVx1_ASAP7_75t_L g16560 ( 
.A(n_16371),
.Y(n_16560)
);

INVx1_ASAP7_75t_L g16561 ( 
.A(n_16372),
.Y(n_16561)
);

HB1xp67_ASAP7_75t_L g16562 ( 
.A(n_16322),
.Y(n_16562)
);

BUFx3_ASAP7_75t_L g16563 ( 
.A(n_16340),
.Y(n_16563)
);

INVx1_ASAP7_75t_SL g16564 ( 
.A(n_16487),
.Y(n_16564)
);

INVxp67_ASAP7_75t_L g16565 ( 
.A(n_16090),
.Y(n_16565)
);

INVx1_ASAP7_75t_L g16566 ( 
.A(n_16373),
.Y(n_16566)
);

INVx2_ASAP7_75t_L g16567 ( 
.A(n_16277),
.Y(n_16567)
);

INVx1_ASAP7_75t_L g16568 ( 
.A(n_16091),
.Y(n_16568)
);

INVx1_ASAP7_75t_L g16569 ( 
.A(n_16101),
.Y(n_16569)
);

AND2x2_ASAP7_75t_L g16570 ( 
.A(n_16204),
.B(n_15785),
.Y(n_16570)
);

HB1xp67_ASAP7_75t_L g16571 ( 
.A(n_16133),
.Y(n_16571)
);

INVx5_ASAP7_75t_L g16572 ( 
.A(n_16382),
.Y(n_16572)
);

AO21x2_ASAP7_75t_L g16573 ( 
.A1(n_16183),
.A2(n_15873),
.B(n_16019),
.Y(n_16573)
);

INVx2_ASAP7_75t_L g16574 ( 
.A(n_16085),
.Y(n_16574)
);

INVx1_ASAP7_75t_L g16575 ( 
.A(n_16111),
.Y(n_16575)
);

AND2x2_ASAP7_75t_L g16576 ( 
.A(n_16118),
.B(n_15877),
.Y(n_16576)
);

INVx1_ASAP7_75t_L g16577 ( 
.A(n_16114),
.Y(n_16577)
);

INVx1_ASAP7_75t_L g16578 ( 
.A(n_16123),
.Y(n_16578)
);

HB1xp67_ASAP7_75t_L g16579 ( 
.A(n_16448),
.Y(n_16579)
);

INVx2_ASAP7_75t_L g16580 ( 
.A(n_16107),
.Y(n_16580)
);

AO21x2_ASAP7_75t_L g16581 ( 
.A1(n_16117),
.A2(n_16040),
.B(n_15762),
.Y(n_16581)
);

OR2x2_ASAP7_75t_L g16582 ( 
.A(n_16320),
.B(n_15740),
.Y(n_16582)
);

INVx1_ASAP7_75t_L g16583 ( 
.A(n_16128),
.Y(n_16583)
);

INVx2_ASAP7_75t_L g16584 ( 
.A(n_16298),
.Y(n_16584)
);

INVx1_ASAP7_75t_L g16585 ( 
.A(n_16132),
.Y(n_16585)
);

CKINVDCx5p33_ASAP7_75t_R g16586 ( 
.A(n_16106),
.Y(n_16586)
);

NAND2xp5_ASAP7_75t_L g16587 ( 
.A(n_16266),
.B(n_16271),
.Y(n_16587)
);

INVx1_ASAP7_75t_L g16588 ( 
.A(n_16146),
.Y(n_16588)
);

INVx4_ASAP7_75t_SL g16589 ( 
.A(n_16330),
.Y(n_16589)
);

OAI21x1_ASAP7_75t_L g16590 ( 
.A1(n_16150),
.A2(n_15835),
.B(n_15826),
.Y(n_16590)
);

INVx2_ASAP7_75t_L g16591 ( 
.A(n_16434),
.Y(n_16591)
);

INVx3_ASAP7_75t_L g16592 ( 
.A(n_16279),
.Y(n_16592)
);

NAND2xp5_ASAP7_75t_L g16593 ( 
.A(n_16345),
.B(n_15740),
.Y(n_16593)
);

INVx1_ASAP7_75t_L g16594 ( 
.A(n_16148),
.Y(n_16594)
);

AO21x2_ASAP7_75t_L g16595 ( 
.A1(n_16137),
.A2(n_15850),
.B(n_15809),
.Y(n_16595)
);

BUFx2_ASAP7_75t_L g16596 ( 
.A(n_16104),
.Y(n_16596)
);

INVx2_ASAP7_75t_L g16597 ( 
.A(n_16323),
.Y(n_16597)
);

INVx1_ASAP7_75t_L g16598 ( 
.A(n_16178),
.Y(n_16598)
);

NAND2xp5_ASAP7_75t_L g16599 ( 
.A(n_16358),
.B(n_15936),
.Y(n_16599)
);

AOI21x1_ASAP7_75t_L g16600 ( 
.A1(n_16099),
.A2(n_16122),
.B(n_16417),
.Y(n_16600)
);

INVx1_ASAP7_75t_L g16601 ( 
.A(n_16190),
.Y(n_16601)
);

HB1xp67_ASAP7_75t_L g16602 ( 
.A(n_16514),
.Y(n_16602)
);

AND2x2_ASAP7_75t_L g16603 ( 
.A(n_16203),
.B(n_16110),
.Y(n_16603)
);

NAND2xp5_ASAP7_75t_L g16604 ( 
.A(n_16432),
.B(n_15936),
.Y(n_16604)
);

INVx1_ASAP7_75t_L g16605 ( 
.A(n_16199),
.Y(n_16605)
);

NAND2xp5_ASAP7_75t_L g16606 ( 
.A(n_16286),
.B(n_15955),
.Y(n_16606)
);

INVx2_ASAP7_75t_L g16607 ( 
.A(n_16392),
.Y(n_16607)
);

INVx1_ASAP7_75t_L g16608 ( 
.A(n_16208),
.Y(n_16608)
);

OAI22xp5_ASAP7_75t_L g16609 ( 
.A1(n_16295),
.A2(n_15949),
.B1(n_15861),
.B2(n_16051),
.Y(n_16609)
);

OAI21xp5_ASAP7_75t_L g16610 ( 
.A1(n_16187),
.A2(n_16044),
.B(n_15897),
.Y(n_16610)
);

INVx2_ASAP7_75t_L g16611 ( 
.A(n_16370),
.Y(n_16611)
);

INVx1_ASAP7_75t_L g16612 ( 
.A(n_16223),
.Y(n_16612)
);

INVx1_ASAP7_75t_L g16613 ( 
.A(n_16238),
.Y(n_16613)
);

INVx2_ASAP7_75t_L g16614 ( 
.A(n_16370),
.Y(n_16614)
);

OAI221xp5_ASAP7_75t_L g16615 ( 
.A1(n_16289),
.A2(n_15955),
.B1(n_16051),
.B2(n_16054),
.C(n_15905),
.Y(n_16615)
);

BUFx6f_ASAP7_75t_L g16616 ( 
.A(n_16211),
.Y(n_16616)
);

HB1xp67_ASAP7_75t_SL g16617 ( 
.A(n_16349),
.Y(n_16617)
);

OAI21x1_ASAP7_75t_L g16618 ( 
.A1(n_16186),
.A2(n_15837),
.B(n_15858),
.Y(n_16618)
);

BUFx2_ASAP7_75t_L g16619 ( 
.A(n_16156),
.Y(n_16619)
);

INVx1_ASAP7_75t_L g16620 ( 
.A(n_16239),
.Y(n_16620)
);

INVx1_ASAP7_75t_L g16621 ( 
.A(n_16241),
.Y(n_16621)
);

OAI21x1_ASAP7_75t_L g16622 ( 
.A1(n_16143),
.A2(n_15868),
.B(n_15864),
.Y(n_16622)
);

OAI21x1_ASAP7_75t_L g16623 ( 
.A1(n_16088),
.A2(n_15906),
.B(n_15893),
.Y(n_16623)
);

INVx1_ASAP7_75t_L g16624 ( 
.A(n_16252),
.Y(n_16624)
);

INVx1_ASAP7_75t_L g16625 ( 
.A(n_16254),
.Y(n_16625)
);

AOI22xp33_ASAP7_75t_L g16626 ( 
.A1(n_16222),
.A2(n_15926),
.B1(n_15928),
.B2(n_15925),
.Y(n_16626)
);

AND2x4_ASAP7_75t_L g16627 ( 
.A(n_16176),
.B(n_15929),
.Y(n_16627)
);

INVx1_ASAP7_75t_L g16628 ( 
.A(n_16261),
.Y(n_16628)
);

NOR2xp33_ASAP7_75t_L g16629 ( 
.A(n_16216),
.B(n_15937),
.Y(n_16629)
);

INVx2_ASAP7_75t_L g16630 ( 
.A(n_16217),
.Y(n_16630)
);

HB1xp67_ASAP7_75t_L g16631 ( 
.A(n_16521),
.Y(n_16631)
);

CKINVDCx5p33_ASAP7_75t_R g16632 ( 
.A(n_16125),
.Y(n_16632)
);

INVx1_ASAP7_75t_L g16633 ( 
.A(n_16262),
.Y(n_16633)
);

NAND2xp5_ASAP7_75t_L g16634 ( 
.A(n_16498),
.B(n_15938),
.Y(n_16634)
);

INVx1_ASAP7_75t_L g16635 ( 
.A(n_16285),
.Y(n_16635)
);

INVx1_ASAP7_75t_L g16636 ( 
.A(n_16290),
.Y(n_16636)
);

INVx1_ASAP7_75t_L g16637 ( 
.A(n_16304),
.Y(n_16637)
);

INVx1_ASAP7_75t_L g16638 ( 
.A(n_16311),
.Y(n_16638)
);

OAI21x1_ASAP7_75t_L g16639 ( 
.A1(n_16413),
.A2(n_15942),
.B(n_15941),
.Y(n_16639)
);

INVx2_ASAP7_75t_L g16640 ( 
.A(n_16511),
.Y(n_16640)
);

INVx2_ASAP7_75t_L g16641 ( 
.A(n_16391),
.Y(n_16641)
);

INVx2_ASAP7_75t_L g16642 ( 
.A(n_16449),
.Y(n_16642)
);

AOI22xp33_ASAP7_75t_L g16643 ( 
.A1(n_16222),
.A2(n_16054),
.B1(n_2226),
.B2(n_2224),
.Y(n_16643)
);

AND2x2_ASAP7_75t_L g16644 ( 
.A(n_16131),
.B(n_2225),
.Y(n_16644)
);

INVx2_ASAP7_75t_L g16645 ( 
.A(n_16452),
.Y(n_16645)
);

AOI22xp33_ASAP7_75t_SL g16646 ( 
.A1(n_16364),
.A2(n_16288),
.B1(n_16283),
.B2(n_16153),
.Y(n_16646)
);

INVx2_ASAP7_75t_L g16647 ( 
.A(n_16455),
.Y(n_16647)
);

OR2x2_ASAP7_75t_L g16648 ( 
.A(n_16362),
.B(n_2225),
.Y(n_16648)
);

INVx2_ASAP7_75t_L g16649 ( 
.A(n_16382),
.Y(n_16649)
);

INVx2_ASAP7_75t_SL g16650 ( 
.A(n_16279),
.Y(n_16650)
);

BUFx2_ASAP7_75t_L g16651 ( 
.A(n_16156),
.Y(n_16651)
);

INVx2_ASAP7_75t_L g16652 ( 
.A(n_16154),
.Y(n_16652)
);

INVx1_ASAP7_75t_L g16653 ( 
.A(n_16316),
.Y(n_16653)
);

INVx1_ASAP7_75t_L g16654 ( 
.A(n_16428),
.Y(n_16654)
);

INVx1_ASAP7_75t_L g16655 ( 
.A(n_16401),
.Y(n_16655)
);

INVx1_ASAP7_75t_L g16656 ( 
.A(n_16403),
.Y(n_16656)
);

INVx1_ASAP7_75t_L g16657 ( 
.A(n_16420),
.Y(n_16657)
);

INVx1_ASAP7_75t_SL g16658 ( 
.A(n_16453),
.Y(n_16658)
);

HB1xp67_ASAP7_75t_L g16659 ( 
.A(n_16475),
.Y(n_16659)
);

AND2x4_ASAP7_75t_L g16660 ( 
.A(n_16188),
.B(n_2226),
.Y(n_16660)
);

INVx1_ASAP7_75t_L g16661 ( 
.A(n_16237),
.Y(n_16661)
);

HB1xp67_ASAP7_75t_L g16662 ( 
.A(n_16480),
.Y(n_16662)
);

BUFx3_ASAP7_75t_L g16663 ( 
.A(n_16161),
.Y(n_16663)
);

AO21x2_ASAP7_75t_L g16664 ( 
.A1(n_16297),
.A2(n_2227),
.B(n_2228),
.Y(n_16664)
);

INVx1_ASAP7_75t_L g16665 ( 
.A(n_16233),
.Y(n_16665)
);

INVx1_ASAP7_75t_L g16666 ( 
.A(n_16402),
.Y(n_16666)
);

CKINVDCx5p33_ASAP7_75t_R g16667 ( 
.A(n_16129),
.Y(n_16667)
);

BUFx3_ASAP7_75t_L g16668 ( 
.A(n_16466),
.Y(n_16668)
);

INVx2_ASAP7_75t_L g16669 ( 
.A(n_16151),
.Y(n_16669)
);

OAI21x1_ASAP7_75t_L g16670 ( 
.A1(n_16162),
.A2(n_2228),
.B(n_2229),
.Y(n_16670)
);

AOI22xp33_ASAP7_75t_L g16671 ( 
.A1(n_16243),
.A2(n_2231),
.B1(n_2229),
.B2(n_2230),
.Y(n_16671)
);

INVx3_ASAP7_75t_L g16672 ( 
.A(n_16215),
.Y(n_16672)
);

OR2x2_ASAP7_75t_L g16673 ( 
.A(n_16145),
.B(n_2231),
.Y(n_16673)
);

INVxp67_ASAP7_75t_L g16674 ( 
.A(n_16437),
.Y(n_16674)
);

INVx1_ASAP7_75t_L g16675 ( 
.A(n_16170),
.Y(n_16675)
);

AND2x4_ASAP7_75t_L g16676 ( 
.A(n_16092),
.B(n_2232),
.Y(n_16676)
);

AOI22xp33_ASAP7_75t_SL g16677 ( 
.A1(n_16087),
.A2(n_2234),
.B1(n_2232),
.B2(n_2233),
.Y(n_16677)
);

CKINVDCx20_ASAP7_75t_R g16678 ( 
.A(n_16460),
.Y(n_16678)
);

INVx2_ASAP7_75t_L g16679 ( 
.A(n_16151),
.Y(n_16679)
);

INVx1_ASAP7_75t_L g16680 ( 
.A(n_16100),
.Y(n_16680)
);

INVx1_ASAP7_75t_L g16681 ( 
.A(n_16422),
.Y(n_16681)
);

INVx2_ASAP7_75t_L g16682 ( 
.A(n_16253),
.Y(n_16682)
);

INVx1_ASAP7_75t_L g16683 ( 
.A(n_16374),
.Y(n_16683)
);

INVx1_ASAP7_75t_SL g16684 ( 
.A(n_16366),
.Y(n_16684)
);

INVx2_ASAP7_75t_L g16685 ( 
.A(n_16253),
.Y(n_16685)
);

AND2x4_ASAP7_75t_L g16686 ( 
.A(n_16275),
.B(n_2233),
.Y(n_16686)
);

BUFx2_ASAP7_75t_L g16687 ( 
.A(n_16388),
.Y(n_16687)
);

NAND2xp5_ASAP7_75t_L g16688 ( 
.A(n_16493),
.B(n_2234),
.Y(n_16688)
);

NOR2x1_ASAP7_75t_L g16689 ( 
.A(n_16407),
.B(n_2235),
.Y(n_16689)
);

INVx1_ASAP7_75t_L g16690 ( 
.A(n_16387),
.Y(n_16690)
);

AND2x2_ASAP7_75t_L g16691 ( 
.A(n_16127),
.B(n_2236),
.Y(n_16691)
);

BUFx2_ASAP7_75t_L g16692 ( 
.A(n_16229),
.Y(n_16692)
);

INVx2_ASAP7_75t_L g16693 ( 
.A(n_16272),
.Y(n_16693)
);

INVx1_ASAP7_75t_L g16694 ( 
.A(n_16175),
.Y(n_16694)
);

INVx3_ASAP7_75t_L g16695 ( 
.A(n_16272),
.Y(n_16695)
);

INVx1_ASAP7_75t_L g16696 ( 
.A(n_16414),
.Y(n_16696)
);

OA21x2_ASAP7_75t_L g16697 ( 
.A1(n_16201),
.A2(n_2236),
.B(n_2237),
.Y(n_16697)
);

NOR2xp67_ASAP7_75t_SL g16698 ( 
.A(n_16181),
.B(n_16166),
.Y(n_16698)
);

INVx1_ASAP7_75t_L g16699 ( 
.A(n_16214),
.Y(n_16699)
);

OAI21x1_ASAP7_75t_L g16700 ( 
.A1(n_16321),
.A2(n_2237),
.B(n_2238),
.Y(n_16700)
);

BUFx3_ASAP7_75t_L g16701 ( 
.A(n_16351),
.Y(n_16701)
);

INVx2_ASAP7_75t_L g16702 ( 
.A(n_16126),
.Y(n_16702)
);

INVx1_ASAP7_75t_L g16703 ( 
.A(n_16173),
.Y(n_16703)
);

INVx1_ASAP7_75t_L g16704 ( 
.A(n_16180),
.Y(n_16704)
);

BUFx2_ASAP7_75t_L g16705 ( 
.A(n_16139),
.Y(n_16705)
);

INVx1_ASAP7_75t_L g16706 ( 
.A(n_16194),
.Y(n_16706)
);

INVx2_ASAP7_75t_L g16707 ( 
.A(n_16485),
.Y(n_16707)
);

INVx2_ASAP7_75t_L g16708 ( 
.A(n_16141),
.Y(n_16708)
);

INVx2_ASAP7_75t_L g16709 ( 
.A(n_16184),
.Y(n_16709)
);

BUFx6f_ASAP7_75t_L g16710 ( 
.A(n_16368),
.Y(n_16710)
);

INVx3_ASAP7_75t_L g16711 ( 
.A(n_16478),
.Y(n_16711)
);

BUFx6f_ASAP7_75t_L g16712 ( 
.A(n_16333),
.Y(n_16712)
);

INVx3_ASAP7_75t_L g16713 ( 
.A(n_16459),
.Y(n_16713)
);

INVx3_ASAP7_75t_L g16714 ( 
.A(n_16473),
.Y(n_16714)
);

AOI22xp5_ASAP7_75t_SL g16715 ( 
.A1(n_16105),
.A2(n_2240),
.B1(n_2238),
.B2(n_2239),
.Y(n_16715)
);

INVx2_ASAP7_75t_L g16716 ( 
.A(n_16189),
.Y(n_16716)
);

INVx1_ASAP7_75t_L g16717 ( 
.A(n_16198),
.Y(n_16717)
);

INVx2_ASAP7_75t_L g16718 ( 
.A(n_16250),
.Y(n_16718)
);

INVx2_ASAP7_75t_L g16719 ( 
.A(n_16134),
.Y(n_16719)
);

NAND2xp5_ASAP7_75t_L g16720 ( 
.A(n_16454),
.B(n_16492),
.Y(n_16720)
);

INVx1_ASAP7_75t_L g16721 ( 
.A(n_16210),
.Y(n_16721)
);

HB1xp67_ASAP7_75t_L g16722 ( 
.A(n_16425),
.Y(n_16722)
);

INVx2_ASAP7_75t_SL g16723 ( 
.A(n_16376),
.Y(n_16723)
);

INVx1_ASAP7_75t_L g16724 ( 
.A(n_16226),
.Y(n_16724)
);

OAI21x1_ASAP7_75t_L g16725 ( 
.A1(n_16221),
.A2(n_2239),
.B(n_2240),
.Y(n_16725)
);

AND2x2_ASAP7_75t_L g16726 ( 
.A(n_16260),
.B(n_2241),
.Y(n_16726)
);

INVx1_ASAP7_75t_L g16727 ( 
.A(n_16234),
.Y(n_16727)
);

AOI22xp33_ASAP7_75t_SL g16728 ( 
.A1(n_16164),
.A2(n_2243),
.B1(n_2241),
.B2(n_2242),
.Y(n_16728)
);

INVx1_ASAP7_75t_L g16729 ( 
.A(n_16248),
.Y(n_16729)
);

OR2x2_ASAP7_75t_L g16730 ( 
.A(n_16465),
.B(n_2243),
.Y(n_16730)
);

OAI21x1_ASAP7_75t_L g16731 ( 
.A1(n_16179),
.A2(n_2244),
.B(n_2245),
.Y(n_16731)
);

INVx3_ASAP7_75t_L g16732 ( 
.A(n_16479),
.Y(n_16732)
);

INVx2_ASAP7_75t_L g16733 ( 
.A(n_16158),
.Y(n_16733)
);

AOI22xp33_ASAP7_75t_L g16734 ( 
.A1(n_16144),
.A2(n_2248),
.B1(n_2245),
.B2(n_2246),
.Y(n_16734)
);

INVx2_ASAP7_75t_L g16735 ( 
.A(n_16256),
.Y(n_16735)
);

INVx2_ASAP7_75t_L g16736 ( 
.A(n_16259),
.Y(n_16736)
);

BUFx6f_ASAP7_75t_L g16737 ( 
.A(n_16433),
.Y(n_16737)
);

INVx2_ASAP7_75t_L g16738 ( 
.A(n_16326),
.Y(n_16738)
);

AOI22xp33_ASAP7_75t_L g16739 ( 
.A1(n_16113),
.A2(n_2250),
.B1(n_2248),
.B2(n_2249),
.Y(n_16739)
);

AND2x2_ASAP7_75t_L g16740 ( 
.A(n_16264),
.B(n_2249),
.Y(n_16740)
);

INVx3_ASAP7_75t_L g16741 ( 
.A(n_16447),
.Y(n_16741)
);

INVx1_ASAP7_75t_L g16742 ( 
.A(n_16343),
.Y(n_16742)
);

INVx2_ASAP7_75t_L g16743 ( 
.A(n_16360),
.Y(n_16743)
);

OA21x2_ASAP7_75t_L g16744 ( 
.A1(n_16251),
.A2(n_2251),
.B(n_2252),
.Y(n_16744)
);

INVx1_ASAP7_75t_L g16745 ( 
.A(n_16102),
.Y(n_16745)
);

NAND2x1p5_ASAP7_75t_L g16746 ( 
.A(n_16249),
.B(n_2251),
.Y(n_16746)
);

AOI22xp5_ASAP7_75t_L g16747 ( 
.A1(n_16383),
.A2(n_2255),
.B1(n_2253),
.B2(n_2254),
.Y(n_16747)
);

INVx1_ASAP7_75t_L g16748 ( 
.A(n_16415),
.Y(n_16748)
);

AND2x2_ASAP7_75t_L g16749 ( 
.A(n_16513),
.B(n_2253),
.Y(n_16749)
);

OR2x2_ASAP7_75t_L g16750 ( 
.A(n_16218),
.B(n_2254),
.Y(n_16750)
);

NOR2xp33_ASAP7_75t_L g16751 ( 
.A(n_16435),
.B(n_2255),
.Y(n_16751)
);

OR2x2_ASAP7_75t_L g16752 ( 
.A(n_16112),
.B(n_2256),
.Y(n_16752)
);

NAND2xp5_ASAP7_75t_L g16753 ( 
.A(n_16486),
.B(n_2256),
.Y(n_16753)
);

INVx2_ASAP7_75t_SL g16754 ( 
.A(n_16332),
.Y(n_16754)
);

INVx1_ASAP7_75t_L g16755 ( 
.A(n_16227),
.Y(n_16755)
);

INVx2_ASAP7_75t_L g16756 ( 
.A(n_16209),
.Y(n_16756)
);

INVx3_ASAP7_75t_L g16757 ( 
.A(n_16329),
.Y(n_16757)
);

INVx1_ASAP7_75t_L g16758 ( 
.A(n_16494),
.Y(n_16758)
);

INVx4_ASAP7_75t_L g16759 ( 
.A(n_16421),
.Y(n_16759)
);

HB1xp67_ASAP7_75t_L g16760 ( 
.A(n_16171),
.Y(n_16760)
);

INVx1_ASAP7_75t_L g16761 ( 
.A(n_16303),
.Y(n_16761)
);

INVx3_ASAP7_75t_L g16762 ( 
.A(n_16446),
.Y(n_16762)
);

HB1xp67_ASAP7_75t_L g16763 ( 
.A(n_16202),
.Y(n_16763)
);

AND2x4_ASAP7_75t_L g16764 ( 
.A(n_16228),
.B(n_2257),
.Y(n_16764)
);

OAI21xp5_ASAP7_75t_L g16765 ( 
.A1(n_16315),
.A2(n_16185),
.B(n_16236),
.Y(n_16765)
);

BUFx2_ASAP7_75t_L g16766 ( 
.A(n_16424),
.Y(n_16766)
);

INVx1_ASAP7_75t_SL g16767 ( 
.A(n_16509),
.Y(n_16767)
);

INVx1_ASAP7_75t_L g16768 ( 
.A(n_16483),
.Y(n_16768)
);

INVx2_ASAP7_75t_L g16769 ( 
.A(n_16474),
.Y(n_16769)
);

INVx1_ASAP7_75t_L g16770 ( 
.A(n_16488),
.Y(n_16770)
);

INVx1_ASAP7_75t_L g16771 ( 
.A(n_16406),
.Y(n_16771)
);

INVx2_ASAP7_75t_L g16772 ( 
.A(n_16519),
.Y(n_16772)
);

AOI22xp33_ASAP7_75t_L g16773 ( 
.A1(n_16274),
.A2(n_16276),
.B1(n_16386),
.B2(n_16152),
.Y(n_16773)
);

OAI21x1_ASAP7_75t_L g16774 ( 
.A1(n_16089),
.A2(n_2258),
.B(n_2259),
.Y(n_16774)
);

CKINVDCx5p33_ASAP7_75t_R g16775 ( 
.A(n_16467),
.Y(n_16775)
);

INVx2_ASAP7_75t_SL g16776 ( 
.A(n_16393),
.Y(n_16776)
);

BUFx2_ASAP7_75t_SL g16777 ( 
.A(n_16445),
.Y(n_16777)
);

HB1xp67_ASAP7_75t_L g16778 ( 
.A(n_16235),
.Y(n_16778)
);

AND2x2_ASAP7_75t_L g16779 ( 
.A(n_16182),
.B(n_2258),
.Y(n_16779)
);

INVx1_ASAP7_75t_L g16780 ( 
.A(n_16396),
.Y(n_16780)
);

BUFx12f_ASAP7_75t_L g16781 ( 
.A(n_16467),
.Y(n_16781)
);

AO21x2_ASAP7_75t_L g16782 ( 
.A1(n_16119),
.A2(n_2259),
.B(n_2260),
.Y(n_16782)
);

BUFx2_ASAP7_75t_L g16783 ( 
.A(n_16276),
.Y(n_16783)
);

HB1xp67_ASAP7_75t_L g16784 ( 
.A(n_16515),
.Y(n_16784)
);

INVx1_ASAP7_75t_L g16785 ( 
.A(n_16397),
.Y(n_16785)
);

OA21x2_ASAP7_75t_L g16786 ( 
.A1(n_16244),
.A2(n_2260),
.B(n_2261),
.Y(n_16786)
);

INVx1_ASAP7_75t_L g16787 ( 
.A(n_16192),
.Y(n_16787)
);

AND2x2_ASAP7_75t_L g16788 ( 
.A(n_16167),
.B(n_2261),
.Y(n_16788)
);

INVx3_ASAP7_75t_SL g16789 ( 
.A(n_16390),
.Y(n_16789)
);

INVx1_ASAP7_75t_L g16790 ( 
.A(n_16205),
.Y(n_16790)
);

INVx1_ASAP7_75t_L g16791 ( 
.A(n_16327),
.Y(n_16791)
);

INVx1_ASAP7_75t_L g16792 ( 
.A(n_16312),
.Y(n_16792)
);

OR2x2_ASAP7_75t_L g16793 ( 
.A(n_16242),
.B(n_16293),
.Y(n_16793)
);

NAND2x1p5_ASAP7_75t_L g16794 ( 
.A(n_16240),
.B(n_16313),
.Y(n_16794)
);

INVx2_ASAP7_75t_L g16795 ( 
.A(n_16457),
.Y(n_16795)
);

NAND2xp5_ASAP7_75t_L g16796 ( 
.A(n_16431),
.B(n_2262),
.Y(n_16796)
);

INVx3_ASAP7_75t_L g16797 ( 
.A(n_16172),
.Y(n_16797)
);

INVx1_ASAP7_75t_L g16798 ( 
.A(n_16347),
.Y(n_16798)
);

HB1xp67_ASAP7_75t_L g16799 ( 
.A(n_16461),
.Y(n_16799)
);

INVx1_ASAP7_75t_L g16800 ( 
.A(n_16361),
.Y(n_16800)
);

HB1xp67_ASAP7_75t_L g16801 ( 
.A(n_16093),
.Y(n_16801)
);

NOR2xp33_ASAP7_75t_L g16802 ( 
.A(n_16193),
.B(n_2262),
.Y(n_16802)
);

INVx2_ASAP7_75t_L g16803 ( 
.A(n_16245),
.Y(n_16803)
);

INVx2_ASAP7_75t_SL g16804 ( 
.A(n_16439),
.Y(n_16804)
);

CKINVDCx20_ASAP7_75t_R g16805 ( 
.A(n_16416),
.Y(n_16805)
);

OR2x2_ASAP7_75t_L g16806 ( 
.A(n_16157),
.B(n_2263),
.Y(n_16806)
);

HB1xp67_ASAP7_75t_L g16807 ( 
.A(n_16213),
.Y(n_16807)
);

INVx2_ASAP7_75t_L g16808 ( 
.A(n_16231),
.Y(n_16808)
);

INVx2_ASAP7_75t_L g16809 ( 
.A(n_16381),
.Y(n_16809)
);

INVx1_ASAP7_75t_L g16810 ( 
.A(n_16365),
.Y(n_16810)
);

AND2x2_ASAP7_75t_L g16811 ( 
.A(n_16224),
.B(n_2263),
.Y(n_16811)
);

AND2x2_ASAP7_75t_L g16812 ( 
.A(n_16094),
.B(n_16196),
.Y(n_16812)
);

INVx1_ASAP7_75t_L g16813 ( 
.A(n_16379),
.Y(n_16813)
);

OAI21xp5_ASAP7_75t_L g16814 ( 
.A1(n_16097),
.A2(n_2264),
.B(n_2265),
.Y(n_16814)
);

OR2x2_ASAP7_75t_L g16815 ( 
.A(n_16307),
.B(n_2264),
.Y(n_16815)
);

INVx2_ASAP7_75t_SL g16816 ( 
.A(n_16451),
.Y(n_16816)
);

HB1xp67_ASAP7_75t_L g16817 ( 
.A(n_16121),
.Y(n_16817)
);

AND2x4_ASAP7_75t_L g16818 ( 
.A(n_16342),
.B(n_2265),
.Y(n_16818)
);

INVx1_ASAP7_75t_L g16819 ( 
.A(n_16380),
.Y(n_16819)
);

INVx1_ASAP7_75t_L g16820 ( 
.A(n_16385),
.Y(n_16820)
);

INVx1_ASAP7_75t_L g16821 ( 
.A(n_16389),
.Y(n_16821)
);

INVxp33_ASAP7_75t_L g16822 ( 
.A(n_16219),
.Y(n_16822)
);

AOI21x1_ASAP7_75t_L g16823 ( 
.A1(n_16296),
.A2(n_2266),
.B(n_2267),
.Y(n_16823)
);

BUFx3_ASAP7_75t_L g16824 ( 
.A(n_16427),
.Y(n_16824)
);

INVx1_ASAP7_75t_L g16825 ( 
.A(n_16470),
.Y(n_16825)
);

INVx2_ASAP7_75t_L g16826 ( 
.A(n_16247),
.Y(n_16826)
);

INVx1_ASAP7_75t_L g16827 ( 
.A(n_16469),
.Y(n_16827)
);

INVx1_ASAP7_75t_L g16828 ( 
.A(n_16310),
.Y(n_16828)
);

INVx1_ASAP7_75t_L g16829 ( 
.A(n_16344),
.Y(n_16829)
);

INVx1_ASAP7_75t_L g16830 ( 
.A(n_16348),
.Y(n_16830)
);

INVx2_ASAP7_75t_L g16831 ( 
.A(n_16384),
.Y(n_16831)
);

AOI21x1_ASAP7_75t_L g16832 ( 
.A1(n_16341),
.A2(n_2267),
.B(n_2268),
.Y(n_16832)
);

INVx3_ASAP7_75t_L g16833 ( 
.A(n_16456),
.Y(n_16833)
);

BUFx2_ASAP7_75t_L g16834 ( 
.A(n_16490),
.Y(n_16834)
);

INVx2_ASAP7_75t_L g16835 ( 
.A(n_16507),
.Y(n_16835)
);

INVx1_ASAP7_75t_L g16836 ( 
.A(n_16369),
.Y(n_16836)
);

OAI21x1_ASAP7_75t_L g16837 ( 
.A1(n_16149),
.A2(n_2268),
.B(n_2269),
.Y(n_16837)
);

INVx1_ASAP7_75t_L g16838 ( 
.A(n_16334),
.Y(n_16838)
);

AND2x2_ASAP7_75t_L g16839 ( 
.A(n_16294),
.B(n_16335),
.Y(n_16839)
);

INVx1_ASAP7_75t_L g16840 ( 
.A(n_16450),
.Y(n_16840)
);

INVx1_ASAP7_75t_L g16841 ( 
.A(n_16462),
.Y(n_16841)
);

INVx2_ASAP7_75t_SL g16842 ( 
.A(n_16300),
.Y(n_16842)
);

AND2x2_ASAP7_75t_L g16843 ( 
.A(n_16378),
.B(n_2269),
.Y(n_16843)
);

INVx3_ASAP7_75t_L g16844 ( 
.A(n_16305),
.Y(n_16844)
);

INVx2_ASAP7_75t_L g16845 ( 
.A(n_16246),
.Y(n_16845)
);

INVx2_ASAP7_75t_L g16846 ( 
.A(n_16436),
.Y(n_16846)
);

OR2x2_ASAP7_75t_L g16847 ( 
.A(n_16263),
.B(n_2270),
.Y(n_16847)
);

INVx1_ASAP7_75t_L g16848 ( 
.A(n_16400),
.Y(n_16848)
);

AO21x1_ASAP7_75t_SL g16849 ( 
.A1(n_16501),
.A2(n_2270),
.B(n_2271),
.Y(n_16849)
);

INVx1_ASAP7_75t_L g16850 ( 
.A(n_16499),
.Y(n_16850)
);

AO31x2_ASAP7_75t_L g16851 ( 
.A1(n_16440),
.A2(n_2273),
.A3(n_2271),
.B(n_2272),
.Y(n_16851)
);

AOI22xp33_ASAP7_75t_L g16852 ( 
.A1(n_16258),
.A2(n_2274),
.B1(n_2272),
.B2(n_2273),
.Y(n_16852)
);

AOI22xp5_ASAP7_75t_L g16853 ( 
.A1(n_16207),
.A2(n_2276),
.B1(n_2274),
.B2(n_2275),
.Y(n_16853)
);

INVx1_ASAP7_75t_L g16854 ( 
.A(n_16292),
.Y(n_16854)
);

INVx1_ASAP7_75t_L g16855 ( 
.A(n_16325),
.Y(n_16855)
);

INVx2_ASAP7_75t_L g16856 ( 
.A(n_16505),
.Y(n_16856)
);

INVx2_ASAP7_75t_SL g16857 ( 
.A(n_16506),
.Y(n_16857)
);

INVx1_ASAP7_75t_L g16858 ( 
.A(n_16458),
.Y(n_16858)
);

INVx1_ASAP7_75t_L g16859 ( 
.A(n_16308),
.Y(n_16859)
);

INVx2_ASAP7_75t_L g16860 ( 
.A(n_16282),
.Y(n_16860)
);

INVx1_ASAP7_75t_L g16861 ( 
.A(n_16267),
.Y(n_16861)
);

INVx3_ASAP7_75t_L g16862 ( 
.A(n_16463),
.Y(n_16862)
);

OAI22xp5_ASAP7_75t_L g16863 ( 
.A1(n_16120),
.A2(n_2278),
.B1(n_2275),
.B2(n_2277),
.Y(n_16863)
);

INVx1_ASAP7_75t_L g16864 ( 
.A(n_16270),
.Y(n_16864)
);

AND2x4_ASAP7_75t_L g16865 ( 
.A(n_16398),
.B(n_2277),
.Y(n_16865)
);

INVx4_ASAP7_75t_L g16866 ( 
.A(n_16489),
.Y(n_16866)
);

AND2x2_ASAP7_75t_L g16867 ( 
.A(n_16257),
.B(n_2278),
.Y(n_16867)
);

BUFx6f_ASAP7_75t_L g16868 ( 
.A(n_16502),
.Y(n_16868)
);

INVx2_ASAP7_75t_L g16869 ( 
.A(n_16503),
.Y(n_16869)
);

INVx2_ASAP7_75t_L g16870 ( 
.A(n_16476),
.Y(n_16870)
);

NOR2xp33_ASAP7_75t_L g16871 ( 
.A(n_16496),
.B(n_2279),
.Y(n_16871)
);

INVx1_ASAP7_75t_L g16872 ( 
.A(n_16442),
.Y(n_16872)
);

OAI22xp33_ASAP7_75t_L g16873 ( 
.A1(n_16287),
.A2(n_2281),
.B1(n_2279),
.B2(n_2280),
.Y(n_16873)
);

AND2x4_ASAP7_75t_L g16874 ( 
.A(n_16408),
.B(n_2280),
.Y(n_16874)
);

HB1xp67_ASAP7_75t_L g16875 ( 
.A(n_16265),
.Y(n_16875)
);

INVx2_ASAP7_75t_L g16876 ( 
.A(n_16510),
.Y(n_16876)
);

INVx2_ASAP7_75t_L g16877 ( 
.A(n_16484),
.Y(n_16877)
);

INVx1_ASAP7_75t_L g16878 ( 
.A(n_16443),
.Y(n_16878)
);

INVx2_ASAP7_75t_L g16879 ( 
.A(n_16477),
.Y(n_16879)
);

INVx2_ASAP7_75t_L g16880 ( 
.A(n_16426),
.Y(n_16880)
);

INVx2_ASAP7_75t_L g16881 ( 
.A(n_16269),
.Y(n_16881)
);

OR2x2_ASAP7_75t_L g16882 ( 
.A(n_16418),
.B(n_2281),
.Y(n_16882)
);

INVx1_ASAP7_75t_SL g16883 ( 
.A(n_16116),
.Y(n_16883)
);

BUFx2_ASAP7_75t_L g16884 ( 
.A(n_16444),
.Y(n_16884)
);

NAND3xp33_ASAP7_75t_L g16885 ( 
.A(n_16098),
.B(n_2282),
.C(n_2283),
.Y(n_16885)
);

INVx2_ASAP7_75t_L g16886 ( 
.A(n_16280),
.Y(n_16886)
);

NAND2xp5_ASAP7_75t_L g16887 ( 
.A(n_16500),
.B(n_2283),
.Y(n_16887)
);

AO31x2_ASAP7_75t_L g16888 ( 
.A1(n_16377),
.A2(n_2286),
.A3(n_2284),
.B(n_2285),
.Y(n_16888)
);

AOI22xp5_ASAP7_75t_L g16889 ( 
.A1(n_16177),
.A2(n_2286),
.B1(n_2284),
.B2(n_2285),
.Y(n_16889)
);

CKINVDCx20_ASAP7_75t_R g16890 ( 
.A(n_16409),
.Y(n_16890)
);

INVx1_ASAP7_75t_L g16891 ( 
.A(n_16429),
.Y(n_16891)
);

INVx2_ASAP7_75t_L g16892 ( 
.A(n_16324),
.Y(n_16892)
);

OA21x2_ASAP7_75t_L g16893 ( 
.A1(n_16142),
.A2(n_2287),
.B(n_2288),
.Y(n_16893)
);

AND2x4_ASAP7_75t_L g16894 ( 
.A(n_16363),
.B(n_2288),
.Y(n_16894)
);

OAI21xp5_ASAP7_75t_L g16895 ( 
.A1(n_16354),
.A2(n_16135),
.B(n_16353),
.Y(n_16895)
);

BUFx2_ASAP7_75t_L g16896 ( 
.A(n_16163),
.Y(n_16896)
);

OAI21x1_ASAP7_75t_L g16897 ( 
.A1(n_16115),
.A2(n_16147),
.B(n_16464),
.Y(n_16897)
);

INVx3_ASAP7_75t_L g16898 ( 
.A(n_16508),
.Y(n_16898)
);

BUFx2_ASAP7_75t_L g16899 ( 
.A(n_16159),
.Y(n_16899)
);

HB1xp67_ASAP7_75t_L g16900 ( 
.A(n_16562),
.Y(n_16900)
);

BUFx3_ASAP7_75t_L g16901 ( 
.A(n_16550),
.Y(n_16901)
);

OAI21x1_ASAP7_75t_L g16902 ( 
.A1(n_16600),
.A2(n_16130),
.B(n_16410),
.Y(n_16902)
);

CKINVDCx12_ASAP7_75t_R g16903 ( 
.A(n_16715),
.Y(n_16903)
);

AND2x2_ASAP7_75t_L g16904 ( 
.A(n_16522),
.B(n_16495),
.Y(n_16904)
);

CKINVDCx16_ASAP7_75t_R g16905 ( 
.A(n_16781),
.Y(n_16905)
);

OR2x6_ASAP7_75t_L g16906 ( 
.A(n_16777),
.B(n_16411),
.Y(n_16906)
);

AND2x2_ASAP7_75t_L g16907 ( 
.A(n_16640),
.B(n_16530),
.Y(n_16907)
);

OR2x6_ASAP7_75t_L g16908 ( 
.A(n_16687),
.B(n_16306),
.Y(n_16908)
);

NOR3xp33_ASAP7_75t_SL g16909 ( 
.A(n_16765),
.B(n_16405),
.C(n_16399),
.Y(n_16909)
);

CKINVDCx5p33_ASAP7_75t_R g16910 ( 
.A(n_16537),
.Y(n_16910)
);

INVx4_ASAP7_75t_SL g16911 ( 
.A(n_16528),
.Y(n_16911)
);

NAND2xp5_ASAP7_75t_L g16912 ( 
.A(n_16853),
.B(n_16359),
.Y(n_16912)
);

INVx2_ASAP7_75t_L g16913 ( 
.A(n_16529),
.Y(n_16913)
);

INVx2_ASAP7_75t_L g16914 ( 
.A(n_16668),
.Y(n_16914)
);

AND2x2_ASAP7_75t_L g16915 ( 
.A(n_16559),
.B(n_16468),
.Y(n_16915)
);

INVx2_ASAP7_75t_L g16916 ( 
.A(n_16572),
.Y(n_16916)
);

AOI22xp33_ASAP7_75t_L g16917 ( 
.A1(n_16896),
.A2(n_16168),
.B1(n_16155),
.B2(n_16206),
.Y(n_16917)
);

OA21x2_ASAP7_75t_L g16918 ( 
.A1(n_16773),
.A2(n_16350),
.B(n_16319),
.Y(n_16918)
);

INVx4_ASAP7_75t_L g16919 ( 
.A(n_16572),
.Y(n_16919)
);

HB1xp67_ASAP7_75t_L g16920 ( 
.A(n_16527),
.Y(n_16920)
);

INVx2_ASAP7_75t_L g16921 ( 
.A(n_16616),
.Y(n_16921)
);

OAI22xp5_ASAP7_75t_L g16922 ( 
.A1(n_16692),
.A2(n_16212),
.B1(n_16302),
.B2(n_16317),
.Y(n_16922)
);

AOI22xp33_ASAP7_75t_L g16923 ( 
.A1(n_16698),
.A2(n_16284),
.B1(n_16497),
.B2(n_16472),
.Y(n_16923)
);

CKINVDCx5p33_ASAP7_75t_R g16924 ( 
.A(n_16667),
.Y(n_16924)
);

INVx2_ASAP7_75t_L g16925 ( 
.A(n_16616),
.Y(n_16925)
);

NAND3xp33_ASAP7_75t_SL g16926 ( 
.A(n_16884),
.B(n_16124),
.C(n_16518),
.Y(n_16926)
);

OR2x6_ASAP7_75t_L g16927 ( 
.A(n_16535),
.B(n_16367),
.Y(n_16927)
);

AND2x2_ASAP7_75t_L g16928 ( 
.A(n_16552),
.B(n_16281),
.Y(n_16928)
);

NOR3xp33_ASAP7_75t_SL g16929 ( 
.A(n_16556),
.B(n_16504),
.C(n_16299),
.Y(n_16929)
);

INVx1_ASAP7_75t_L g16930 ( 
.A(n_16763),
.Y(n_16930)
);

BUFx4f_ASAP7_75t_SL g16931 ( 
.A(n_16678),
.Y(n_16931)
);

AND2x2_ASAP7_75t_L g16932 ( 
.A(n_16684),
.B(n_16339),
.Y(n_16932)
);

AO31x2_ASAP7_75t_L g16933 ( 
.A1(n_16705),
.A2(n_16471),
.A3(n_16338),
.B(n_16352),
.Y(n_16933)
);

INVx1_ASAP7_75t_L g16934 ( 
.A(n_16549),
.Y(n_16934)
);

OAI22xp33_ASAP7_75t_SL g16935 ( 
.A1(n_16617),
.A2(n_16419),
.B1(n_16395),
.B2(n_16512),
.Y(n_16935)
);

NAND2xp5_ASAP7_75t_L g16936 ( 
.A(n_16677),
.B(n_16291),
.Y(n_16936)
);

BUFx8_ASAP7_75t_SL g16937 ( 
.A(n_16597),
.Y(n_16937)
);

AND2x4_ASAP7_75t_L g16938 ( 
.A(n_16650),
.B(n_16526),
.Y(n_16938)
);

INVx3_ASAP7_75t_L g16939 ( 
.A(n_16563),
.Y(n_16939)
);

BUFx3_ASAP7_75t_L g16940 ( 
.A(n_16663),
.Y(n_16940)
);

BUFx6f_ASAP7_75t_L g16941 ( 
.A(n_16660),
.Y(n_16941)
);

NOR2xp33_ASAP7_75t_R g16942 ( 
.A(n_16775),
.B(n_2289),
.Y(n_16942)
);

INVx1_ASAP7_75t_L g16943 ( 
.A(n_16579),
.Y(n_16943)
);

AOI22xp33_ASAP7_75t_L g16944 ( 
.A1(n_16899),
.A2(n_16517),
.B1(n_16491),
.B2(n_16481),
.Y(n_16944)
);

INVx3_ASAP7_75t_L g16945 ( 
.A(n_16710),
.Y(n_16945)
);

NOR2xp33_ASAP7_75t_R g16946 ( 
.A(n_16586),
.B(n_16632),
.Y(n_16946)
);

NOR2xp33_ASAP7_75t_R g16947 ( 
.A(n_16797),
.B(n_2289),
.Y(n_16947)
);

INVx1_ASAP7_75t_L g16948 ( 
.A(n_16758),
.Y(n_16948)
);

INVx3_ASAP7_75t_L g16949 ( 
.A(n_16710),
.Y(n_16949)
);

INVx2_ASAP7_75t_L g16950 ( 
.A(n_16592),
.Y(n_16950)
);

INVxp67_ASAP7_75t_SL g16951 ( 
.A(n_16746),
.Y(n_16951)
);

AND2x2_ASAP7_75t_L g16952 ( 
.A(n_16596),
.B(n_16268),
.Y(n_16952)
);

NAND2xp33_ASAP7_75t_SL g16953 ( 
.A(n_16805),
.B(n_16516),
.Y(n_16953)
);

OR2x2_ASAP7_75t_L g16954 ( 
.A(n_16582),
.B(n_16394),
.Y(n_16954)
);

AO31x2_ASAP7_75t_L g16955 ( 
.A1(n_16783),
.A2(n_16520),
.A3(n_16441),
.B(n_16423),
.Y(n_16955)
);

AOI21xp5_ASAP7_75t_L g16956 ( 
.A1(n_16895),
.A2(n_16225),
.B(n_16375),
.Y(n_16956)
);

AND2x2_ASAP7_75t_L g16957 ( 
.A(n_16672),
.B(n_2290),
.Y(n_16957)
);

NAND2xp5_ASAP7_75t_L g16958 ( 
.A(n_16834),
.B(n_16691),
.Y(n_16958)
);

NAND2xp33_ASAP7_75t_SL g16959 ( 
.A(n_16609),
.B(n_16482),
.Y(n_16959)
);

BUFx2_ASAP7_75t_L g16960 ( 
.A(n_16551),
.Y(n_16960)
);

OA21x2_ASAP7_75t_L g16961 ( 
.A1(n_16565),
.A2(n_2290),
.B(n_2291),
.Y(n_16961)
);

INVx2_ASAP7_75t_SL g16962 ( 
.A(n_16712),
.Y(n_16962)
);

NAND2xp33_ASAP7_75t_R g16963 ( 
.A(n_16893),
.B(n_2291),
.Y(n_16963)
);

AND2x4_ASAP7_75t_SL g16964 ( 
.A(n_16759),
.B(n_16712),
.Y(n_16964)
);

CKINVDCx20_ASAP7_75t_R g16965 ( 
.A(n_16890),
.Y(n_16965)
);

AND2x2_ASAP7_75t_L g16966 ( 
.A(n_16713),
.B(n_2292),
.Y(n_16966)
);

AND2x4_ASAP7_75t_L g16967 ( 
.A(n_16649),
.B(n_2293),
.Y(n_16967)
);

INVx3_ASAP7_75t_L g16968 ( 
.A(n_16701),
.Y(n_16968)
);

BUFx2_ASAP7_75t_L g16969 ( 
.A(n_16794),
.Y(n_16969)
);

INVx1_ASAP7_75t_L g16970 ( 
.A(n_16768),
.Y(n_16970)
);

INVx1_ASAP7_75t_L g16971 ( 
.A(n_16770),
.Y(n_16971)
);

NOR2xp33_ASAP7_75t_R g16972 ( 
.A(n_16898),
.B(n_2293),
.Y(n_16972)
);

NAND2xp33_ASAP7_75t_R g16973 ( 
.A(n_16786),
.B(n_2294),
.Y(n_16973)
);

INVx2_ASAP7_75t_L g16974 ( 
.A(n_16543),
.Y(n_16974)
);

OR2x6_ASAP7_75t_L g16975 ( 
.A(n_16814),
.B(n_2294),
.Y(n_16975)
);

INVx2_ASAP7_75t_L g16976 ( 
.A(n_16737),
.Y(n_16976)
);

BUFx6f_ASAP7_75t_L g16977 ( 
.A(n_16676),
.Y(n_16977)
);

NOR2xp33_ASAP7_75t_R g16978 ( 
.A(n_16757),
.B(n_2295),
.Y(n_16978)
);

AOI22xp33_ASAP7_75t_L g16979 ( 
.A1(n_16865),
.A2(n_2297),
.B1(n_2295),
.B2(n_2296),
.Y(n_16979)
);

INVxp67_ASAP7_75t_L g16980 ( 
.A(n_16689),
.Y(n_16980)
);

CKINVDCx5p33_ASAP7_75t_R g16981 ( 
.A(n_16589),
.Y(n_16981)
);

INVx1_ASAP7_75t_L g16982 ( 
.A(n_16540),
.Y(n_16982)
);

INVx2_ASAP7_75t_L g16983 ( 
.A(n_16737),
.Y(n_16983)
);

NOR2xp33_ASAP7_75t_R g16984 ( 
.A(n_16762),
.B(n_2297),
.Y(n_16984)
);

INVx1_ASAP7_75t_L g16985 ( 
.A(n_16545),
.Y(n_16985)
);

AND2x2_ASAP7_75t_L g16986 ( 
.A(n_16711),
.B(n_2298),
.Y(n_16986)
);

INVx1_ASAP7_75t_L g16987 ( 
.A(n_16548),
.Y(n_16987)
);

CKINVDCx12_ASAP7_75t_R g16988 ( 
.A(n_16630),
.Y(n_16988)
);

BUFx2_ASAP7_75t_L g16989 ( 
.A(n_16824),
.Y(n_16989)
);

HB1xp67_ASAP7_75t_L g16990 ( 
.A(n_16741),
.Y(n_16990)
);

AO31x2_ASAP7_75t_L g16991 ( 
.A1(n_16587),
.A2(n_2300),
.A3(n_2298),
.B(n_2299),
.Y(n_16991)
);

INVx2_ASAP7_75t_L g16992 ( 
.A(n_16868),
.Y(n_16992)
);

AND2x2_ASAP7_75t_L g16993 ( 
.A(n_16567),
.B(n_2300),
.Y(n_16993)
);

NOR2xp33_ASAP7_75t_R g16994 ( 
.A(n_16658),
.B(n_16564),
.Y(n_16994)
);

NAND2xp33_ASAP7_75t_R g16995 ( 
.A(n_16744),
.B(n_2301),
.Y(n_16995)
);

INVx4_ASAP7_75t_L g16996 ( 
.A(n_16589),
.Y(n_16996)
);

AND2x6_ASAP7_75t_L g16997 ( 
.A(n_16764),
.B(n_2301),
.Y(n_16997)
);

CKINVDCx16_ASAP7_75t_R g16998 ( 
.A(n_16874),
.Y(n_16998)
);

OAI21x1_ASAP7_75t_L g16999 ( 
.A1(n_16555),
.A2(n_2302),
.B(n_2303),
.Y(n_16999)
);

AND2x4_ASAP7_75t_SL g17000 ( 
.A(n_16546),
.B(n_2302),
.Y(n_17000)
);

CKINVDCx8_ASAP7_75t_R g17001 ( 
.A(n_16818),
.Y(n_17001)
);

OR2x2_ASAP7_75t_L g17002 ( 
.A(n_16606),
.B(n_16825),
.Y(n_17002)
);

AND2x2_ASAP7_75t_L g17003 ( 
.A(n_16580),
.B(n_16574),
.Y(n_17003)
);

OAI21xp5_ASAP7_75t_L g17004 ( 
.A1(n_16897),
.A2(n_2303),
.B(n_2304),
.Y(n_17004)
);

NAND2xp33_ASAP7_75t_R g17005 ( 
.A(n_16697),
.B(n_2304),
.Y(n_17005)
);

NAND2xp5_ASAP7_75t_L g17006 ( 
.A(n_16892),
.B(n_2305),
.Y(n_17006)
);

CKINVDCx8_ASAP7_75t_R g17007 ( 
.A(n_16686),
.Y(n_17007)
);

OR2x6_ASAP7_75t_L g17008 ( 
.A(n_16885),
.B(n_2305),
.Y(n_17008)
);

INVx1_ASAP7_75t_L g17009 ( 
.A(n_16553),
.Y(n_17009)
);

AO31x2_ASAP7_75t_L g17010 ( 
.A1(n_16599),
.A2(n_2309),
.A3(n_2307),
.B(n_2308),
.Y(n_17010)
);

CKINVDCx5p33_ASAP7_75t_R g17011 ( 
.A(n_16883),
.Y(n_17011)
);

INVx4_ASAP7_75t_L g17012 ( 
.A(n_16695),
.Y(n_17012)
);

NOR2xp33_ASAP7_75t_L g17013 ( 
.A(n_16822),
.B(n_2307),
.Y(n_17013)
);

INVx2_ASAP7_75t_L g17014 ( 
.A(n_16868),
.Y(n_17014)
);

NOR2xp33_ASAP7_75t_R g17015 ( 
.A(n_16823),
.B(n_2308),
.Y(n_17015)
);

INVx1_ASAP7_75t_L g17016 ( 
.A(n_16557),
.Y(n_17016)
);

NAND2x1p5_ASAP7_75t_L g17017 ( 
.A(n_16619),
.B(n_2309),
.Y(n_17017)
);

NOR3xp33_ASAP7_75t_SL g17018 ( 
.A(n_16615),
.B(n_2310),
.C(n_2311),
.Y(n_17018)
);

NAND2xp5_ASAP7_75t_L g17019 ( 
.A(n_16855),
.B(n_2311),
.Y(n_17019)
);

NAND2xp5_ASAP7_75t_L g17020 ( 
.A(n_16674),
.B(n_16857),
.Y(n_17020)
);

AND2x2_ASAP7_75t_L g17021 ( 
.A(n_16603),
.B(n_2312),
.Y(n_17021)
);

NOR2xp67_ASAP7_75t_L g17022 ( 
.A(n_16722),
.B(n_16866),
.Y(n_17022)
);

HB1xp67_ASAP7_75t_L g17023 ( 
.A(n_16760),
.Y(n_17023)
);

AND2x4_ASAP7_75t_L g17024 ( 
.A(n_16584),
.B(n_2312),
.Y(n_17024)
);

AOI22xp33_ASAP7_75t_L g17025 ( 
.A1(n_16646),
.A2(n_2315),
.B1(n_2313),
.B2(n_2314),
.Y(n_17025)
);

AO31x2_ASAP7_75t_L g17026 ( 
.A1(n_16593),
.A2(n_2315),
.A3(n_2313),
.B(n_2314),
.Y(n_17026)
);

INVxp33_ASAP7_75t_SL g17027 ( 
.A(n_16751),
.Y(n_17027)
);

AND2x2_ASAP7_75t_L g17028 ( 
.A(n_16651),
.B(n_2316),
.Y(n_17028)
);

INVx2_ASAP7_75t_L g17029 ( 
.A(n_16833),
.Y(n_17029)
);

AND2x4_ASAP7_75t_L g17030 ( 
.A(n_16591),
.B(n_2316),
.Y(n_17030)
);

INVx1_ASAP7_75t_L g17031 ( 
.A(n_16560),
.Y(n_17031)
);

HB1xp67_ASAP7_75t_L g17032 ( 
.A(n_16602),
.Y(n_17032)
);

AND2x2_ASAP7_75t_L g17033 ( 
.A(n_16525),
.B(n_2317),
.Y(n_17033)
);

NAND2xp33_ASAP7_75t_R g17034 ( 
.A(n_16531),
.B(n_2317),
.Y(n_17034)
);

OR2x6_ASAP7_75t_L g17035 ( 
.A(n_16804),
.B(n_2318),
.Y(n_17035)
);

AND2x2_ASAP7_75t_L g17036 ( 
.A(n_16839),
.B(n_2318),
.Y(n_17036)
);

AND2x4_ASAP7_75t_L g17037 ( 
.A(n_16554),
.B(n_2320),
.Y(n_17037)
);

NAND2xp33_ASAP7_75t_R g17038 ( 
.A(n_16788),
.B(n_2320),
.Y(n_17038)
);

NOR3xp33_ASAP7_75t_SL g17039 ( 
.A(n_16873),
.B(n_2321),
.C(n_2322),
.Y(n_17039)
);

INVxp67_ASAP7_75t_L g17040 ( 
.A(n_16849),
.Y(n_17040)
);

INVx3_ASAP7_75t_L g17041 ( 
.A(n_16862),
.Y(n_17041)
);

OR2x2_ASAP7_75t_L g17042 ( 
.A(n_16793),
.B(n_2321),
.Y(n_17042)
);

NAND3xp33_ASAP7_75t_L g17043 ( 
.A(n_16643),
.B(n_2322),
.C(n_2323),
.Y(n_17043)
);

AND2x2_ASAP7_75t_L g17044 ( 
.A(n_16809),
.B(n_2323),
.Y(n_17044)
);

INVx3_ASAP7_75t_L g17045 ( 
.A(n_16547),
.Y(n_17045)
);

AND2x2_ASAP7_75t_L g17046 ( 
.A(n_16879),
.B(n_2324),
.Y(n_17046)
);

NOR2xp33_ASAP7_75t_R g17047 ( 
.A(n_16832),
.B(n_2325),
.Y(n_17047)
);

O2A1O1Ixp5_ASAP7_75t_SL g17048 ( 
.A1(n_16748),
.A2(n_2327),
.B(n_2325),
.C(n_2326),
.Y(n_17048)
);

NAND2xp5_ASAP7_75t_L g17049 ( 
.A(n_16644),
.B(n_2326),
.Y(n_17049)
);

AND2x2_ASAP7_75t_L g17050 ( 
.A(n_16776),
.B(n_2327),
.Y(n_17050)
);

OAI21xp5_ASAP7_75t_L g17051 ( 
.A1(n_16610),
.A2(n_2329),
.B(n_2330),
.Y(n_17051)
);

NAND2xp33_ASAP7_75t_R g17052 ( 
.A(n_16894),
.B(n_2329),
.Y(n_17052)
);

INVx1_ASAP7_75t_L g17053 ( 
.A(n_16561),
.Y(n_17053)
);

CKINVDCx16_ASAP7_75t_R g17054 ( 
.A(n_16754),
.Y(n_17054)
);

AND2x2_ASAP7_75t_L g17055 ( 
.A(n_16835),
.B(n_16877),
.Y(n_17055)
);

AOI22xp33_ASAP7_75t_L g17056 ( 
.A1(n_16581),
.A2(n_2332),
.B1(n_2330),
.B2(n_2331),
.Y(n_17056)
);

INVx1_ASAP7_75t_L g17057 ( 
.A(n_16566),
.Y(n_17057)
);

A2O1A1Ixp33_ASAP7_75t_L g17058 ( 
.A1(n_16889),
.A2(n_2333),
.B(n_2331),
.C(n_2332),
.Y(n_17058)
);

INVx1_ASAP7_75t_L g17059 ( 
.A(n_16846),
.Y(n_17059)
);

INVx2_ASAP7_75t_SL g17060 ( 
.A(n_16789),
.Y(n_17060)
);

NAND2xp33_ASAP7_75t_R g17061 ( 
.A(n_16779),
.B(n_2333),
.Y(n_17061)
);

INVx2_ASAP7_75t_L g17062 ( 
.A(n_16844),
.Y(n_17062)
);

NAND2xp33_ASAP7_75t_R g17063 ( 
.A(n_16749),
.B(n_2334),
.Y(n_17063)
);

NAND2x1_ASAP7_75t_L g17064 ( 
.A(n_16826),
.B(n_2334),
.Y(n_17064)
);

INVx3_ASAP7_75t_L g17065 ( 
.A(n_16714),
.Y(n_17065)
);

BUFx3_ASAP7_75t_L g17066 ( 
.A(n_16611),
.Y(n_17066)
);

AND2x2_ASAP7_75t_L g17067 ( 
.A(n_16541),
.B(n_16718),
.Y(n_17067)
);

BUFx3_ASAP7_75t_L g17068 ( 
.A(n_16614),
.Y(n_17068)
);

INVx2_ASAP7_75t_L g17069 ( 
.A(n_16669),
.Y(n_17069)
);

AOI22xp33_ASAP7_75t_SL g17070 ( 
.A1(n_16827),
.A2(n_2337),
.B1(n_2335),
.B2(n_2336),
.Y(n_17070)
);

OR2x6_ASAP7_75t_L g17071 ( 
.A(n_16816),
.B(n_2335),
.Y(n_17071)
);

CKINVDCx16_ASAP7_75t_R g17072 ( 
.A(n_16863),
.Y(n_17072)
);

OR2x6_ASAP7_75t_L g17073 ( 
.A(n_16869),
.B(n_2336),
.Y(n_17073)
);

INVx2_ASAP7_75t_L g17074 ( 
.A(n_16679),
.Y(n_17074)
);

NAND2xp33_ASAP7_75t_R g17075 ( 
.A(n_16811),
.B(n_2338),
.Y(n_17075)
);

INVx1_ASAP7_75t_L g17076 ( 
.A(n_16571),
.Y(n_17076)
);

INVx3_ASAP7_75t_L g17077 ( 
.A(n_16732),
.Y(n_17077)
);

INVx1_ASAP7_75t_L g17078 ( 
.A(n_16761),
.Y(n_17078)
);

INVx2_ASAP7_75t_L g17079 ( 
.A(n_16682),
.Y(n_17079)
);

AOI22xp33_ASAP7_75t_SL g17080 ( 
.A1(n_16886),
.A2(n_2340),
.B1(n_2338),
.B2(n_2339),
.Y(n_17080)
);

AND2x2_ASAP7_75t_L g17081 ( 
.A(n_16880),
.B(n_2340),
.Y(n_17081)
);

INVx1_ASAP7_75t_L g17082 ( 
.A(n_16771),
.Y(n_17082)
);

NOR2xp33_ASAP7_75t_R g17083 ( 
.A(n_16648),
.B(n_2341),
.Y(n_17083)
);

INVx2_ASAP7_75t_L g17084 ( 
.A(n_16685),
.Y(n_17084)
);

NOR3xp33_ASAP7_75t_SL g17085 ( 
.A(n_16720),
.B(n_2341),
.C(n_2342),
.Y(n_17085)
);

AND2x2_ASAP7_75t_L g17086 ( 
.A(n_16607),
.B(n_2343),
.Y(n_17086)
);

BUFx3_ASAP7_75t_L g17087 ( 
.A(n_16693),
.Y(n_17087)
);

NOR2xp33_ASAP7_75t_R g17088 ( 
.A(n_16726),
.B(n_2343),
.Y(n_17088)
);

HB1xp67_ASAP7_75t_L g17089 ( 
.A(n_16631),
.Y(n_17089)
);

INVx1_ASAP7_75t_L g17090 ( 
.A(n_16666),
.Y(n_17090)
);

AND2x2_ASAP7_75t_L g17091 ( 
.A(n_16570),
.B(n_2344),
.Y(n_17091)
);

INVx2_ASAP7_75t_L g17092 ( 
.A(n_16723),
.Y(n_17092)
);

AND2x4_ASAP7_75t_L g17093 ( 
.A(n_16842),
.B(n_2344),
.Y(n_17093)
);

NAND2xp5_ASAP7_75t_L g17094 ( 
.A(n_16740),
.B(n_2345),
.Y(n_17094)
);

CKINVDCx5p33_ASAP7_75t_R g17095 ( 
.A(n_16802),
.Y(n_17095)
);

INVx1_ASAP7_75t_L g17096 ( 
.A(n_16568),
.Y(n_17096)
);

OR2x6_ASAP7_75t_L g17097 ( 
.A(n_16870),
.B(n_2345),
.Y(n_17097)
);

CKINVDCx5p33_ASAP7_75t_R g17098 ( 
.A(n_16867),
.Y(n_17098)
);

CKINVDCx5p33_ASAP7_75t_R g17099 ( 
.A(n_16728),
.Y(n_17099)
);

NOR3xp33_ASAP7_75t_SL g17100 ( 
.A(n_16604),
.B(n_2346),
.C(n_2347),
.Y(n_17100)
);

AOI22xp33_ASAP7_75t_SL g17101 ( 
.A1(n_16538),
.A2(n_2348),
.B1(n_2346),
.B2(n_2347),
.Y(n_17101)
);

BUFx2_ASAP7_75t_L g17102 ( 
.A(n_16766),
.Y(n_17102)
);

AND2x2_ASAP7_75t_L g17103 ( 
.A(n_16767),
.B(n_2348),
.Y(n_17103)
);

BUFx2_ASAP7_75t_L g17104 ( 
.A(n_16558),
.Y(n_17104)
);

NOR3xp33_ASAP7_75t_SL g17105 ( 
.A(n_16629),
.B(n_2349),
.C(n_2350),
.Y(n_17105)
);

HB1xp67_ASAP7_75t_L g17106 ( 
.A(n_16659),
.Y(n_17106)
);

HB1xp67_ASAP7_75t_L g17107 ( 
.A(n_16662),
.Y(n_17107)
);

CKINVDCx20_ASAP7_75t_R g17108 ( 
.A(n_16843),
.Y(n_17108)
);

INVx2_ASAP7_75t_L g17109 ( 
.A(n_16831),
.Y(n_17109)
);

NOR2xp33_ASAP7_75t_L g17110 ( 
.A(n_16856),
.B(n_2349),
.Y(n_17110)
);

INVx1_ASAP7_75t_L g17111 ( 
.A(n_16569),
.Y(n_17111)
);

OR2x6_ASAP7_75t_L g17112 ( 
.A(n_16876),
.B(n_2350),
.Y(n_17112)
);

CKINVDCx5p33_ASAP7_75t_R g17113 ( 
.A(n_16881),
.Y(n_17113)
);

NOR2xp33_ASAP7_75t_R g17114 ( 
.A(n_16887),
.B(n_2351),
.Y(n_17114)
);

NAND2xp33_ASAP7_75t_R g17115 ( 
.A(n_16796),
.B(n_2351),
.Y(n_17115)
);

INVx1_ASAP7_75t_L g17116 ( 
.A(n_16575),
.Y(n_17116)
);

INVx1_ASAP7_75t_L g17117 ( 
.A(n_16577),
.Y(n_17117)
);

NAND2xp5_ASAP7_75t_L g17118 ( 
.A(n_16828),
.B(n_2352),
.Y(n_17118)
);

NOR3xp33_ASAP7_75t_SL g17119 ( 
.A(n_16864),
.B(n_2353),
.C(n_2354),
.Y(n_17119)
);

BUFx3_ASAP7_75t_L g17120 ( 
.A(n_16829),
.Y(n_17120)
);

NOR2xp33_ASAP7_75t_R g17121 ( 
.A(n_16815),
.B(n_2353),
.Y(n_17121)
);

INVx1_ASAP7_75t_L g17122 ( 
.A(n_16578),
.Y(n_17122)
);

HB1xp67_ASAP7_75t_L g17123 ( 
.A(n_16778),
.Y(n_17123)
);

CKINVDCx16_ASAP7_75t_R g17124 ( 
.A(n_16747),
.Y(n_17124)
);

HB1xp67_ASAP7_75t_L g17125 ( 
.A(n_16801),
.Y(n_17125)
);

CKINVDCx16_ASAP7_75t_R g17126 ( 
.A(n_16664),
.Y(n_17126)
);

INVx3_ASAP7_75t_L g17127 ( 
.A(n_16709),
.Y(n_17127)
);

OR2x2_ASAP7_75t_L g17128 ( 
.A(n_16544),
.B(n_2354),
.Y(n_17128)
);

AND2x2_ASAP7_75t_L g17129 ( 
.A(n_16780),
.B(n_2355),
.Y(n_17129)
);

XOR2xp5_ASAP7_75t_L g17130 ( 
.A(n_16830),
.B(n_2355),
.Y(n_17130)
);

OAI22xp33_ASAP7_75t_SL g17131 ( 
.A1(n_16730),
.A2(n_2358),
.B1(n_2356),
.B2(n_2357),
.Y(n_17131)
);

AND2x2_ASAP7_75t_L g17132 ( 
.A(n_16785),
.B(n_2356),
.Y(n_17132)
);

INVx2_ASAP7_75t_L g17133 ( 
.A(n_16756),
.Y(n_17133)
);

NOR2x1_ASAP7_75t_SL g17134 ( 
.A(n_16782),
.B(n_2357),
.Y(n_17134)
);

NOR2xp33_ASAP7_75t_L g17135 ( 
.A(n_16858),
.B(n_2358),
.Y(n_17135)
);

INVx3_ASAP7_75t_SL g17136 ( 
.A(n_16673),
.Y(n_17136)
);

BUFx2_ASAP7_75t_L g17137 ( 
.A(n_16576),
.Y(n_17137)
);

INVx1_ASAP7_75t_L g17138 ( 
.A(n_16583),
.Y(n_17138)
);

OR2x4_ASAP7_75t_L g17139 ( 
.A(n_16840),
.B(n_2359),
.Y(n_17139)
);

OR2x2_ASAP7_75t_L g17140 ( 
.A(n_16806),
.B(n_2360),
.Y(n_17140)
);

HB1xp67_ASAP7_75t_L g17141 ( 
.A(n_16799),
.Y(n_17141)
);

AND2x4_ASAP7_75t_SL g17142 ( 
.A(n_16627),
.B(n_2360),
.Y(n_17142)
);

INVx1_ASAP7_75t_L g17143 ( 
.A(n_16585),
.Y(n_17143)
);

CKINVDCx20_ASAP7_75t_R g17144 ( 
.A(n_16836),
.Y(n_17144)
);

CKINVDCx8_ASAP7_75t_R g17145 ( 
.A(n_16871),
.Y(n_17145)
);

NOR2xp33_ASAP7_75t_R g17146 ( 
.A(n_16847),
.B(n_2361),
.Y(n_17146)
);

INVx2_ASAP7_75t_L g17147 ( 
.A(n_16716),
.Y(n_17147)
);

INVx4_ASAP7_75t_SL g17148 ( 
.A(n_16851),
.Y(n_17148)
);

AOI22xp33_ASAP7_75t_L g17149 ( 
.A1(n_16652),
.A2(n_2363),
.B1(n_2361),
.B2(n_2362),
.Y(n_17149)
);

HB1xp67_ASAP7_75t_L g17150 ( 
.A(n_16784),
.Y(n_17150)
);

NAND2xp5_ASAP7_75t_L g17151 ( 
.A(n_16838),
.B(n_2362),
.Y(n_17151)
);

CKINVDCx16_ASAP7_75t_R g17152 ( 
.A(n_16882),
.Y(n_17152)
);

NAND3xp33_ASAP7_75t_L g17153 ( 
.A(n_16852),
.B(n_2363),
.C(n_2364),
.Y(n_17153)
);

OR2x2_ASAP7_75t_L g17154 ( 
.A(n_16841),
.B(n_2364),
.Y(n_17154)
);

AO31x2_ASAP7_75t_L g17155 ( 
.A1(n_16753),
.A2(n_2368),
.A3(n_2365),
.B(n_2366),
.Y(n_17155)
);

INVx1_ASAP7_75t_L g17156 ( 
.A(n_16588),
.Y(n_17156)
);

HB1xp67_ASAP7_75t_L g17157 ( 
.A(n_16807),
.Y(n_17157)
);

INVx1_ASAP7_75t_L g17158 ( 
.A(n_16594),
.Y(n_17158)
);

NOR2xp33_ASAP7_75t_L g17159 ( 
.A(n_16872),
.B(n_2366),
.Y(n_17159)
);

OR2x6_ASAP7_75t_L g17160 ( 
.A(n_16837),
.B(n_2368),
.Y(n_17160)
);

INVx1_ASAP7_75t_L g17161 ( 
.A(n_16598),
.Y(n_17161)
);

INVx2_ASAP7_75t_L g17162 ( 
.A(n_16733),
.Y(n_17162)
);

NAND2x1_ASAP7_75t_L g17163 ( 
.A(n_16708),
.B(n_2369),
.Y(n_17163)
);

HB1xp67_ASAP7_75t_L g17164 ( 
.A(n_16573),
.Y(n_17164)
);

OAI22xp5_ASAP7_75t_L g17165 ( 
.A1(n_16626),
.A2(n_2372),
.B1(n_2370),
.B2(n_2371),
.Y(n_17165)
);

AND2x2_ASAP7_75t_L g17166 ( 
.A(n_16642),
.B(n_2370),
.Y(n_17166)
);

NAND2xp33_ASAP7_75t_SL g17167 ( 
.A(n_16671),
.B(n_2371),
.Y(n_17167)
);

AOI22xp33_ASAP7_75t_L g17168 ( 
.A1(n_16641),
.A2(n_2374),
.B1(n_2372),
.B2(n_2373),
.Y(n_17168)
);

INVx1_ASAP7_75t_L g17169 ( 
.A(n_16601),
.Y(n_17169)
);

INVx2_ASAP7_75t_L g17170 ( 
.A(n_16702),
.Y(n_17170)
);

NAND2xp5_ASAP7_75t_L g17171 ( 
.A(n_16998),
.B(n_16791),
.Y(n_17171)
);

NOR2x1_ASAP7_75t_R g17172 ( 
.A(n_16910),
.B(n_16688),
.Y(n_17172)
);

INVx4_ASAP7_75t_L g17173 ( 
.A(n_16996),
.Y(n_17173)
);

BUFx2_ASAP7_75t_L g17174 ( 
.A(n_17011),
.Y(n_17174)
);

HB1xp67_ASAP7_75t_L g17175 ( 
.A(n_17102),
.Y(n_17175)
);

AND2x2_ASAP7_75t_L g17176 ( 
.A(n_16907),
.B(n_16645),
.Y(n_17176)
);

INVx2_ASAP7_75t_L g17177 ( 
.A(n_16919),
.Y(n_17177)
);

AND2x4_ASAP7_75t_L g17178 ( 
.A(n_16901),
.B(n_16647),
.Y(n_17178)
);

INVx2_ASAP7_75t_L g17179 ( 
.A(n_16941),
.Y(n_17179)
);

OR2x6_ASAP7_75t_L g17180 ( 
.A(n_16916),
.B(n_17060),
.Y(n_17180)
);

O2A1O1Ixp33_ASAP7_75t_SL g17181 ( 
.A1(n_16980),
.A2(n_16752),
.B(n_16750),
.C(n_16817),
.Y(n_17181)
);

AOI22xp33_ASAP7_75t_L g17182 ( 
.A1(n_16959),
.A2(n_16745),
.B1(n_16680),
.B2(n_16860),
.Y(n_17182)
);

OAI21x1_ASAP7_75t_L g17183 ( 
.A1(n_16902),
.A2(n_16590),
.B(n_16523),
.Y(n_17183)
);

AND2x4_ASAP7_75t_L g17184 ( 
.A(n_16911),
.B(n_16707),
.Y(n_17184)
);

OAI21xp5_ASAP7_75t_L g17185 ( 
.A1(n_16956),
.A2(n_16618),
.B(n_16533),
.Y(n_17185)
);

A2O1A1Ixp33_ASAP7_75t_L g17186 ( 
.A1(n_17018),
.A2(n_16774),
.B(n_16700),
.C(n_16731),
.Y(n_17186)
);

AND2x2_ASAP7_75t_L g17187 ( 
.A(n_16905),
.B(n_17054),
.Y(n_17187)
);

AOI21xp5_ASAP7_75t_SL g17188 ( 
.A1(n_16926),
.A2(n_16542),
.B(n_16595),
.Y(n_17188)
);

AO32x1_ASAP7_75t_L g17189 ( 
.A1(n_16922),
.A2(n_16755),
.A3(n_16536),
.B1(n_16539),
.B2(n_16532),
.Y(n_17189)
);

INVx1_ASAP7_75t_SL g17190 ( 
.A(n_16931),
.Y(n_17190)
);

INVx5_ASAP7_75t_L g17191 ( 
.A(n_16937),
.Y(n_17191)
);

AND4x1_ASAP7_75t_L g17192 ( 
.A(n_17025),
.B(n_16739),
.C(n_16734),
.D(n_16848),
.Y(n_17192)
);

AND2x4_ASAP7_75t_L g17193 ( 
.A(n_16940),
.B(n_16769),
.Y(n_17193)
);

AND2x4_ASAP7_75t_L g17194 ( 
.A(n_16914),
.B(n_16654),
.Y(n_17194)
);

OAI22xp5_ASAP7_75t_SL g17195 ( 
.A1(n_16903),
.A2(n_16850),
.B1(n_16891),
.B2(n_16878),
.Y(n_17195)
);

NAND2xp5_ASAP7_75t_L g17196 ( 
.A(n_16960),
.B(n_16861),
.Y(n_17196)
);

OR2x2_ASAP7_75t_L g17197 ( 
.A(n_16958),
.B(n_16875),
.Y(n_17197)
);

AND2x2_ASAP7_75t_L g17198 ( 
.A(n_16904),
.B(n_16812),
.Y(n_17198)
);

OA21x2_ASAP7_75t_L g17199 ( 
.A1(n_16936),
.A2(n_16524),
.B(n_16657),
.Y(n_17199)
);

AOI21xp5_ASAP7_75t_L g17200 ( 
.A1(n_16912),
.A2(n_16953),
.B(n_17051),
.Y(n_17200)
);

OAI21xp5_ASAP7_75t_L g17201 ( 
.A1(n_17056),
.A2(n_16623),
.B(n_16670),
.Y(n_17201)
);

INVx3_ASAP7_75t_L g17202 ( 
.A(n_17001),
.Y(n_17202)
);

OAI22xp5_ASAP7_75t_L g17203 ( 
.A1(n_17126),
.A2(n_16634),
.B1(n_16859),
.B2(n_16854),
.Y(n_17203)
);

AND2x2_ASAP7_75t_L g17204 ( 
.A(n_16939),
.B(n_16792),
.Y(n_17204)
);

A2O1A1Ixp33_ASAP7_75t_L g17205 ( 
.A1(n_16909),
.A2(n_16534),
.B(n_16725),
.C(n_16787),
.Y(n_17205)
);

AND2x2_ASAP7_75t_L g17206 ( 
.A(n_16915),
.B(n_16798),
.Y(n_17206)
);

OA21x2_ASAP7_75t_L g17207 ( 
.A1(n_17004),
.A2(n_16696),
.B(n_16772),
.Y(n_17207)
);

AND2x2_ASAP7_75t_L g17208 ( 
.A(n_16990),
.B(n_16800),
.Y(n_17208)
);

INVx2_ASAP7_75t_L g17209 ( 
.A(n_16941),
.Y(n_17209)
);

BUFx3_ASAP7_75t_L g17210 ( 
.A(n_16981),
.Y(n_17210)
);

INVx1_ASAP7_75t_L g17211 ( 
.A(n_16920),
.Y(n_17211)
);

HB1xp67_ASAP7_75t_L g17212 ( 
.A(n_17022),
.Y(n_17212)
);

NOR2x1_ASAP7_75t_SL g17213 ( 
.A(n_17160),
.B(n_16795),
.Y(n_17213)
);

OAI21xp5_ASAP7_75t_L g17214 ( 
.A1(n_16929),
.A2(n_16923),
.B(n_16918),
.Y(n_17214)
);

NAND2xp5_ASAP7_75t_SL g17215 ( 
.A(n_17072),
.B(n_16803),
.Y(n_17215)
);

AOI21xp5_ASAP7_75t_L g17216 ( 
.A1(n_16935),
.A2(n_16813),
.B(n_16810),
.Y(n_17216)
);

OAI22xp5_ASAP7_75t_SL g17217 ( 
.A1(n_17124),
.A2(n_16819),
.B1(n_16821),
.B2(n_16820),
.Y(n_17217)
);

OAI221xp5_ASAP7_75t_L g17218 ( 
.A1(n_16917),
.A2(n_17034),
.B1(n_16944),
.B2(n_16975),
.C(n_17100),
.Y(n_17218)
);

O2A1O1Ixp33_ASAP7_75t_L g17219 ( 
.A1(n_17165),
.A2(n_16790),
.B(n_16699),
.C(n_16681),
.Y(n_17219)
);

A2O1A1Ixp33_ASAP7_75t_L g17220 ( 
.A1(n_17085),
.A2(n_17099),
.B(n_17043),
.C(n_17040),
.Y(n_17220)
);

AO21x2_ASAP7_75t_L g17221 ( 
.A1(n_17164),
.A2(n_16675),
.B(n_16694),
.Y(n_17221)
);

AND2x2_ASAP7_75t_L g17222 ( 
.A(n_16913),
.B(n_16735),
.Y(n_17222)
);

OA21x2_ASAP7_75t_L g17223 ( 
.A1(n_16999),
.A2(n_16719),
.B(n_16622),
.Y(n_17223)
);

AND2x4_ASAP7_75t_L g17224 ( 
.A(n_16938),
.B(n_16736),
.Y(n_17224)
);

INVxp67_ASAP7_75t_SL g17225 ( 
.A(n_16965),
.Y(n_17225)
);

OA21x2_ASAP7_75t_L g17226 ( 
.A1(n_16969),
.A2(n_16639),
.B(n_16655),
.Y(n_17226)
);

NOR2xp33_ASAP7_75t_L g17227 ( 
.A(n_17027),
.B(n_16665),
.Y(n_17227)
);

OAI221xp5_ASAP7_75t_L g17228 ( 
.A1(n_16975),
.A2(n_16845),
.B1(n_16683),
.B2(n_16704),
.C(n_16703),
.Y(n_17228)
);

INVx4_ASAP7_75t_L g17229 ( 
.A(n_16924),
.Y(n_17229)
);

INVx2_ASAP7_75t_L g17230 ( 
.A(n_16977),
.Y(n_17230)
);

INVx5_ASAP7_75t_L g17231 ( 
.A(n_16997),
.Y(n_17231)
);

AND2x2_ASAP7_75t_SL g17232 ( 
.A(n_17152),
.B(n_16738),
.Y(n_17232)
);

OA21x2_ASAP7_75t_L g17233 ( 
.A1(n_16951),
.A2(n_16656),
.B(n_16690),
.Y(n_17233)
);

AO21x2_ASAP7_75t_L g17234 ( 
.A1(n_17019),
.A2(n_17006),
.B(n_16972),
.Y(n_17234)
);

OAI22xp5_ASAP7_75t_L g17235 ( 
.A1(n_17008),
.A2(n_16808),
.B1(n_16743),
.B2(n_16706),
.Y(n_17235)
);

AND2x4_ASAP7_75t_L g17236 ( 
.A(n_16921),
.B(n_16925),
.Y(n_17236)
);

HB1xp67_ASAP7_75t_L g17237 ( 
.A(n_16900),
.Y(n_17237)
);

INVx1_ASAP7_75t_L g17238 ( 
.A(n_17141),
.Y(n_17238)
);

OAI21xp5_ASAP7_75t_L g17239 ( 
.A1(n_17058),
.A2(n_16721),
.B(n_16717),
.Y(n_17239)
);

AND2x2_ASAP7_75t_L g17240 ( 
.A(n_16968),
.B(n_16724),
.Y(n_17240)
);

NOR2xp33_ASAP7_75t_L g17241 ( 
.A(n_16977),
.B(n_16727),
.Y(n_17241)
);

NAND2xp5_ASAP7_75t_L g17242 ( 
.A(n_17134),
.B(n_16729),
.Y(n_17242)
);

A2O1A1Ixp33_ASAP7_75t_L g17243 ( 
.A1(n_17039),
.A2(n_16608),
.B(n_16612),
.C(n_16605),
.Y(n_17243)
);

OA21x2_ASAP7_75t_L g17244 ( 
.A1(n_17020),
.A2(n_16742),
.B(n_16620),
.Y(n_17244)
);

AOI22xp5_ASAP7_75t_L g17245 ( 
.A1(n_16973),
.A2(n_16661),
.B1(n_16621),
.B2(n_16624),
.Y(n_17245)
);

NOR2xp33_ASAP7_75t_L g17246 ( 
.A(n_16945),
.B(n_16613),
.Y(n_17246)
);

AND2x6_ASAP7_75t_L g17247 ( 
.A(n_17028),
.B(n_16625),
.Y(n_17247)
);

OR2x2_ASAP7_75t_L g17248 ( 
.A(n_16974),
.B(n_17076),
.Y(n_17248)
);

AND2x2_ASAP7_75t_L g17249 ( 
.A(n_16949),
.B(n_16628),
.Y(n_17249)
);

AND2x2_ASAP7_75t_L g17250 ( 
.A(n_17012),
.B(n_16633),
.Y(n_17250)
);

BUFx2_ASAP7_75t_L g17251 ( 
.A(n_16994),
.Y(n_17251)
);

AND2x2_ASAP7_75t_L g17252 ( 
.A(n_16964),
.B(n_16635),
.Y(n_17252)
);

AND2x2_ASAP7_75t_L g17253 ( 
.A(n_16989),
.B(n_16636),
.Y(n_17253)
);

AND2x2_ASAP7_75t_L g17254 ( 
.A(n_16962),
.B(n_16637),
.Y(n_17254)
);

AOI221xp5_ASAP7_75t_L g17255 ( 
.A1(n_16934),
.A2(n_16653),
.B1(n_16638),
.B2(n_16851),
.C(n_16888),
.Y(n_17255)
);

BUFx3_ASAP7_75t_L g17256 ( 
.A(n_16997),
.Y(n_17256)
);

AO32x2_ASAP7_75t_L g17257 ( 
.A1(n_16988),
.A2(n_17115),
.A3(n_17148),
.B1(n_16995),
.B2(n_17144),
.Y(n_17257)
);

AO32x2_ASAP7_75t_L g17258 ( 
.A1(n_17005),
.A2(n_16888),
.A3(n_2375),
.B1(n_2373),
.B2(n_2374),
.Y(n_17258)
);

BUFx12f_ASAP7_75t_L g17259 ( 
.A(n_16997),
.Y(n_17259)
);

AOI221x1_ASAP7_75t_SL g17260 ( 
.A1(n_16930),
.A2(n_17078),
.B1(n_17082),
.B2(n_17092),
.C(n_17059),
.Y(n_17260)
);

NAND2xp5_ASAP7_75t_L g17261 ( 
.A(n_17033),
.B(n_2376),
.Y(n_17261)
);

AO21x2_ASAP7_75t_L g17262 ( 
.A1(n_17047),
.A2(n_2377),
.B(n_2378),
.Y(n_17262)
);

NAND2xp5_ASAP7_75t_L g17263 ( 
.A(n_16932),
.B(n_2377),
.Y(n_17263)
);

AND2x4_ASAP7_75t_SL g17264 ( 
.A(n_17041),
.B(n_2378),
.Y(n_17264)
);

INVx1_ASAP7_75t_L g17265 ( 
.A(n_17123),
.Y(n_17265)
);

O2A1O1Ixp5_ASAP7_75t_SL g17266 ( 
.A1(n_16943),
.A2(n_2381),
.B(n_2379),
.C(n_2380),
.Y(n_17266)
);

OR2x6_ASAP7_75t_L g17267 ( 
.A(n_17017),
.B(n_2379),
.Y(n_17267)
);

AO32x2_ASAP7_75t_L g17268 ( 
.A1(n_16954),
.A2(n_2383),
.A3(n_2380),
.B1(n_2382),
.B2(n_2384),
.Y(n_17268)
);

AND2x4_ASAP7_75t_L g17269 ( 
.A(n_16950),
.B(n_17066),
.Y(n_17269)
);

AND2x2_ASAP7_75t_L g17270 ( 
.A(n_17003),
.B(n_17136),
.Y(n_17270)
);

AND2x2_ASAP7_75t_L g17271 ( 
.A(n_17065),
.B(n_2382),
.Y(n_17271)
);

OR2x2_ASAP7_75t_L g17272 ( 
.A(n_17137),
.B(n_2383),
.Y(n_17272)
);

NOR4xp25_ASAP7_75t_SL g17273 ( 
.A(n_16963),
.B(n_2386),
.C(n_2384),
.D(n_2385),
.Y(n_17273)
);

A2O1A1Ixp33_ASAP7_75t_L g17274 ( 
.A1(n_17105),
.A2(n_2387),
.B(n_2385),
.C(n_2386),
.Y(n_17274)
);

OA21x2_ASAP7_75t_L g17275 ( 
.A1(n_16992),
.A2(n_2388),
.B(n_2389),
.Y(n_17275)
);

OAI221xp5_ASAP7_75t_L g17276 ( 
.A1(n_17145),
.A2(n_2390),
.B1(n_2388),
.B2(n_2389),
.C(n_2391),
.Y(n_17276)
);

NAND3xp33_ASAP7_75t_L g17277 ( 
.A(n_17070),
.B(n_2390),
.C(n_2391),
.Y(n_17277)
);

AND2x4_ASAP7_75t_L g17278 ( 
.A(n_17068),
.B(n_17087),
.Y(n_17278)
);

OR2x2_ASAP7_75t_L g17279 ( 
.A(n_17002),
.B(n_2392),
.Y(n_17279)
);

HB1xp67_ASAP7_75t_L g17280 ( 
.A(n_17125),
.Y(n_17280)
);

AO21x2_ASAP7_75t_L g17281 ( 
.A1(n_17015),
.A2(n_2392),
.B(n_2393),
.Y(n_17281)
);

NAND2xp5_ASAP7_75t_L g17282 ( 
.A(n_17023),
.B(n_2393),
.Y(n_17282)
);

AND2x2_ASAP7_75t_L g17283 ( 
.A(n_17077),
.B(n_2394),
.Y(n_17283)
);

INVx2_ASAP7_75t_L g17284 ( 
.A(n_17142),
.Y(n_17284)
);

NAND2xp5_ASAP7_75t_L g17285 ( 
.A(n_17091),
.B(n_2394),
.Y(n_17285)
);

OR2x2_ASAP7_75t_L g17286 ( 
.A(n_17104),
.B(n_2395),
.Y(n_17286)
);

BUFx6f_ASAP7_75t_L g17287 ( 
.A(n_16967),
.Y(n_17287)
);

AND2x4_ASAP7_75t_L g17288 ( 
.A(n_17014),
.B(n_2395),
.Y(n_17288)
);

INVx2_ASAP7_75t_L g17289 ( 
.A(n_17108),
.Y(n_17289)
);

OR2x6_ASAP7_75t_L g17290 ( 
.A(n_17073),
.B(n_2396),
.Y(n_17290)
);

A2O1A1Ixp33_ASAP7_75t_L g17291 ( 
.A1(n_17167),
.A2(n_2398),
.B(n_2396),
.C(n_2397),
.Y(n_17291)
);

INVx2_ASAP7_75t_L g17292 ( 
.A(n_16976),
.Y(n_17292)
);

OAI211xp5_ASAP7_75t_L g17293 ( 
.A1(n_17101),
.A2(n_2399),
.B(n_2397),
.C(n_2398),
.Y(n_17293)
);

AND2x2_ASAP7_75t_L g17294 ( 
.A(n_16983),
.B(n_2399),
.Y(n_17294)
);

BUFx3_ASAP7_75t_L g17295 ( 
.A(n_17007),
.Y(n_17295)
);

NOR2x1_ASAP7_75t_SL g17296 ( 
.A(n_17160),
.B(n_2400),
.Y(n_17296)
);

AND2x4_ASAP7_75t_L g17297 ( 
.A(n_17045),
.B(n_2400),
.Y(n_17297)
);

AND2x2_ASAP7_75t_L g17298 ( 
.A(n_17055),
.B(n_2401),
.Y(n_17298)
);

NOR2xp33_ASAP7_75t_L g17299 ( 
.A(n_17098),
.B(n_2401),
.Y(n_17299)
);

NAND2xp5_ASAP7_75t_L g17300 ( 
.A(n_16961),
.B(n_2402),
.Y(n_17300)
);

NAND2xp5_ASAP7_75t_L g17301 ( 
.A(n_16955),
.B(n_2402),
.Y(n_17301)
);

NOR2x1_ASAP7_75t_SL g17302 ( 
.A(n_17035),
.B(n_2403),
.Y(n_17302)
);

AND2x2_ASAP7_75t_L g17303 ( 
.A(n_16928),
.B(n_17029),
.Y(n_17303)
);

AND2x2_ASAP7_75t_L g17304 ( 
.A(n_17067),
.B(n_2403),
.Y(n_17304)
);

AND2x2_ASAP7_75t_L g17305 ( 
.A(n_17062),
.B(n_2404),
.Y(n_17305)
);

INVx2_ASAP7_75t_SL g17306 ( 
.A(n_17000),
.Y(n_17306)
);

INVx2_ASAP7_75t_L g17307 ( 
.A(n_17035),
.Y(n_17307)
);

INVx2_ASAP7_75t_L g17308 ( 
.A(n_17071),
.Y(n_17308)
);

OAI21xp5_ASAP7_75t_L g17309 ( 
.A1(n_16906),
.A2(n_2405),
.B(n_2406),
.Y(n_17309)
);

AND2x2_ASAP7_75t_L g17310 ( 
.A(n_17127),
.B(n_2405),
.Y(n_17310)
);

OA21x2_ASAP7_75t_L g17311 ( 
.A1(n_16952),
.A2(n_2406),
.B(n_2407),
.Y(n_17311)
);

NAND2xp5_ASAP7_75t_L g17312 ( 
.A(n_16955),
.B(n_2407),
.Y(n_17312)
);

BUFx12f_ASAP7_75t_L g17313 ( 
.A(n_17113),
.Y(n_17313)
);

NOR2xp33_ASAP7_75t_L g17314 ( 
.A(n_17095),
.B(n_17139),
.Y(n_17314)
);

NAND2xp5_ASAP7_75t_L g17315 ( 
.A(n_16933),
.B(n_2408),
.Y(n_17315)
);

INVx1_ASAP7_75t_L g17316 ( 
.A(n_17150),
.Y(n_17316)
);

INVx1_ASAP7_75t_L g17317 ( 
.A(n_17032),
.Y(n_17317)
);

OA21x2_ASAP7_75t_L g17318 ( 
.A1(n_17133),
.A2(n_2409),
.B(n_2410),
.Y(n_17318)
);

INVx1_ASAP7_75t_L g17319 ( 
.A(n_17089),
.Y(n_17319)
);

NOR2xp33_ASAP7_75t_L g17320 ( 
.A(n_17042),
.B(n_17140),
.Y(n_17320)
);

OA21x2_ASAP7_75t_L g17321 ( 
.A1(n_17147),
.A2(n_2411),
.B(n_2412),
.Y(n_17321)
);

BUFx2_ASAP7_75t_L g17322 ( 
.A(n_16947),
.Y(n_17322)
);

AND2x4_ASAP7_75t_L g17323 ( 
.A(n_17120),
.B(n_2411),
.Y(n_17323)
);

BUFx4f_ASAP7_75t_SL g17324 ( 
.A(n_16966),
.Y(n_17324)
);

INVx1_ASAP7_75t_L g17325 ( 
.A(n_17106),
.Y(n_17325)
);

AND2x2_ASAP7_75t_L g17326 ( 
.A(n_17069),
.B(n_2412),
.Y(n_17326)
);

A2O1A1Ixp33_ASAP7_75t_L g17327 ( 
.A1(n_17119),
.A2(n_2415),
.B(n_2413),
.C(n_2414),
.Y(n_17327)
);

NAND2xp5_ASAP7_75t_SL g17328 ( 
.A(n_17131),
.B(n_2413),
.Y(n_17328)
);

NOR2xp33_ASAP7_75t_L g17329 ( 
.A(n_17128),
.B(n_2414),
.Y(n_17329)
);

A2O1A1Ixp33_ASAP7_75t_L g17330 ( 
.A1(n_17064),
.A2(n_2417),
.B(n_2415),
.C(n_2416),
.Y(n_17330)
);

OR2x2_ASAP7_75t_L g17331 ( 
.A(n_17109),
.B(n_2416),
.Y(n_17331)
);

INVxp67_ASAP7_75t_L g17332 ( 
.A(n_17038),
.Y(n_17332)
);

BUFx12f_ASAP7_75t_L g17333 ( 
.A(n_17030),
.Y(n_17333)
);

NOR2xp33_ASAP7_75t_L g17334 ( 
.A(n_17118),
.B(n_2417),
.Y(n_17334)
);

INVx1_ASAP7_75t_L g17335 ( 
.A(n_17107),
.Y(n_17335)
);

O2A1O1Ixp33_ASAP7_75t_L g17336 ( 
.A1(n_17008),
.A2(n_2420),
.B(n_2418),
.C(n_2419),
.Y(n_17336)
);

AND2x2_ASAP7_75t_L g17337 ( 
.A(n_17074),
.B(n_2418),
.Y(n_17337)
);

INVx1_ASAP7_75t_L g17338 ( 
.A(n_17157),
.Y(n_17338)
);

A2O1A1Ixp33_ASAP7_75t_L g17339 ( 
.A1(n_17153),
.A2(n_17163),
.B(n_16979),
.C(n_17080),
.Y(n_17339)
);

AOI22xp5_ASAP7_75t_SL g17340 ( 
.A1(n_17130),
.A2(n_2421),
.B1(n_2419),
.B2(n_2420),
.Y(n_17340)
);

INVx1_ASAP7_75t_L g17341 ( 
.A(n_16948),
.Y(n_17341)
);

INVx3_ASAP7_75t_L g17342 ( 
.A(n_17093),
.Y(n_17342)
);

AND2x2_ASAP7_75t_L g17343 ( 
.A(n_17079),
.B(n_2422),
.Y(n_17343)
);

OR2x2_ASAP7_75t_L g17344 ( 
.A(n_16933),
.B(n_2422),
.Y(n_17344)
);

OAI21xp5_ASAP7_75t_L g17345 ( 
.A1(n_16906),
.A2(n_2423),
.B(n_2424),
.Y(n_17345)
);

OR2x2_ASAP7_75t_L g17346 ( 
.A(n_17084),
.B(n_2423),
.Y(n_17346)
);

INVxp67_ASAP7_75t_L g17347 ( 
.A(n_17063),
.Y(n_17347)
);

INVx1_ASAP7_75t_L g17348 ( 
.A(n_16970),
.Y(n_17348)
);

OR2x2_ASAP7_75t_L g17349 ( 
.A(n_16908),
.B(n_2424),
.Y(n_17349)
);

O2A1O1Ixp5_ASAP7_75t_L g17350 ( 
.A1(n_17162),
.A2(n_2427),
.B(n_2425),
.C(n_2426),
.Y(n_17350)
);

CKINVDCx5p33_ASAP7_75t_R g17351 ( 
.A(n_16946),
.Y(n_17351)
);

AOI21xp5_ASAP7_75t_L g17352 ( 
.A1(n_16908),
.A2(n_2426),
.B(n_2427),
.Y(n_17352)
);

AND2x2_ASAP7_75t_L g17353 ( 
.A(n_17036),
.B(n_2428),
.Y(n_17353)
);

NOR2xp67_ASAP7_75t_L g17354 ( 
.A(n_17170),
.B(n_2428),
.Y(n_17354)
);

NOR2x1_ASAP7_75t_SL g17355 ( 
.A(n_17071),
.B(n_2429),
.Y(n_17355)
);

OAI21xp5_ASAP7_75t_L g17356 ( 
.A1(n_16927),
.A2(n_2429),
.B(n_2430),
.Y(n_17356)
);

AND2x2_ASAP7_75t_L g17357 ( 
.A(n_17021),
.B(n_2430),
.Y(n_17357)
);

BUFx12f_ASAP7_75t_L g17358 ( 
.A(n_17024),
.Y(n_17358)
);

NAND2xp5_ASAP7_75t_L g17359 ( 
.A(n_17103),
.B(n_2431),
.Y(n_17359)
);

OAI21xp5_ASAP7_75t_L g17360 ( 
.A1(n_16927),
.A2(n_2432),
.B(n_2433),
.Y(n_17360)
);

AND2x2_ASAP7_75t_L g17361 ( 
.A(n_16957),
.B(n_2432),
.Y(n_17361)
);

AND2x4_ASAP7_75t_L g17362 ( 
.A(n_16993),
.B(n_2434),
.Y(n_17362)
);

INVx1_ASAP7_75t_L g17363 ( 
.A(n_16971),
.Y(n_17363)
);

NAND4xp25_ASAP7_75t_L g17364 ( 
.A(n_17061),
.B(n_17075),
.C(n_17052),
.D(n_17013),
.Y(n_17364)
);

AOI22xp5_ASAP7_75t_L g17365 ( 
.A1(n_17135),
.A2(n_2436),
.B1(n_2434),
.B2(n_2435),
.Y(n_17365)
);

AOI21xp5_ASAP7_75t_L g17366 ( 
.A1(n_17159),
.A2(n_2436),
.B(n_2437),
.Y(n_17366)
);

O2A1O1Ixp33_ASAP7_75t_SL g17367 ( 
.A1(n_17049),
.A2(n_2440),
.B(n_2438),
.C(n_2439),
.Y(n_17367)
);

NOR2x1_ASAP7_75t_SL g17368 ( 
.A(n_17073),
.B(n_2438),
.Y(n_17368)
);

NOR2xp33_ASAP7_75t_L g17369 ( 
.A(n_17151),
.B(n_2439),
.Y(n_17369)
);

AND2x2_ASAP7_75t_L g17370 ( 
.A(n_17129),
.B(n_2440),
.Y(n_17370)
);

NAND2xp5_ASAP7_75t_L g17371 ( 
.A(n_17110),
.B(n_2441),
.Y(n_17371)
);

AND2x4_ASAP7_75t_L g17372 ( 
.A(n_16986),
.B(n_2441),
.Y(n_17372)
);

HB1xp67_ASAP7_75t_L g17373 ( 
.A(n_17097),
.Y(n_17373)
);

HB1xp67_ASAP7_75t_L g17374 ( 
.A(n_17097),
.Y(n_17374)
);

OAI21xp5_ASAP7_75t_L g17375 ( 
.A1(n_17168),
.A2(n_2442),
.B(n_2443),
.Y(n_17375)
);

BUFx12f_ASAP7_75t_L g17376 ( 
.A(n_17037),
.Y(n_17376)
);

INVx1_ASAP7_75t_L g17377 ( 
.A(n_17237),
.Y(n_17377)
);

AOI221xp5_ASAP7_75t_L g17378 ( 
.A1(n_17188),
.A2(n_16982),
.B1(n_17009),
.B2(n_16987),
.C(n_16985),
.Y(n_17378)
);

INVx1_ASAP7_75t_L g17379 ( 
.A(n_17280),
.Y(n_17379)
);

NAND2xp5_ASAP7_75t_L g17380 ( 
.A(n_17332),
.B(n_17132),
.Y(n_17380)
);

INVx1_ASAP7_75t_L g17381 ( 
.A(n_17175),
.Y(n_17381)
);

HB1xp67_ASAP7_75t_L g17382 ( 
.A(n_17322),
.Y(n_17382)
);

BUFx3_ASAP7_75t_L g17383 ( 
.A(n_17313),
.Y(n_17383)
);

BUFx3_ASAP7_75t_L g17384 ( 
.A(n_17191),
.Y(n_17384)
);

NAND2xp5_ASAP7_75t_L g17385 ( 
.A(n_17347),
.B(n_17247),
.Y(n_17385)
);

INVx1_ASAP7_75t_L g17386 ( 
.A(n_17265),
.Y(n_17386)
);

NAND2xp5_ASAP7_75t_L g17387 ( 
.A(n_17247),
.B(n_17050),
.Y(n_17387)
);

AND2x2_ASAP7_75t_L g17388 ( 
.A(n_17187),
.B(n_17086),
.Y(n_17388)
);

AND2x2_ASAP7_75t_L g17389 ( 
.A(n_17191),
.B(n_17112),
.Y(n_17389)
);

INVx2_ASAP7_75t_L g17390 ( 
.A(n_17180),
.Y(n_17390)
);

AO21x2_ASAP7_75t_L g17391 ( 
.A1(n_17301),
.A2(n_16984),
.B(n_16978),
.Y(n_17391)
);

INVx2_ASAP7_75t_L g17392 ( 
.A(n_17180),
.Y(n_17392)
);

HB1xp67_ASAP7_75t_L g17393 ( 
.A(n_17231),
.Y(n_17393)
);

INVx3_ASAP7_75t_L g17394 ( 
.A(n_17173),
.Y(n_17394)
);

INVx2_ASAP7_75t_SL g17395 ( 
.A(n_17231),
.Y(n_17395)
);

INVx2_ASAP7_75t_L g17396 ( 
.A(n_17295),
.Y(n_17396)
);

INVx2_ASAP7_75t_L g17397 ( 
.A(n_17202),
.Y(n_17397)
);

AND2x2_ASAP7_75t_L g17398 ( 
.A(n_17190),
.B(n_17251),
.Y(n_17398)
);

INVx1_ASAP7_75t_L g17399 ( 
.A(n_17338),
.Y(n_17399)
);

INVx2_ASAP7_75t_L g17400 ( 
.A(n_17210),
.Y(n_17400)
);

INVx5_ASAP7_75t_L g17401 ( 
.A(n_17259),
.Y(n_17401)
);

INVx1_ASAP7_75t_L g17402 ( 
.A(n_17211),
.Y(n_17402)
);

BUFx3_ASAP7_75t_L g17403 ( 
.A(n_17333),
.Y(n_17403)
);

INVx2_ASAP7_75t_L g17404 ( 
.A(n_17256),
.Y(n_17404)
);

INVx3_ASAP7_75t_L g17405 ( 
.A(n_17278),
.Y(n_17405)
);

NAND2xp5_ASAP7_75t_L g17406 ( 
.A(n_17247),
.B(n_17166),
.Y(n_17406)
);

AND2x2_ASAP7_75t_L g17407 ( 
.A(n_17174),
.B(n_17112),
.Y(n_17407)
);

AOI22xp33_ASAP7_75t_L g17408 ( 
.A1(n_17195),
.A2(n_17090),
.B1(n_17114),
.B2(n_17016),
.Y(n_17408)
);

HB1xp67_ASAP7_75t_L g17409 ( 
.A(n_17373),
.Y(n_17409)
);

INVx2_ASAP7_75t_L g17410 ( 
.A(n_17287),
.Y(n_17410)
);

NOR2xp67_ASAP7_75t_L g17411 ( 
.A(n_17212),
.B(n_17306),
.Y(n_17411)
);

OR2x2_ASAP7_75t_L g17412 ( 
.A(n_17364),
.B(n_17154),
.Y(n_17412)
);

AND2x4_ASAP7_75t_L g17413 ( 
.A(n_17225),
.B(n_17046),
.Y(n_17413)
);

NAND2xp5_ASAP7_75t_L g17414 ( 
.A(n_17289),
.B(n_17010),
.Y(n_17414)
);

AOI322xp5_ASAP7_75t_L g17415 ( 
.A1(n_17312),
.A2(n_17149),
.A3(n_17031),
.B1(n_17053),
.B2(n_17057),
.C1(n_17116),
.C2(n_17111),
.Y(n_17415)
);

INVx2_ASAP7_75t_L g17416 ( 
.A(n_17287),
.Y(n_17416)
);

HB1xp67_ASAP7_75t_L g17417 ( 
.A(n_17374),
.Y(n_17417)
);

OR2x2_ASAP7_75t_L g17418 ( 
.A(n_17171),
.B(n_17096),
.Y(n_17418)
);

BUFx2_ASAP7_75t_L g17419 ( 
.A(n_17358),
.Y(n_17419)
);

AND2x2_ASAP7_75t_L g17420 ( 
.A(n_17232),
.B(n_17081),
.Y(n_17420)
);

AND2x2_ASAP7_75t_L g17421 ( 
.A(n_17198),
.B(n_16942),
.Y(n_17421)
);

INVx2_ASAP7_75t_L g17422 ( 
.A(n_17270),
.Y(n_17422)
);

INVx1_ASAP7_75t_L g17423 ( 
.A(n_17317),
.Y(n_17423)
);

INVx3_ASAP7_75t_L g17424 ( 
.A(n_17184),
.Y(n_17424)
);

INVx2_ASAP7_75t_L g17425 ( 
.A(n_17324),
.Y(n_17425)
);

OAI31xp33_ASAP7_75t_SL g17426 ( 
.A1(n_17214),
.A2(n_17122),
.A3(n_17138),
.B(n_17117),
.Y(n_17426)
);

INVx1_ASAP7_75t_L g17427 ( 
.A(n_17319),
.Y(n_17427)
);

AND2x2_ASAP7_75t_L g17428 ( 
.A(n_17176),
.B(n_17088),
.Y(n_17428)
);

OAI221xp5_ASAP7_75t_L g17429 ( 
.A1(n_17218),
.A2(n_17156),
.B1(n_17161),
.B2(n_17158),
.C(n_17143),
.Y(n_17429)
);

INVxp67_ASAP7_75t_SL g17430 ( 
.A(n_17302),
.Y(n_17430)
);

OR2x2_ASAP7_75t_L g17431 ( 
.A(n_17307),
.B(n_17169),
.Y(n_17431)
);

AND2x2_ASAP7_75t_L g17432 ( 
.A(n_17308),
.B(n_17044),
.Y(n_17432)
);

NAND2xp5_ASAP7_75t_L g17433 ( 
.A(n_17262),
.B(n_17010),
.Y(n_17433)
);

AND2x2_ASAP7_75t_L g17434 ( 
.A(n_17177),
.B(n_17342),
.Y(n_17434)
);

INVx2_ASAP7_75t_L g17435 ( 
.A(n_17355),
.Y(n_17435)
);

INVx2_ASAP7_75t_SL g17436 ( 
.A(n_17264),
.Y(n_17436)
);

AND2x2_ASAP7_75t_L g17437 ( 
.A(n_17284),
.B(n_17146),
.Y(n_17437)
);

NOR2x1_ASAP7_75t_SL g17438 ( 
.A(n_17267),
.B(n_17094),
.Y(n_17438)
);

AND2x2_ASAP7_75t_L g17439 ( 
.A(n_17269),
.B(n_17083),
.Y(n_17439)
);

BUFx3_ASAP7_75t_L g17440 ( 
.A(n_17376),
.Y(n_17440)
);

INVx1_ASAP7_75t_L g17441 ( 
.A(n_17325),
.Y(n_17441)
);

AND2x2_ASAP7_75t_L g17442 ( 
.A(n_17230),
.B(n_17121),
.Y(n_17442)
);

INVx1_ASAP7_75t_L g17443 ( 
.A(n_17335),
.Y(n_17443)
);

INVx2_ASAP7_75t_L g17444 ( 
.A(n_17368),
.Y(n_17444)
);

INVx1_ASAP7_75t_L g17445 ( 
.A(n_17238),
.Y(n_17445)
);

HB1xp67_ASAP7_75t_L g17446 ( 
.A(n_17233),
.Y(n_17446)
);

INVx8_ASAP7_75t_L g17447 ( 
.A(n_17351),
.Y(n_17447)
);

INVx2_ASAP7_75t_L g17448 ( 
.A(n_17213),
.Y(n_17448)
);

AND2x2_ASAP7_75t_SL g17449 ( 
.A(n_17344),
.B(n_17315),
.Y(n_17449)
);

INVx1_ASAP7_75t_L g17450 ( 
.A(n_17286),
.Y(n_17450)
);

AND2x2_ASAP7_75t_L g17451 ( 
.A(n_17303),
.B(n_17179),
.Y(n_17451)
);

INVx2_ASAP7_75t_L g17452 ( 
.A(n_17296),
.Y(n_17452)
);

BUFx3_ASAP7_75t_L g17453 ( 
.A(n_17178),
.Y(n_17453)
);

AND2x4_ASAP7_75t_L g17454 ( 
.A(n_17209),
.B(n_17155),
.Y(n_17454)
);

INVx4_ASAP7_75t_L g17455 ( 
.A(n_17229),
.Y(n_17455)
);

INVx1_ASAP7_75t_L g17456 ( 
.A(n_17208),
.Y(n_17456)
);

NAND2xp5_ASAP7_75t_L g17457 ( 
.A(n_17281),
.B(n_17026),
.Y(n_17457)
);

NAND2xp5_ASAP7_75t_L g17458 ( 
.A(n_17245),
.B(n_17026),
.Y(n_17458)
);

AND2x2_ASAP7_75t_L g17459 ( 
.A(n_17206),
.B(n_17155),
.Y(n_17459)
);

OR2x2_ASAP7_75t_L g17460 ( 
.A(n_17248),
.B(n_16991),
.Y(n_17460)
);

INVx1_ASAP7_75t_L g17461 ( 
.A(n_17331),
.Y(n_17461)
);

INVx1_ASAP7_75t_L g17462 ( 
.A(n_17316),
.Y(n_17462)
);

NAND2xp5_ASAP7_75t_L g17463 ( 
.A(n_17193),
.B(n_17220),
.Y(n_17463)
);

BUFx2_ASAP7_75t_L g17464 ( 
.A(n_17257),
.Y(n_17464)
);

INVx1_ASAP7_75t_L g17465 ( 
.A(n_17346),
.Y(n_17465)
);

INVx1_ASAP7_75t_L g17466 ( 
.A(n_17326),
.Y(n_17466)
);

INVx1_ASAP7_75t_L g17467 ( 
.A(n_17337),
.Y(n_17467)
);

INVx1_ASAP7_75t_L g17468 ( 
.A(n_17343),
.Y(n_17468)
);

AND2x2_ASAP7_75t_L g17469 ( 
.A(n_17236),
.B(n_16991),
.Y(n_17469)
);

HB1xp67_ASAP7_75t_L g17470 ( 
.A(n_17354),
.Y(n_17470)
);

INVx2_ASAP7_75t_L g17471 ( 
.A(n_17267),
.Y(n_17471)
);

AO21x2_ASAP7_75t_L g17472 ( 
.A1(n_17200),
.A2(n_17263),
.B(n_17352),
.Y(n_17472)
);

INVx1_ASAP7_75t_L g17473 ( 
.A(n_17298),
.Y(n_17473)
);

CKINVDCx16_ASAP7_75t_R g17474 ( 
.A(n_17217),
.Y(n_17474)
);

INVxp67_ASAP7_75t_SL g17475 ( 
.A(n_17172),
.Y(n_17475)
);

AND2x2_ASAP7_75t_L g17476 ( 
.A(n_17252),
.B(n_17048),
.Y(n_17476)
);

AND2x2_ASAP7_75t_L g17477 ( 
.A(n_17257),
.B(n_2442),
.Y(n_17477)
);

OA21x2_ASAP7_75t_L g17478 ( 
.A1(n_17185),
.A2(n_2443),
.B(n_2444),
.Y(n_17478)
);

BUFx3_ASAP7_75t_L g17479 ( 
.A(n_17224),
.Y(n_17479)
);

AND2x2_ASAP7_75t_L g17480 ( 
.A(n_17204),
.B(n_2444),
.Y(n_17480)
);

INVx2_ASAP7_75t_SL g17481 ( 
.A(n_17253),
.Y(n_17481)
);

INVx1_ASAP7_75t_L g17482 ( 
.A(n_17304),
.Y(n_17482)
);

OR2x2_ASAP7_75t_L g17483 ( 
.A(n_17197),
.B(n_2445),
.Y(n_17483)
);

INVx3_ASAP7_75t_L g17484 ( 
.A(n_17297),
.Y(n_17484)
);

AND2x2_ASAP7_75t_L g17485 ( 
.A(n_17240),
.B(n_2445),
.Y(n_17485)
);

AND2x2_ASAP7_75t_SL g17486 ( 
.A(n_17199),
.B(n_2446),
.Y(n_17486)
);

INVx1_ASAP7_75t_L g17487 ( 
.A(n_17282),
.Y(n_17487)
);

INVx2_ASAP7_75t_L g17488 ( 
.A(n_17290),
.Y(n_17488)
);

OR2x2_ASAP7_75t_L g17489 ( 
.A(n_17196),
.B(n_2446),
.Y(n_17489)
);

HB1xp67_ASAP7_75t_L g17490 ( 
.A(n_17221),
.Y(n_17490)
);

INVx1_ASAP7_75t_L g17491 ( 
.A(n_17272),
.Y(n_17491)
);

AND2x2_ASAP7_75t_L g17492 ( 
.A(n_17222),
.B(n_2447),
.Y(n_17492)
);

AOI22xp33_ASAP7_75t_L g17493 ( 
.A1(n_17215),
.A2(n_2449),
.B1(n_2447),
.B2(n_2448),
.Y(n_17493)
);

NAND2xp5_ASAP7_75t_L g17494 ( 
.A(n_17273),
.B(n_2448),
.Y(n_17494)
);

INVx1_ASAP7_75t_L g17495 ( 
.A(n_17310),
.Y(n_17495)
);

INVx3_ASAP7_75t_L g17496 ( 
.A(n_17194),
.Y(n_17496)
);

BUFx6f_ASAP7_75t_L g17497 ( 
.A(n_17323),
.Y(n_17497)
);

AND2x2_ASAP7_75t_L g17498 ( 
.A(n_17314),
.B(n_2449),
.Y(n_17498)
);

INVx1_ASAP7_75t_L g17499 ( 
.A(n_17305),
.Y(n_17499)
);

OR2x2_ASAP7_75t_L g17500 ( 
.A(n_17242),
.B(n_2450),
.Y(n_17500)
);

AND2x2_ASAP7_75t_L g17501 ( 
.A(n_17254),
.B(n_2451),
.Y(n_17501)
);

INVx1_ASAP7_75t_L g17502 ( 
.A(n_17294),
.Y(n_17502)
);

NOR2xp33_ASAP7_75t_L g17503 ( 
.A(n_17328),
.B(n_2451),
.Y(n_17503)
);

AND2x2_ASAP7_75t_L g17504 ( 
.A(n_17250),
.B(n_17292),
.Y(n_17504)
);

INVx1_ASAP7_75t_L g17505 ( 
.A(n_17359),
.Y(n_17505)
);

INVx2_ASAP7_75t_L g17506 ( 
.A(n_17290),
.Y(n_17506)
);

NOR2xp67_ASAP7_75t_L g17507 ( 
.A(n_17349),
.B(n_17228),
.Y(n_17507)
);

INVx1_ASAP7_75t_L g17508 ( 
.A(n_17261),
.Y(n_17508)
);

INVx1_ASAP7_75t_SL g17509 ( 
.A(n_17340),
.Y(n_17509)
);

NAND2xp5_ASAP7_75t_L g17510 ( 
.A(n_17260),
.B(n_2452),
.Y(n_17510)
);

OR2x2_ASAP7_75t_L g17511 ( 
.A(n_17234),
.B(n_2452),
.Y(n_17511)
);

NAND2xp5_ASAP7_75t_L g17512 ( 
.A(n_17339),
.B(n_2453),
.Y(n_17512)
);

NAND2xp5_ASAP7_75t_L g17513 ( 
.A(n_17311),
.B(n_2453),
.Y(n_17513)
);

INVx1_ASAP7_75t_L g17514 ( 
.A(n_17285),
.Y(n_17514)
);

INVx1_ASAP7_75t_L g17515 ( 
.A(n_17271),
.Y(n_17515)
);

INVx1_ASAP7_75t_L g17516 ( 
.A(n_17283),
.Y(n_17516)
);

INVx1_ASAP7_75t_L g17517 ( 
.A(n_17370),
.Y(n_17517)
);

NAND2xp5_ASAP7_75t_L g17518 ( 
.A(n_17320),
.B(n_2454),
.Y(n_17518)
);

AND2x2_ASAP7_75t_L g17519 ( 
.A(n_17249),
.B(n_2454),
.Y(n_17519)
);

BUFx3_ASAP7_75t_L g17520 ( 
.A(n_17372),
.Y(n_17520)
);

INVx3_ASAP7_75t_L g17521 ( 
.A(n_17288),
.Y(n_17521)
);

INVx1_ASAP7_75t_L g17522 ( 
.A(n_17268),
.Y(n_17522)
);

INVx1_ASAP7_75t_L g17523 ( 
.A(n_17268),
.Y(n_17523)
);

INVx3_ASAP7_75t_L g17524 ( 
.A(n_17362),
.Y(n_17524)
);

INVx1_ASAP7_75t_L g17525 ( 
.A(n_17341),
.Y(n_17525)
);

INVx2_ASAP7_75t_L g17526 ( 
.A(n_17183),
.Y(n_17526)
);

HB1xp67_ASAP7_75t_L g17527 ( 
.A(n_17275),
.Y(n_17527)
);

AND2x4_ASAP7_75t_L g17528 ( 
.A(n_17241),
.B(n_2455),
.Y(n_17528)
);

AND2x4_ASAP7_75t_SL g17529 ( 
.A(n_17361),
.B(n_2455),
.Y(n_17529)
);

INVx1_ASAP7_75t_L g17530 ( 
.A(n_17348),
.Y(n_17530)
);

INVx1_ASAP7_75t_L g17531 ( 
.A(n_17363),
.Y(n_17531)
);

HB1xp67_ASAP7_75t_L g17532 ( 
.A(n_17318),
.Y(n_17532)
);

INVx1_ASAP7_75t_L g17533 ( 
.A(n_17279),
.Y(n_17533)
);

AND2x2_ASAP7_75t_L g17534 ( 
.A(n_17389),
.B(n_17246),
.Y(n_17534)
);

NAND2xp5_ASAP7_75t_L g17535 ( 
.A(n_17464),
.B(n_17182),
.Y(n_17535)
);

NAND3xp33_ASAP7_75t_L g17536 ( 
.A(n_17378),
.B(n_17203),
.C(n_17255),
.Y(n_17536)
);

AND2x2_ASAP7_75t_L g17537 ( 
.A(n_17384),
.B(n_17227),
.Y(n_17537)
);

OAI221xp5_ASAP7_75t_L g17538 ( 
.A1(n_17426),
.A2(n_17201),
.B1(n_17205),
.B2(n_17186),
.C(n_17356),
.Y(n_17538)
);

AND2x2_ASAP7_75t_L g17539 ( 
.A(n_17401),
.B(n_17309),
.Y(n_17539)
);

NOR2xp33_ASAP7_75t_L g17540 ( 
.A(n_17401),
.B(n_17405),
.Y(n_17540)
);

AND2x2_ASAP7_75t_L g17541 ( 
.A(n_17398),
.B(n_17345),
.Y(n_17541)
);

NAND2xp5_ASAP7_75t_L g17542 ( 
.A(n_17509),
.B(n_17243),
.Y(n_17542)
);

OAI221xp5_ASAP7_75t_L g17543 ( 
.A1(n_17408),
.A2(n_17360),
.B1(n_17239),
.B2(n_17216),
.C(n_17219),
.Y(n_17543)
);

NAND2xp5_ASAP7_75t_L g17544 ( 
.A(n_17477),
.B(n_17430),
.Y(n_17544)
);

NAND2xp5_ASAP7_75t_L g17545 ( 
.A(n_17411),
.B(n_17235),
.Y(n_17545)
);

OAI21xp5_ASAP7_75t_L g17546 ( 
.A1(n_17486),
.A2(n_17277),
.B(n_17336),
.Y(n_17546)
);

NAND3xp33_ASAP7_75t_L g17547 ( 
.A(n_17490),
.B(n_17181),
.C(n_17244),
.Y(n_17547)
);

OAI221xp5_ASAP7_75t_L g17548 ( 
.A1(n_17512),
.A2(n_17291),
.B1(n_17192),
.B2(n_17207),
.C(n_17274),
.Y(n_17548)
);

NOR2xp33_ASAP7_75t_L g17549 ( 
.A(n_17419),
.B(n_17329),
.Y(n_17549)
);

NAND2xp5_ASAP7_75t_SL g17550 ( 
.A(n_17474),
.B(n_17350),
.Y(n_17550)
);

NAND3xp33_ASAP7_75t_L g17551 ( 
.A(n_17433),
.B(n_17293),
.C(n_17327),
.Y(n_17551)
);

AND2x2_ASAP7_75t_L g17552 ( 
.A(n_17421),
.B(n_17353),
.Y(n_17552)
);

INVx1_ASAP7_75t_L g17553 ( 
.A(n_17382),
.Y(n_17553)
);

NAND3xp33_ASAP7_75t_L g17554 ( 
.A(n_17457),
.B(n_17330),
.C(n_17366),
.Y(n_17554)
);

AOI22xp33_ASAP7_75t_L g17555 ( 
.A1(n_17390),
.A2(n_17226),
.B1(n_17223),
.B2(n_17375),
.Y(n_17555)
);

NAND3xp33_ASAP7_75t_L g17556 ( 
.A(n_17446),
.B(n_17300),
.C(n_17365),
.Y(n_17556)
);

NAND3xp33_ASAP7_75t_L g17557 ( 
.A(n_17527),
.B(n_17276),
.C(n_17321),
.Y(n_17557)
);

NAND3xp33_ASAP7_75t_L g17558 ( 
.A(n_17532),
.B(n_17367),
.C(n_17266),
.Y(n_17558)
);

NAND2xp5_ASAP7_75t_SL g17559 ( 
.A(n_17452),
.B(n_17299),
.Y(n_17559)
);

NOR2xp33_ASAP7_75t_SL g17560 ( 
.A(n_17407),
.B(n_17357),
.Y(n_17560)
);

AOI22xp33_ASAP7_75t_L g17561 ( 
.A1(n_17392),
.A2(n_17334),
.B1(n_17369),
.B2(n_17189),
.Y(n_17561)
);

NAND3xp33_ASAP7_75t_L g17562 ( 
.A(n_17510),
.B(n_17189),
.C(n_17371),
.Y(n_17562)
);

AOI221xp5_ASAP7_75t_L g17563 ( 
.A1(n_17429),
.A2(n_17258),
.B1(n_2458),
.B2(n_2456),
.C(n_2457),
.Y(n_17563)
);

OAI22xp5_ASAP7_75t_L g17564 ( 
.A1(n_17522),
.A2(n_17258),
.B1(n_2458),
.B2(n_2456),
.Y(n_17564)
);

NAND2xp5_ASAP7_75t_L g17565 ( 
.A(n_17435),
.B(n_17409),
.Y(n_17565)
);

AND2x4_ASAP7_75t_L g17566 ( 
.A(n_17395),
.B(n_2457),
.Y(n_17566)
);

NOR2xp33_ASAP7_75t_R g17567 ( 
.A(n_17424),
.B(n_2459),
.Y(n_17567)
);

NAND2xp5_ASAP7_75t_L g17568 ( 
.A(n_17417),
.B(n_2459),
.Y(n_17568)
);

AND2x2_ASAP7_75t_L g17569 ( 
.A(n_17388),
.B(n_2460),
.Y(n_17569)
);

NOR3xp33_ASAP7_75t_L g17570 ( 
.A(n_17475),
.B(n_2460),
.C(n_2461),
.Y(n_17570)
);

NAND2xp5_ASAP7_75t_L g17571 ( 
.A(n_17444),
.B(n_2461),
.Y(n_17571)
);

NAND4xp25_ASAP7_75t_L g17572 ( 
.A(n_17463),
.B(n_2464),
.C(n_2462),
.D(n_2463),
.Y(n_17572)
);

NAND2xp5_ASAP7_75t_SL g17573 ( 
.A(n_17497),
.B(n_2462),
.Y(n_17573)
);

NAND2xp5_ASAP7_75t_L g17574 ( 
.A(n_17523),
.B(n_2463),
.Y(n_17574)
);

AOI22xp33_ASAP7_75t_L g17575 ( 
.A1(n_17397),
.A2(n_2466),
.B1(n_2464),
.B2(n_2465),
.Y(n_17575)
);

NAND3xp33_ASAP7_75t_L g17576 ( 
.A(n_17458),
.B(n_17415),
.C(n_17470),
.Y(n_17576)
);

OAI221xp5_ASAP7_75t_SL g17577 ( 
.A1(n_17511),
.A2(n_2467),
.B1(n_2465),
.B2(n_2466),
.C(n_2468),
.Y(n_17577)
);

OAI21xp5_ASAP7_75t_SL g17578 ( 
.A1(n_17420),
.A2(n_2467),
.B(n_2468),
.Y(n_17578)
);

AND2x2_ASAP7_75t_L g17579 ( 
.A(n_17439),
.B(n_2469),
.Y(n_17579)
);

NAND2xp5_ASAP7_75t_L g17580 ( 
.A(n_17393),
.B(n_2469),
.Y(n_17580)
);

AOI22xp33_ASAP7_75t_L g17581 ( 
.A1(n_17396),
.A2(n_17453),
.B1(n_17422),
.B2(n_17440),
.Y(n_17581)
);

OAI211xp5_ASAP7_75t_L g17582 ( 
.A1(n_17478),
.A2(n_2472),
.B(n_2470),
.C(n_2471),
.Y(n_17582)
);

AND2x2_ASAP7_75t_L g17583 ( 
.A(n_17403),
.B(n_2470),
.Y(n_17583)
);

NAND2xp5_ASAP7_75t_L g17584 ( 
.A(n_17481),
.B(n_2471),
.Y(n_17584)
);

NAND2xp5_ASAP7_75t_L g17585 ( 
.A(n_17437),
.B(n_2472),
.Y(n_17585)
);

AND2x2_ASAP7_75t_L g17586 ( 
.A(n_17383),
.B(n_2473),
.Y(n_17586)
);

OAI22xp5_ASAP7_75t_L g17587 ( 
.A1(n_17436),
.A2(n_2475),
.B1(n_2473),
.B2(n_2474),
.Y(n_17587)
);

NAND3xp33_ASAP7_75t_L g17588 ( 
.A(n_17448),
.B(n_2475),
.C(n_2476),
.Y(n_17588)
);

OA21x2_ASAP7_75t_L g17589 ( 
.A1(n_17385),
.A2(n_2476),
.B(n_2477),
.Y(n_17589)
);

AND2x2_ASAP7_75t_L g17590 ( 
.A(n_17428),
.B(n_2477),
.Y(n_17590)
);

NAND4xp25_ASAP7_75t_L g17591 ( 
.A(n_17507),
.B(n_2480),
.C(n_2478),
.D(n_2479),
.Y(n_17591)
);

NAND2xp5_ASAP7_75t_L g17592 ( 
.A(n_17449),
.B(n_2478),
.Y(n_17592)
);

NAND4xp25_ASAP7_75t_L g17593 ( 
.A(n_17380),
.B(n_2481),
.C(n_2479),
.D(n_2480),
.Y(n_17593)
);

NOR2xp33_ASAP7_75t_L g17594 ( 
.A(n_17394),
.B(n_2481),
.Y(n_17594)
);

NAND2xp5_ASAP7_75t_L g17595 ( 
.A(n_17488),
.B(n_2482),
.Y(n_17595)
);

OAI21xp5_ASAP7_75t_L g17596 ( 
.A1(n_17387),
.A2(n_2482),
.B(n_2483),
.Y(n_17596)
);

AND2x2_ASAP7_75t_L g17597 ( 
.A(n_17442),
.B(n_17434),
.Y(n_17597)
);

OAI21xp33_ASAP7_75t_L g17598 ( 
.A1(n_17479),
.A2(n_2483),
.B(n_2484),
.Y(n_17598)
);

NAND2xp5_ASAP7_75t_L g17599 ( 
.A(n_17506),
.B(n_2484),
.Y(n_17599)
);

AOI22xp33_ASAP7_75t_L g17600 ( 
.A1(n_17400),
.A2(n_2487),
.B1(n_2485),
.B2(n_2486),
.Y(n_17600)
);

NAND2xp5_ASAP7_75t_L g17601 ( 
.A(n_17496),
.B(n_2485),
.Y(n_17601)
);

NAND3xp33_ASAP7_75t_L g17602 ( 
.A(n_17381),
.B(n_2487),
.C(n_2488),
.Y(n_17602)
);

NAND2xp5_ASAP7_75t_L g17603 ( 
.A(n_17521),
.B(n_17471),
.Y(n_17603)
);

INVx1_ASAP7_75t_L g17604 ( 
.A(n_17377),
.Y(n_17604)
);

AND2x2_ASAP7_75t_L g17605 ( 
.A(n_17451),
.B(n_17425),
.Y(n_17605)
);

AND2x2_ASAP7_75t_L g17606 ( 
.A(n_17391),
.B(n_2488),
.Y(n_17606)
);

INVx1_ASAP7_75t_L g17607 ( 
.A(n_17379),
.Y(n_17607)
);

NAND2xp5_ASAP7_75t_L g17608 ( 
.A(n_17413),
.B(n_2489),
.Y(n_17608)
);

NAND2xp5_ASAP7_75t_L g17609 ( 
.A(n_17524),
.B(n_2489),
.Y(n_17609)
);

NAND4xp25_ASAP7_75t_L g17610 ( 
.A(n_17412),
.B(n_17455),
.C(n_17410),
.D(n_17416),
.Y(n_17610)
);

AOI22xp33_ASAP7_75t_L g17611 ( 
.A1(n_17404),
.A2(n_2492),
.B1(n_2490),
.B2(n_2491),
.Y(n_17611)
);

NAND3xp33_ASAP7_75t_L g17612 ( 
.A(n_17497),
.B(n_2490),
.C(n_2491),
.Y(n_17612)
);

NAND2xp5_ASAP7_75t_L g17613 ( 
.A(n_17484),
.B(n_2492),
.Y(n_17613)
);

OAI221xp5_ASAP7_75t_L g17614 ( 
.A1(n_17493),
.A2(n_2495),
.B1(n_2493),
.B2(n_2494),
.C(n_2496),
.Y(n_17614)
);

OAI221xp5_ASAP7_75t_L g17615 ( 
.A1(n_17406),
.A2(n_2495),
.B1(n_2493),
.B2(n_2494),
.C(n_2496),
.Y(n_17615)
);

AND2x2_ASAP7_75t_L g17616 ( 
.A(n_17504),
.B(n_2497),
.Y(n_17616)
);

OAI221xp5_ASAP7_75t_SL g17617 ( 
.A1(n_17460),
.A2(n_2499),
.B1(n_2497),
.B2(n_2498),
.C(n_2500),
.Y(n_17617)
);

OAI21xp5_ASAP7_75t_L g17618 ( 
.A1(n_17494),
.A2(n_2498),
.B(n_2499),
.Y(n_17618)
);

AND2x2_ASAP7_75t_L g17619 ( 
.A(n_17432),
.B(n_2500),
.Y(n_17619)
);

NAND2xp5_ASAP7_75t_SL g17620 ( 
.A(n_17459),
.B(n_2501),
.Y(n_17620)
);

NOR2xp33_ASAP7_75t_L g17621 ( 
.A(n_17447),
.B(n_2501),
.Y(n_17621)
);

AND2x2_ASAP7_75t_L g17622 ( 
.A(n_17438),
.B(n_2502),
.Y(n_17622)
);

NAND2xp5_ASAP7_75t_SL g17623 ( 
.A(n_17520),
.B(n_2503),
.Y(n_17623)
);

AND2x2_ASAP7_75t_L g17624 ( 
.A(n_17498),
.B(n_2503),
.Y(n_17624)
);

AOI221x1_ASAP7_75t_SL g17625 ( 
.A1(n_17456),
.A2(n_17414),
.B1(n_17402),
.B2(n_17399),
.C(n_17386),
.Y(n_17625)
);

OAI22xp5_ASAP7_75t_L g17626 ( 
.A1(n_17473),
.A2(n_2506),
.B1(n_2504),
.B2(n_2505),
.Y(n_17626)
);

NAND3xp33_ASAP7_75t_L g17627 ( 
.A(n_17423),
.B(n_2504),
.C(n_2505),
.Y(n_17627)
);

NAND2xp5_ASAP7_75t_L g17628 ( 
.A(n_17501),
.B(n_2506),
.Y(n_17628)
);

AND2x2_ASAP7_75t_L g17629 ( 
.A(n_17517),
.B(n_2508),
.Y(n_17629)
);

NAND2xp5_ASAP7_75t_L g17630 ( 
.A(n_17469),
.B(n_2509),
.Y(n_17630)
);

NAND2xp5_ASAP7_75t_L g17631 ( 
.A(n_17492),
.B(n_2509),
.Y(n_17631)
);

NAND3xp33_ASAP7_75t_L g17632 ( 
.A(n_17427),
.B(n_2510),
.C(n_2511),
.Y(n_17632)
);

NAND2xp5_ASAP7_75t_L g17633 ( 
.A(n_17519),
.B(n_2510),
.Y(n_17633)
);

AND2x2_ASAP7_75t_L g17634 ( 
.A(n_17515),
.B(n_2511),
.Y(n_17634)
);

OAI21xp5_ASAP7_75t_SL g17635 ( 
.A1(n_17476),
.A2(n_2512),
.B(n_2513),
.Y(n_17635)
);

AND2x2_ASAP7_75t_L g17636 ( 
.A(n_17516),
.B(n_2512),
.Y(n_17636)
);

OAI22xp5_ASAP7_75t_L g17637 ( 
.A1(n_17482),
.A2(n_2516),
.B1(n_2513),
.B2(n_2514),
.Y(n_17637)
);

AND2x2_ASAP7_75t_L g17638 ( 
.A(n_17502),
.B(n_2514),
.Y(n_17638)
);

AND2x2_ASAP7_75t_L g17639 ( 
.A(n_17499),
.B(n_2516),
.Y(n_17639)
);

AND2x2_ASAP7_75t_L g17640 ( 
.A(n_17495),
.B(n_2517),
.Y(n_17640)
);

NAND4xp25_ASAP7_75t_L g17641 ( 
.A(n_17418),
.B(n_2519),
.C(n_2517),
.D(n_2518),
.Y(n_17641)
);

NAND2xp5_ASAP7_75t_L g17642 ( 
.A(n_17485),
.B(n_2518),
.Y(n_17642)
);

NAND2xp5_ASAP7_75t_L g17643 ( 
.A(n_17480),
.B(n_2519),
.Y(n_17643)
);

AOI221xp5_ASAP7_75t_L g17644 ( 
.A1(n_17441),
.A2(n_2522),
.B1(n_2520),
.B2(n_2521),
.C(n_2523),
.Y(n_17644)
);

OA21x2_ASAP7_75t_L g17645 ( 
.A1(n_17513),
.A2(n_2521),
.B(n_2522),
.Y(n_17645)
);

NOR3xp33_ASAP7_75t_L g17646 ( 
.A(n_17461),
.B(n_2523),
.C(n_2524),
.Y(n_17646)
);

AND2x2_ASAP7_75t_L g17647 ( 
.A(n_17491),
.B(n_17466),
.Y(n_17647)
);

AND2x2_ASAP7_75t_L g17648 ( 
.A(n_17467),
.B(n_2524),
.Y(n_17648)
);

AND2x2_ASAP7_75t_L g17649 ( 
.A(n_17468),
.B(n_2525),
.Y(n_17649)
);

INVx1_ASAP7_75t_L g17650 ( 
.A(n_17431),
.Y(n_17650)
);

BUFx2_ASAP7_75t_SL g17651 ( 
.A(n_17528),
.Y(n_17651)
);

OAI21xp33_ASAP7_75t_L g17652 ( 
.A1(n_17508),
.A2(n_2525),
.B(n_2526),
.Y(n_17652)
);

OAI221xp5_ASAP7_75t_SL g17653 ( 
.A1(n_17526),
.A2(n_17462),
.B1(n_17445),
.B2(n_17443),
.C(n_17500),
.Y(n_17653)
);

NOR2xp33_ASAP7_75t_L g17654 ( 
.A(n_17447),
.B(n_2526),
.Y(n_17654)
);

AND2x2_ASAP7_75t_L g17655 ( 
.A(n_17450),
.B(n_2527),
.Y(n_17655)
);

NAND2xp5_ASAP7_75t_L g17656 ( 
.A(n_17533),
.B(n_2527),
.Y(n_17656)
);

NAND2xp5_ASAP7_75t_L g17657 ( 
.A(n_17454),
.B(n_2528),
.Y(n_17657)
);

NOR2xp33_ASAP7_75t_L g17658 ( 
.A(n_17483),
.B(n_2528),
.Y(n_17658)
);

NAND2xp5_ASAP7_75t_L g17659 ( 
.A(n_17465),
.B(n_2529),
.Y(n_17659)
);

NAND2xp5_ASAP7_75t_L g17660 ( 
.A(n_17472),
.B(n_2529),
.Y(n_17660)
);

NAND2xp5_ASAP7_75t_L g17661 ( 
.A(n_17503),
.B(n_2530),
.Y(n_17661)
);

NAND2xp5_ASAP7_75t_L g17662 ( 
.A(n_17505),
.B(n_2530),
.Y(n_17662)
);

OAI21xp33_ASAP7_75t_SL g17663 ( 
.A1(n_17525),
.A2(n_2531),
.B(n_2532),
.Y(n_17663)
);

AOI22xp33_ASAP7_75t_L g17664 ( 
.A1(n_17514),
.A2(n_2534),
.B1(n_2531),
.B2(n_2533),
.Y(n_17664)
);

NAND3xp33_ASAP7_75t_L g17665 ( 
.A(n_17487),
.B(n_17531),
.C(n_17530),
.Y(n_17665)
);

AND2x2_ASAP7_75t_L g17666 ( 
.A(n_17529),
.B(n_2535),
.Y(n_17666)
);

AND2x2_ASAP7_75t_L g17667 ( 
.A(n_17534),
.B(n_17489),
.Y(n_17667)
);

OR2x6_ASAP7_75t_L g17668 ( 
.A(n_17651),
.B(n_17518),
.Y(n_17668)
);

INVx2_ASAP7_75t_SL g17669 ( 
.A(n_17566),
.Y(n_17669)
);

A2O1A1Ixp33_ASAP7_75t_L g17670 ( 
.A1(n_17547),
.A2(n_2537),
.B(n_2535),
.C(n_2536),
.Y(n_17670)
);

NAND3xp33_ASAP7_75t_L g17671 ( 
.A(n_17536),
.B(n_2536),
.C(n_2537),
.Y(n_17671)
);

NAND2xp5_ASAP7_75t_L g17672 ( 
.A(n_17605),
.B(n_2538),
.Y(n_17672)
);

NAND2xp5_ASAP7_75t_L g17673 ( 
.A(n_17541),
.B(n_2538),
.Y(n_17673)
);

INVxp67_ASAP7_75t_L g17674 ( 
.A(n_17540),
.Y(n_17674)
);

INVx4_ASAP7_75t_SL g17675 ( 
.A(n_17566),
.Y(n_17675)
);

INVx2_ASAP7_75t_SL g17676 ( 
.A(n_17597),
.Y(n_17676)
);

INVx1_ASAP7_75t_L g17677 ( 
.A(n_17565),
.Y(n_17677)
);

NAND2xp5_ASAP7_75t_L g17678 ( 
.A(n_17552),
.B(n_2539),
.Y(n_17678)
);

INVxp67_ASAP7_75t_SL g17679 ( 
.A(n_17544),
.Y(n_17679)
);

NAND2xp5_ASAP7_75t_L g17680 ( 
.A(n_17560),
.B(n_2539),
.Y(n_17680)
);

OAI21x1_ASAP7_75t_L g17681 ( 
.A1(n_17545),
.A2(n_2540),
.B(n_2541),
.Y(n_17681)
);

AOI21xp5_ASAP7_75t_L g17682 ( 
.A1(n_17538),
.A2(n_2541),
.B(n_2542),
.Y(n_17682)
);

AND2x4_ASAP7_75t_L g17683 ( 
.A(n_17537),
.B(n_2542),
.Y(n_17683)
);

INVx2_ASAP7_75t_L g17684 ( 
.A(n_17622),
.Y(n_17684)
);

OR2x2_ASAP7_75t_L g17685 ( 
.A(n_17591),
.B(n_2543),
.Y(n_17685)
);

INVx1_ASAP7_75t_L g17686 ( 
.A(n_17569),
.Y(n_17686)
);

CKINVDCx6p67_ASAP7_75t_R g17687 ( 
.A(n_17583),
.Y(n_17687)
);

INVx4_ASAP7_75t_L g17688 ( 
.A(n_17666),
.Y(n_17688)
);

INVx2_ASAP7_75t_L g17689 ( 
.A(n_17579),
.Y(n_17689)
);

OA21x2_ASAP7_75t_L g17690 ( 
.A1(n_17535),
.A2(n_17576),
.B(n_17550),
.Y(n_17690)
);

AOI21xp33_ASAP7_75t_L g17691 ( 
.A1(n_17543),
.A2(n_2543),
.B(n_2544),
.Y(n_17691)
);

INVx1_ASAP7_75t_L g17692 ( 
.A(n_17553),
.Y(n_17692)
);

NAND2xp5_ASAP7_75t_L g17693 ( 
.A(n_17581),
.B(n_2544),
.Y(n_17693)
);

NOR2xp33_ASAP7_75t_L g17694 ( 
.A(n_17548),
.B(n_2545),
.Y(n_17694)
);

INVx2_ASAP7_75t_L g17695 ( 
.A(n_17586),
.Y(n_17695)
);

OR2x2_ASAP7_75t_L g17696 ( 
.A(n_17542),
.B(n_2545),
.Y(n_17696)
);

AND2x2_ASAP7_75t_L g17697 ( 
.A(n_17539),
.B(n_2546),
.Y(n_17697)
);

INVx4_ASAP7_75t_L g17698 ( 
.A(n_17606),
.Y(n_17698)
);

OR2x6_ASAP7_75t_L g17699 ( 
.A(n_17619),
.B(n_2547),
.Y(n_17699)
);

INVxp67_ASAP7_75t_L g17700 ( 
.A(n_17621),
.Y(n_17700)
);

INVx2_ASAP7_75t_L g17701 ( 
.A(n_17590),
.Y(n_17701)
);

NAND2xp5_ASAP7_75t_L g17702 ( 
.A(n_17564),
.B(n_2547),
.Y(n_17702)
);

INVx2_ASAP7_75t_L g17703 ( 
.A(n_17616),
.Y(n_17703)
);

INVx2_ASAP7_75t_L g17704 ( 
.A(n_17624),
.Y(n_17704)
);

OR2x2_ASAP7_75t_L g17705 ( 
.A(n_17603),
.B(n_17574),
.Y(n_17705)
);

NAND2xp5_ASAP7_75t_L g17706 ( 
.A(n_17654),
.B(n_2548),
.Y(n_17706)
);

INVx2_ASAP7_75t_L g17707 ( 
.A(n_17647),
.Y(n_17707)
);

CKINVDCx20_ASAP7_75t_R g17708 ( 
.A(n_17567),
.Y(n_17708)
);

INVx1_ASAP7_75t_L g17709 ( 
.A(n_17580),
.Y(n_17709)
);

OR2x6_ASAP7_75t_L g17710 ( 
.A(n_17585),
.B(n_2548),
.Y(n_17710)
);

INVx1_ASAP7_75t_L g17711 ( 
.A(n_17571),
.Y(n_17711)
);

A2O1A1Ixp33_ASAP7_75t_L g17712 ( 
.A1(n_17625),
.A2(n_2551),
.B(n_2549),
.C(n_2550),
.Y(n_17712)
);

INVx2_ASAP7_75t_L g17713 ( 
.A(n_17629),
.Y(n_17713)
);

HB1xp67_ASAP7_75t_L g17714 ( 
.A(n_17589),
.Y(n_17714)
);

NAND2xp5_ASAP7_75t_L g17715 ( 
.A(n_17561),
.B(n_2549),
.Y(n_17715)
);

AND2x2_ASAP7_75t_L g17716 ( 
.A(n_17549),
.B(n_2550),
.Y(n_17716)
);

AND2x6_ASAP7_75t_SL g17717 ( 
.A(n_17594),
.B(n_2551),
.Y(n_17717)
);

NAND2xp5_ASAP7_75t_L g17718 ( 
.A(n_17563),
.B(n_2552),
.Y(n_17718)
);

AND2x2_ASAP7_75t_L g17719 ( 
.A(n_17618),
.B(n_2552),
.Y(n_17719)
);

AND2x2_ASAP7_75t_L g17720 ( 
.A(n_17546),
.B(n_2553),
.Y(n_17720)
);

BUFx2_ASAP7_75t_L g17721 ( 
.A(n_17663),
.Y(n_17721)
);

INVx4_ASAP7_75t_L g17722 ( 
.A(n_17655),
.Y(n_17722)
);

BUFx2_ASAP7_75t_L g17723 ( 
.A(n_17589),
.Y(n_17723)
);

OAI21xp5_ASAP7_75t_L g17724 ( 
.A1(n_17551),
.A2(n_2553),
.B(n_2554),
.Y(n_17724)
);

OAI21xp33_ASAP7_75t_L g17725 ( 
.A1(n_17610),
.A2(n_2555),
.B(n_2556),
.Y(n_17725)
);

BUFx2_ASAP7_75t_L g17726 ( 
.A(n_17645),
.Y(n_17726)
);

INVx2_ASAP7_75t_L g17727 ( 
.A(n_17634),
.Y(n_17727)
);

INVx2_ASAP7_75t_L g17728 ( 
.A(n_17636),
.Y(n_17728)
);

OR2x2_ASAP7_75t_L g17729 ( 
.A(n_17592),
.B(n_2555),
.Y(n_17729)
);

HB1xp67_ASAP7_75t_L g17730 ( 
.A(n_17645),
.Y(n_17730)
);

BUFx2_ASAP7_75t_L g17731 ( 
.A(n_17650),
.Y(n_17731)
);

NAND2xp5_ASAP7_75t_L g17732 ( 
.A(n_17635),
.B(n_2556),
.Y(n_17732)
);

INVx1_ASAP7_75t_L g17733 ( 
.A(n_17568),
.Y(n_17733)
);

BUFx3_ASAP7_75t_L g17734 ( 
.A(n_17604),
.Y(n_17734)
);

INVx2_ASAP7_75t_L g17735 ( 
.A(n_17640),
.Y(n_17735)
);

INVx2_ASAP7_75t_L g17736 ( 
.A(n_17638),
.Y(n_17736)
);

AO211x2_ASAP7_75t_L g17737 ( 
.A1(n_17557),
.A2(n_2559),
.B(n_2557),
.C(n_2558),
.Y(n_17737)
);

INVxp67_ASAP7_75t_L g17738 ( 
.A(n_17620),
.Y(n_17738)
);

INVx2_ASAP7_75t_L g17739 ( 
.A(n_17639),
.Y(n_17739)
);

OR2x6_ASAP7_75t_L g17740 ( 
.A(n_17608),
.B(n_2558),
.Y(n_17740)
);

INVx1_ASAP7_75t_L g17741 ( 
.A(n_17613),
.Y(n_17741)
);

OAI21x1_ASAP7_75t_L g17742 ( 
.A1(n_17660),
.A2(n_2559),
.B(n_2560),
.Y(n_17742)
);

INVx2_ASAP7_75t_L g17743 ( 
.A(n_17648),
.Y(n_17743)
);

INVx1_ASAP7_75t_L g17744 ( 
.A(n_17609),
.Y(n_17744)
);

INVx1_ASAP7_75t_SL g17745 ( 
.A(n_17573),
.Y(n_17745)
);

INVx2_ASAP7_75t_L g17746 ( 
.A(n_17649),
.Y(n_17746)
);

INVx2_ASAP7_75t_L g17747 ( 
.A(n_17607),
.Y(n_17747)
);

AOI211xp5_ASAP7_75t_SL g17748 ( 
.A1(n_17653),
.A2(n_2562),
.B(n_2560),
.C(n_2561),
.Y(n_17748)
);

INVx1_ASAP7_75t_L g17749 ( 
.A(n_17628),
.Y(n_17749)
);

AOI21xp33_ASAP7_75t_L g17750 ( 
.A1(n_17556),
.A2(n_2561),
.B(n_2562),
.Y(n_17750)
);

AOI21xp5_ASAP7_75t_L g17751 ( 
.A1(n_17554),
.A2(n_2563),
.B(n_2564),
.Y(n_17751)
);

INVx1_ASAP7_75t_L g17752 ( 
.A(n_17601),
.Y(n_17752)
);

INVx2_ASAP7_75t_L g17753 ( 
.A(n_17584),
.Y(n_17753)
);

OA21x2_ASAP7_75t_L g17754 ( 
.A1(n_17558),
.A2(n_2563),
.B(n_2564),
.Y(n_17754)
);

INVx1_ASAP7_75t_L g17755 ( 
.A(n_17633),
.Y(n_17755)
);

NOR3xp33_ASAP7_75t_L g17756 ( 
.A(n_17559),
.B(n_2565),
.C(n_2566),
.Y(n_17756)
);

AND2x4_ASAP7_75t_L g17757 ( 
.A(n_17612),
.B(n_2565),
.Y(n_17757)
);

OAI21xp33_ASAP7_75t_L g17758 ( 
.A1(n_17555),
.A2(n_17562),
.B(n_17572),
.Y(n_17758)
);

NAND2xp5_ASAP7_75t_SL g17759 ( 
.A(n_17588),
.B(n_2566),
.Y(n_17759)
);

INVx2_ASAP7_75t_L g17760 ( 
.A(n_17631),
.Y(n_17760)
);

INVx2_ASAP7_75t_L g17761 ( 
.A(n_17642),
.Y(n_17761)
);

OR2x2_ASAP7_75t_L g17762 ( 
.A(n_17630),
.B(n_2567),
.Y(n_17762)
);

INVx1_ASAP7_75t_L g17763 ( 
.A(n_17643),
.Y(n_17763)
);

NOR2xp33_ASAP7_75t_L g17764 ( 
.A(n_17578),
.B(n_2567),
.Y(n_17764)
);

OR2x2_ASAP7_75t_L g17765 ( 
.A(n_17656),
.B(n_2568),
.Y(n_17765)
);

BUFx2_ASAP7_75t_L g17766 ( 
.A(n_17657),
.Y(n_17766)
);

NAND2xp5_ASAP7_75t_L g17767 ( 
.A(n_17658),
.B(n_2568),
.Y(n_17767)
);

HB1xp67_ASAP7_75t_L g17768 ( 
.A(n_17623),
.Y(n_17768)
);

INVx1_ASAP7_75t_L g17769 ( 
.A(n_17595),
.Y(n_17769)
);

INVx1_ASAP7_75t_L g17770 ( 
.A(n_17599),
.Y(n_17770)
);

INVx1_ASAP7_75t_L g17771 ( 
.A(n_17659),
.Y(n_17771)
);

NAND2xp5_ASAP7_75t_L g17772 ( 
.A(n_17570),
.B(n_2569),
.Y(n_17772)
);

INVx1_ASAP7_75t_L g17773 ( 
.A(n_17662),
.Y(n_17773)
);

AO21x2_ASAP7_75t_L g17774 ( 
.A1(n_17582),
.A2(n_2569),
.B(n_2570),
.Y(n_17774)
);

AOI211x1_ASAP7_75t_SL g17775 ( 
.A1(n_17665),
.A2(n_2572),
.B(n_2570),
.C(n_2571),
.Y(n_17775)
);

INVx2_ASAP7_75t_L g17776 ( 
.A(n_17661),
.Y(n_17776)
);

INVx3_ASAP7_75t_L g17777 ( 
.A(n_17577),
.Y(n_17777)
);

INVx4_ASAP7_75t_SL g17778 ( 
.A(n_17587),
.Y(n_17778)
);

OAI211xp5_ASAP7_75t_L g17779 ( 
.A1(n_17644),
.A2(n_2574),
.B(n_2571),
.C(n_2573),
.Y(n_17779)
);

BUFx6f_ASAP7_75t_L g17780 ( 
.A(n_17602),
.Y(n_17780)
);

INVx1_ASAP7_75t_L g17781 ( 
.A(n_17627),
.Y(n_17781)
);

HB1xp67_ASAP7_75t_L g17782 ( 
.A(n_17596),
.Y(n_17782)
);

BUFx2_ASAP7_75t_L g17783 ( 
.A(n_17675),
.Y(n_17783)
);

INVx2_ASAP7_75t_L g17784 ( 
.A(n_17675),
.Y(n_17784)
);

BUFx2_ASAP7_75t_L g17785 ( 
.A(n_17708),
.Y(n_17785)
);

HB1xp67_ASAP7_75t_L g17786 ( 
.A(n_17669),
.Y(n_17786)
);

NAND3xp33_ASAP7_75t_L g17787 ( 
.A(n_17748),
.B(n_17617),
.C(n_17646),
.Y(n_17787)
);

AND2x2_ASAP7_75t_L g17788 ( 
.A(n_17676),
.B(n_17687),
.Y(n_17788)
);

NAND3xp33_ASAP7_75t_L g17789 ( 
.A(n_17712),
.B(n_17632),
.C(n_17615),
.Y(n_17789)
);

NAND3xp33_ASAP7_75t_L g17790 ( 
.A(n_17670),
.B(n_17664),
.C(n_17575),
.Y(n_17790)
);

INVx1_ASAP7_75t_SL g17791 ( 
.A(n_17721),
.Y(n_17791)
);

INVx3_ASAP7_75t_L g17792 ( 
.A(n_17688),
.Y(n_17792)
);

AND2x2_ASAP7_75t_L g17793 ( 
.A(n_17667),
.B(n_17598),
.Y(n_17793)
);

XOR2xp5_ASAP7_75t_L g17794 ( 
.A(n_17768),
.B(n_17593),
.Y(n_17794)
);

AOI22xp33_ASAP7_75t_L g17795 ( 
.A1(n_17690),
.A2(n_17641),
.B1(n_17614),
.B2(n_17652),
.Y(n_17795)
);

INVx1_ASAP7_75t_L g17796 ( 
.A(n_17714),
.Y(n_17796)
);

AND2x2_ASAP7_75t_L g17797 ( 
.A(n_17684),
.B(n_17611),
.Y(n_17797)
);

OR2x2_ASAP7_75t_L g17798 ( 
.A(n_17774),
.B(n_17626),
.Y(n_17798)
);

AND2x2_ASAP7_75t_SL g17799 ( 
.A(n_17731),
.B(n_17600),
.Y(n_17799)
);

NOR2xp33_ASAP7_75t_L g17800 ( 
.A(n_17698),
.B(n_17637),
.Y(n_17800)
);

NAND3xp33_ASAP7_75t_L g17801 ( 
.A(n_17758),
.B(n_2573),
.C(n_2574),
.Y(n_17801)
);

AND2x4_ASAP7_75t_L g17802 ( 
.A(n_17689),
.B(n_2575),
.Y(n_17802)
);

INVx2_ASAP7_75t_L g17803 ( 
.A(n_17723),
.Y(n_17803)
);

NAND2xp5_ASAP7_75t_L g17804 ( 
.A(n_17722),
.B(n_2575),
.Y(n_17804)
);

OR2x2_ASAP7_75t_L g17805 ( 
.A(n_17680),
.B(n_17726),
.Y(n_17805)
);

AOI22xp33_ASAP7_75t_SL g17806 ( 
.A1(n_17730),
.A2(n_2578),
.B1(n_2576),
.B2(n_2577),
.Y(n_17806)
);

AND2x2_ASAP7_75t_L g17807 ( 
.A(n_17668),
.B(n_2576),
.Y(n_17807)
);

NAND3xp33_ASAP7_75t_L g17808 ( 
.A(n_17694),
.B(n_2577),
.C(n_2579),
.Y(n_17808)
);

INVx2_ASAP7_75t_L g17809 ( 
.A(n_17699),
.Y(n_17809)
);

NAND3xp33_ASAP7_75t_L g17810 ( 
.A(n_17682),
.B(n_17671),
.C(n_17715),
.Y(n_17810)
);

INVx1_ASAP7_75t_L g17811 ( 
.A(n_17716),
.Y(n_17811)
);

AO21x2_ASAP7_75t_L g17812 ( 
.A1(n_17750),
.A2(n_2579),
.B(n_2580),
.Y(n_17812)
);

AND2x4_ASAP7_75t_L g17813 ( 
.A(n_17707),
.B(n_2580),
.Y(n_17813)
);

AND2x2_ASAP7_75t_L g17814 ( 
.A(n_17668),
.B(n_2581),
.Y(n_17814)
);

INVx1_ASAP7_75t_L g17815 ( 
.A(n_17678),
.Y(n_17815)
);

NAND4xp25_ASAP7_75t_L g17816 ( 
.A(n_17691),
.B(n_17674),
.C(n_17777),
.D(n_17781),
.Y(n_17816)
);

NAND3xp33_ASAP7_75t_L g17817 ( 
.A(n_17738),
.B(n_2581),
.C(n_2582),
.Y(n_17817)
);

NAND3xp33_ASAP7_75t_L g17818 ( 
.A(n_17754),
.B(n_2582),
.C(n_2583),
.Y(n_17818)
);

OR2x2_ASAP7_75t_L g17819 ( 
.A(n_17701),
.B(n_2584),
.Y(n_17819)
);

NAND4xp75_ASAP7_75t_L g17820 ( 
.A(n_17692),
.B(n_17677),
.C(n_17751),
.D(n_17686),
.Y(n_17820)
);

NAND2xp5_ASAP7_75t_L g17821 ( 
.A(n_17778),
.B(n_2584),
.Y(n_17821)
);

NAND4xp75_ASAP7_75t_L g17822 ( 
.A(n_17709),
.B(n_2587),
.C(n_2585),
.D(n_2586),
.Y(n_17822)
);

AOI22xp33_ASAP7_75t_L g17823 ( 
.A1(n_17737),
.A2(n_2587),
.B1(n_2585),
.B2(n_2586),
.Y(n_17823)
);

AND2x4_ASAP7_75t_L g17824 ( 
.A(n_17695),
.B(n_2588),
.Y(n_17824)
);

NAND3xp33_ASAP7_75t_L g17825 ( 
.A(n_17724),
.B(n_2588),
.C(n_2589),
.Y(n_17825)
);

BUFx3_ASAP7_75t_L g17826 ( 
.A(n_17683),
.Y(n_17826)
);

OAI22xp5_ASAP7_75t_L g17827 ( 
.A1(n_17745),
.A2(n_2592),
.B1(n_2589),
.B2(n_2591),
.Y(n_17827)
);

NAND4xp25_ASAP7_75t_L g17828 ( 
.A(n_17705),
.B(n_2594),
.C(n_2591),
.D(n_2593),
.Y(n_17828)
);

OR2x2_ASAP7_75t_L g17829 ( 
.A(n_17696),
.B(n_2593),
.Y(n_17829)
);

NAND3xp33_ASAP7_75t_L g17830 ( 
.A(n_17780),
.B(n_2594),
.C(n_2595),
.Y(n_17830)
);

NAND3xp33_ASAP7_75t_L g17831 ( 
.A(n_17780),
.B(n_2595),
.C(n_2596),
.Y(n_17831)
);

NAND3xp33_ASAP7_75t_L g17832 ( 
.A(n_17756),
.B(n_2596),
.C(n_2597),
.Y(n_17832)
);

NOR2xp33_ASAP7_75t_L g17833 ( 
.A(n_17700),
.B(n_2597),
.Y(n_17833)
);

NOR3xp33_ASAP7_75t_L g17834 ( 
.A(n_17679),
.B(n_2598),
.C(n_2599),
.Y(n_17834)
);

AND2x2_ASAP7_75t_L g17835 ( 
.A(n_17720),
.B(n_2598),
.Y(n_17835)
);

AO21x2_ASAP7_75t_L g17836 ( 
.A1(n_17673),
.A2(n_2599),
.B(n_2600),
.Y(n_17836)
);

INVx1_ASAP7_75t_L g17837 ( 
.A(n_17697),
.Y(n_17837)
);

OR2x2_ASAP7_75t_L g17838 ( 
.A(n_17703),
.B(n_2600),
.Y(n_17838)
);

OA211x2_ASAP7_75t_L g17839 ( 
.A1(n_17725),
.A2(n_2603),
.B(n_2601),
.C(n_2602),
.Y(n_17839)
);

NOR3xp33_ASAP7_75t_L g17840 ( 
.A(n_17704),
.B(n_2601),
.C(n_2602),
.Y(n_17840)
);

NAND3xp33_ASAP7_75t_L g17841 ( 
.A(n_17782),
.B(n_2603),
.C(n_2604),
.Y(n_17841)
);

NOR3xp33_ASAP7_75t_L g17842 ( 
.A(n_17766),
.B(n_2604),
.C(n_2605),
.Y(n_17842)
);

AOI22xp5_ASAP7_75t_L g17843 ( 
.A1(n_17713),
.A2(n_2608),
.B1(n_2605),
.B2(n_2606),
.Y(n_17843)
);

AND2x2_ASAP7_75t_L g17844 ( 
.A(n_17727),
.B(n_17728),
.Y(n_17844)
);

AOI22xp5_ASAP7_75t_L g17845 ( 
.A1(n_17735),
.A2(n_2609),
.B1(n_2606),
.B2(n_2608),
.Y(n_17845)
);

NAND3xp33_ASAP7_75t_L g17846 ( 
.A(n_17747),
.B(n_2609),
.C(n_2610),
.Y(n_17846)
);

OR2x2_ASAP7_75t_L g17847 ( 
.A(n_17693),
.B(n_2611),
.Y(n_17847)
);

AND2x2_ASAP7_75t_L g17848 ( 
.A(n_17736),
.B(n_2612),
.Y(n_17848)
);

AND2x2_ASAP7_75t_L g17849 ( 
.A(n_17739),
.B(n_2612),
.Y(n_17849)
);

OA21x2_ASAP7_75t_L g17850 ( 
.A1(n_17681),
.A2(n_2613),
.B(n_2614),
.Y(n_17850)
);

AOI22xp5_ASAP7_75t_L g17851 ( 
.A1(n_17743),
.A2(n_2616),
.B1(n_2614),
.B2(n_2615),
.Y(n_17851)
);

AOI22xp33_ASAP7_75t_L g17852 ( 
.A1(n_17746),
.A2(n_2617),
.B1(n_2615),
.B2(n_2616),
.Y(n_17852)
);

OR2x2_ASAP7_75t_SL g17853 ( 
.A(n_17753),
.B(n_2618),
.Y(n_17853)
);

NAND2xp5_ASAP7_75t_SL g17854 ( 
.A(n_17757),
.B(n_2618),
.Y(n_17854)
);

NAND2xp5_ASAP7_75t_SL g17855 ( 
.A(n_17734),
.B(n_2619),
.Y(n_17855)
);

NOR3xp33_ASAP7_75t_L g17856 ( 
.A(n_17733),
.B(n_2619),
.C(n_2620),
.Y(n_17856)
);

INVx3_ASAP7_75t_L g17857 ( 
.A(n_17699),
.Y(n_17857)
);

NAND4xp75_ASAP7_75t_L g17858 ( 
.A(n_17711),
.B(n_2622),
.C(n_2620),
.D(n_2621),
.Y(n_17858)
);

NAND2xp5_ASAP7_75t_SL g17859 ( 
.A(n_17702),
.B(n_2621),
.Y(n_17859)
);

AOI22xp33_ASAP7_75t_SL g17860 ( 
.A1(n_17718),
.A2(n_2624),
.B1(n_2622),
.B2(n_2623),
.Y(n_17860)
);

INVx2_ASAP7_75t_L g17861 ( 
.A(n_17762),
.Y(n_17861)
);

AND2x2_ASAP7_75t_L g17862 ( 
.A(n_17719),
.B(n_2623),
.Y(n_17862)
);

NOR3xp33_ASAP7_75t_L g17863 ( 
.A(n_17741),
.B(n_2624),
.C(n_2625),
.Y(n_17863)
);

CKINVDCx5p33_ASAP7_75t_R g17864 ( 
.A(n_17717),
.Y(n_17864)
);

AND2x2_ASAP7_75t_L g17865 ( 
.A(n_17710),
.B(n_2626),
.Y(n_17865)
);

AO21x2_ASAP7_75t_L g17866 ( 
.A1(n_17672),
.A2(n_2627),
.B(n_2629),
.Y(n_17866)
);

AND2x2_ASAP7_75t_L g17867 ( 
.A(n_17710),
.B(n_2627),
.Y(n_17867)
);

OAI211xp5_ASAP7_75t_L g17868 ( 
.A1(n_17779),
.A2(n_2631),
.B(n_2629),
.C(n_2630),
.Y(n_17868)
);

OA21x2_ASAP7_75t_L g17869 ( 
.A1(n_17742),
.A2(n_2630),
.B(n_2631),
.Y(n_17869)
);

NAND3xp33_ASAP7_75t_L g17870 ( 
.A(n_17759),
.B(n_2632),
.C(n_2634),
.Y(n_17870)
);

NAND2xp5_ASAP7_75t_L g17871 ( 
.A(n_17764),
.B(n_2632),
.Y(n_17871)
);

OR2x2_ASAP7_75t_L g17872 ( 
.A(n_17732),
.B(n_2634),
.Y(n_17872)
);

NAND2xp5_ASAP7_75t_L g17873 ( 
.A(n_17775),
.B(n_2635),
.Y(n_17873)
);

NOR3xp33_ASAP7_75t_L g17874 ( 
.A(n_17744),
.B(n_2635),
.C(n_2636),
.Y(n_17874)
);

AND2x2_ASAP7_75t_L g17875 ( 
.A(n_17760),
.B(n_17761),
.Y(n_17875)
);

AOI22xp33_ASAP7_75t_L g17876 ( 
.A1(n_17776),
.A2(n_17749),
.B1(n_17763),
.B2(n_17755),
.Y(n_17876)
);

NAND4xp75_ASAP7_75t_L g17877 ( 
.A(n_17752),
.B(n_2638),
.C(n_2636),
.D(n_2637),
.Y(n_17877)
);

AOI22xp33_ASAP7_75t_L g17878 ( 
.A1(n_17769),
.A2(n_2639),
.B1(n_2637),
.B2(n_2638),
.Y(n_17878)
);

AOI221xp5_ASAP7_75t_L g17879 ( 
.A1(n_17770),
.A2(n_2641),
.B1(n_2639),
.B2(n_2640),
.C(n_2642),
.Y(n_17879)
);

HB1xp67_ASAP7_75t_L g17880 ( 
.A(n_17740),
.Y(n_17880)
);

AOI21xp5_ASAP7_75t_L g17881 ( 
.A1(n_17772),
.A2(n_2640),
.B(n_2641),
.Y(n_17881)
);

AND2x2_ASAP7_75t_L g17882 ( 
.A(n_17740),
.B(n_2643),
.Y(n_17882)
);

OR2x2_ASAP7_75t_L g17883 ( 
.A(n_17685),
.B(n_2643),
.Y(n_17883)
);

AND2x4_ASAP7_75t_L g17884 ( 
.A(n_17771),
.B(n_2644),
.Y(n_17884)
);

NOR3xp33_ASAP7_75t_L g17885 ( 
.A(n_17773),
.B(n_2644),
.C(n_2645),
.Y(n_17885)
);

NAND2xp5_ASAP7_75t_L g17886 ( 
.A(n_17706),
.B(n_17729),
.Y(n_17886)
);

AND2x2_ASAP7_75t_L g17887 ( 
.A(n_17765),
.B(n_2645),
.Y(n_17887)
);

AND2x2_ASAP7_75t_L g17888 ( 
.A(n_17767),
.B(n_2646),
.Y(n_17888)
);

AND2x2_ASAP7_75t_L g17889 ( 
.A(n_17676),
.B(n_2646),
.Y(n_17889)
);

AOI211xp5_ASAP7_75t_L g17890 ( 
.A1(n_17691),
.A2(n_2649),
.B(n_2647),
.C(n_2648),
.Y(n_17890)
);

NAND3xp33_ASAP7_75t_L g17891 ( 
.A(n_17748),
.B(n_2648),
.C(n_2649),
.Y(n_17891)
);

AND2x2_ASAP7_75t_L g17892 ( 
.A(n_17676),
.B(n_2650),
.Y(n_17892)
);

AOI22xp5_ASAP7_75t_L g17893 ( 
.A1(n_17690),
.A2(n_2652),
.B1(n_2650),
.B2(n_2651),
.Y(n_17893)
);

AND2x2_ASAP7_75t_L g17894 ( 
.A(n_17676),
.B(n_2651),
.Y(n_17894)
);

AND2x2_ASAP7_75t_L g17895 ( 
.A(n_17676),
.B(n_2652),
.Y(n_17895)
);

BUFx3_ASAP7_75t_L g17896 ( 
.A(n_17669),
.Y(n_17896)
);

AND2x4_ASAP7_75t_L g17897 ( 
.A(n_17675),
.B(n_2653),
.Y(n_17897)
);

AND2x2_ASAP7_75t_L g17898 ( 
.A(n_17676),
.B(n_2655),
.Y(n_17898)
);

AOI211x1_ASAP7_75t_L g17899 ( 
.A1(n_17758),
.A2(n_2658),
.B(n_2656),
.C(n_2657),
.Y(n_17899)
);

NOR3xp33_ASAP7_75t_L g17900 ( 
.A(n_17758),
.B(n_2656),
.C(n_2657),
.Y(n_17900)
);

OR2x2_ASAP7_75t_L g17901 ( 
.A(n_17669),
.B(n_2658),
.Y(n_17901)
);

OR2x2_ASAP7_75t_L g17902 ( 
.A(n_17669),
.B(n_2659),
.Y(n_17902)
);

AND2x2_ASAP7_75t_L g17903 ( 
.A(n_17676),
.B(n_2660),
.Y(n_17903)
);

OR2x2_ASAP7_75t_L g17904 ( 
.A(n_17669),
.B(n_2660),
.Y(n_17904)
);

NAND3xp33_ASAP7_75t_L g17905 ( 
.A(n_17748),
.B(n_2661),
.C(n_2662),
.Y(n_17905)
);

INVxp67_ASAP7_75t_L g17906 ( 
.A(n_17714),
.Y(n_17906)
);

NAND4xp75_ASAP7_75t_L g17907 ( 
.A(n_17690),
.B(n_2663),
.C(n_2661),
.D(n_2662),
.Y(n_17907)
);

NAND4xp75_ASAP7_75t_L g17908 ( 
.A(n_17690),
.B(n_2665),
.C(n_2663),
.D(n_2664),
.Y(n_17908)
);

AND2x2_ASAP7_75t_L g17909 ( 
.A(n_17788),
.B(n_17791),
.Y(n_17909)
);

INVx2_ASAP7_75t_L g17910 ( 
.A(n_17783),
.Y(n_17910)
);

NOR2x1p5_ASAP7_75t_L g17911 ( 
.A(n_17907),
.B(n_2664),
.Y(n_17911)
);

NAND2xp5_ASAP7_75t_L g17912 ( 
.A(n_17784),
.B(n_2665),
.Y(n_17912)
);

NAND2xp5_ASAP7_75t_L g17913 ( 
.A(n_17786),
.B(n_2666),
.Y(n_17913)
);

AND2x2_ASAP7_75t_L g17914 ( 
.A(n_17785),
.B(n_17896),
.Y(n_17914)
);

INVx2_ASAP7_75t_L g17915 ( 
.A(n_17897),
.Y(n_17915)
);

AND2x4_ASAP7_75t_L g17916 ( 
.A(n_17792),
.B(n_2666),
.Y(n_17916)
);

INVx1_ASAP7_75t_L g17917 ( 
.A(n_17880),
.Y(n_17917)
);

INVx3_ASAP7_75t_L g17918 ( 
.A(n_17826),
.Y(n_17918)
);

NAND2xp5_ASAP7_75t_L g17919 ( 
.A(n_17864),
.B(n_17857),
.Y(n_17919)
);

AND2x4_ASAP7_75t_SL g17920 ( 
.A(n_17809),
.B(n_2667),
.Y(n_17920)
);

AND2x6_ASAP7_75t_SL g17921 ( 
.A(n_17833),
.B(n_17821),
.Y(n_17921)
);

AND2x2_ASAP7_75t_L g17922 ( 
.A(n_17793),
.B(n_2668),
.Y(n_17922)
);

NAND2xp5_ASAP7_75t_L g17923 ( 
.A(n_17803),
.B(n_17807),
.Y(n_17923)
);

OR2x2_ASAP7_75t_L g17924 ( 
.A(n_17853),
.B(n_2668),
.Y(n_17924)
);

AND2x4_ASAP7_75t_L g17925 ( 
.A(n_17837),
.B(n_2669),
.Y(n_17925)
);

NAND2xp5_ASAP7_75t_L g17926 ( 
.A(n_17814),
.B(n_2669),
.Y(n_17926)
);

AND2x4_ASAP7_75t_L g17927 ( 
.A(n_17811),
.B(n_2670),
.Y(n_17927)
);

AND2x4_ASAP7_75t_L g17928 ( 
.A(n_17844),
.B(n_2670),
.Y(n_17928)
);

AND2x2_ASAP7_75t_L g17929 ( 
.A(n_17799),
.B(n_2671),
.Y(n_17929)
);

INVx1_ASAP7_75t_SL g17930 ( 
.A(n_17901),
.Y(n_17930)
);

NAND2xp5_ASAP7_75t_L g17931 ( 
.A(n_17823),
.B(n_2671),
.Y(n_17931)
);

INVx1_ASAP7_75t_L g17932 ( 
.A(n_17796),
.Y(n_17932)
);

OR2x2_ASAP7_75t_L g17933 ( 
.A(n_17798),
.B(n_2672),
.Y(n_17933)
);

INVx1_ASAP7_75t_L g17934 ( 
.A(n_17902),
.Y(n_17934)
);

NAND2xp5_ASAP7_75t_SL g17935 ( 
.A(n_17893),
.B(n_17891),
.Y(n_17935)
);

INVx1_ASAP7_75t_L g17936 ( 
.A(n_17904),
.Y(n_17936)
);

NAND2x1p5_ASAP7_75t_L g17937 ( 
.A(n_17889),
.B(n_17892),
.Y(n_17937)
);

INVx1_ASAP7_75t_L g17938 ( 
.A(n_17894),
.Y(n_17938)
);

NAND2xp5_ASAP7_75t_L g17939 ( 
.A(n_17895),
.B(n_2672),
.Y(n_17939)
);

INVx1_ASAP7_75t_L g17940 ( 
.A(n_17898),
.Y(n_17940)
);

NOR2xp33_ASAP7_75t_L g17941 ( 
.A(n_17787),
.B(n_2673),
.Y(n_17941)
);

INVx1_ASAP7_75t_L g17942 ( 
.A(n_17903),
.Y(n_17942)
);

NAND2xp5_ASAP7_75t_L g17943 ( 
.A(n_17806),
.B(n_2673),
.Y(n_17943)
);

AND2x2_ASAP7_75t_L g17944 ( 
.A(n_17797),
.B(n_17835),
.Y(n_17944)
);

OR2x2_ASAP7_75t_L g17945 ( 
.A(n_17805),
.B(n_2674),
.Y(n_17945)
);

AND2x4_ASAP7_75t_L g17946 ( 
.A(n_17848),
.B(n_2674),
.Y(n_17946)
);

NAND2x1p5_ASAP7_75t_L g17947 ( 
.A(n_17850),
.B(n_2675),
.Y(n_17947)
);

INVxp67_ASAP7_75t_SL g17948 ( 
.A(n_17906),
.Y(n_17948)
);

AND2x4_ASAP7_75t_L g17949 ( 
.A(n_17849),
.B(n_2675),
.Y(n_17949)
);

INVx3_ASAP7_75t_L g17950 ( 
.A(n_17802),
.Y(n_17950)
);

INVx1_ASAP7_75t_L g17951 ( 
.A(n_17882),
.Y(n_17951)
);

INVx1_ASAP7_75t_L g17952 ( 
.A(n_17865),
.Y(n_17952)
);

NAND2xp5_ASAP7_75t_L g17953 ( 
.A(n_17867),
.B(n_2676),
.Y(n_17953)
);

OR2x2_ASAP7_75t_L g17954 ( 
.A(n_17905),
.B(n_2676),
.Y(n_17954)
);

NAND2xp5_ASAP7_75t_L g17955 ( 
.A(n_17899),
.B(n_2677),
.Y(n_17955)
);

AND2x4_ASAP7_75t_L g17956 ( 
.A(n_17875),
.B(n_2677),
.Y(n_17956)
);

INVx1_ASAP7_75t_L g17957 ( 
.A(n_17850),
.Y(n_17957)
);

INVx1_ASAP7_75t_L g17958 ( 
.A(n_17804),
.Y(n_17958)
);

NAND2x1p5_ASAP7_75t_L g17959 ( 
.A(n_17869),
.B(n_2678),
.Y(n_17959)
);

INVx1_ASAP7_75t_L g17960 ( 
.A(n_17862),
.Y(n_17960)
);

HB1xp67_ASAP7_75t_L g17961 ( 
.A(n_17836),
.Y(n_17961)
);

INVxp67_ASAP7_75t_SL g17962 ( 
.A(n_17818),
.Y(n_17962)
);

INVx1_ASAP7_75t_L g17963 ( 
.A(n_17819),
.Y(n_17963)
);

INVx1_ASAP7_75t_L g17964 ( 
.A(n_17838),
.Y(n_17964)
);

INVx1_ASAP7_75t_L g17965 ( 
.A(n_17813),
.Y(n_17965)
);

AND2x2_ASAP7_75t_L g17966 ( 
.A(n_17800),
.B(n_2679),
.Y(n_17966)
);

AND2x2_ASAP7_75t_L g17967 ( 
.A(n_17861),
.B(n_2679),
.Y(n_17967)
);

INVx2_ASAP7_75t_L g17968 ( 
.A(n_17829),
.Y(n_17968)
);

HB1xp67_ASAP7_75t_L g17969 ( 
.A(n_17866),
.Y(n_17969)
);

INVx1_ASAP7_75t_L g17970 ( 
.A(n_17824),
.Y(n_17970)
);

INVx2_ASAP7_75t_L g17971 ( 
.A(n_17883),
.Y(n_17971)
);

OR2x2_ASAP7_75t_L g17972 ( 
.A(n_17816),
.B(n_2680),
.Y(n_17972)
);

NAND2xp5_ASAP7_75t_L g17973 ( 
.A(n_17795),
.B(n_2680),
.Y(n_17973)
);

NAND2xp5_ASAP7_75t_L g17974 ( 
.A(n_17908),
.B(n_2681),
.Y(n_17974)
);

NAND2xp5_ASAP7_75t_L g17975 ( 
.A(n_17887),
.B(n_2681),
.Y(n_17975)
);

OR2x2_ASAP7_75t_L g17976 ( 
.A(n_17789),
.B(n_2682),
.Y(n_17976)
);

AND2x2_ASAP7_75t_L g17977 ( 
.A(n_17888),
.B(n_2683),
.Y(n_17977)
);

NAND2xp5_ASAP7_75t_L g17978 ( 
.A(n_17840),
.B(n_2683),
.Y(n_17978)
);

OR2x6_ASAP7_75t_L g17979 ( 
.A(n_17820),
.B(n_2684),
.Y(n_17979)
);

NAND2xp5_ASAP7_75t_L g17980 ( 
.A(n_17860),
.B(n_2685),
.Y(n_17980)
);

INVx1_ASAP7_75t_L g17981 ( 
.A(n_17794),
.Y(n_17981)
);

INVx1_ASAP7_75t_L g17982 ( 
.A(n_17822),
.Y(n_17982)
);

INVx1_ASAP7_75t_L g17983 ( 
.A(n_17877),
.Y(n_17983)
);

HB1xp67_ASAP7_75t_L g17984 ( 
.A(n_17858),
.Y(n_17984)
);

INVx1_ASAP7_75t_L g17985 ( 
.A(n_17884),
.Y(n_17985)
);

NAND2xp5_ASAP7_75t_L g17986 ( 
.A(n_17900),
.B(n_2685),
.Y(n_17986)
);

OR2x2_ASAP7_75t_L g17987 ( 
.A(n_17812),
.B(n_17810),
.Y(n_17987)
);

INVx2_ASAP7_75t_L g17988 ( 
.A(n_17872),
.Y(n_17988)
);

INVx1_ASAP7_75t_L g17989 ( 
.A(n_17847),
.Y(n_17989)
);

OR2x2_ASAP7_75t_L g17990 ( 
.A(n_17790),
.B(n_2686),
.Y(n_17990)
);

OAI21xp5_ASAP7_75t_L g17991 ( 
.A1(n_17801),
.A2(n_2686),
.B(n_2687),
.Y(n_17991)
);

AND2x2_ASAP7_75t_L g17992 ( 
.A(n_17815),
.B(n_2687),
.Y(n_17992)
);

OR2x2_ASAP7_75t_L g17993 ( 
.A(n_17825),
.B(n_2688),
.Y(n_17993)
);

INVx1_ASAP7_75t_L g17994 ( 
.A(n_17830),
.Y(n_17994)
);

OR2x2_ASAP7_75t_L g17995 ( 
.A(n_17873),
.B(n_2688),
.Y(n_17995)
);

AND2x2_ASAP7_75t_L g17996 ( 
.A(n_17876),
.B(n_2689),
.Y(n_17996)
);

INVx1_ASAP7_75t_L g17997 ( 
.A(n_17831),
.Y(n_17997)
);

AND2x2_ASAP7_75t_L g17998 ( 
.A(n_17854),
.B(n_2689),
.Y(n_17998)
);

OR2x2_ASAP7_75t_L g17999 ( 
.A(n_17808),
.B(n_2690),
.Y(n_17999)
);

AND2x2_ASAP7_75t_L g18000 ( 
.A(n_17834),
.B(n_2690),
.Y(n_18000)
);

INVx2_ASAP7_75t_SL g18001 ( 
.A(n_17855),
.Y(n_18001)
);

INVx1_ASAP7_75t_L g18002 ( 
.A(n_17886),
.Y(n_18002)
);

INVx1_ASAP7_75t_L g18003 ( 
.A(n_17846),
.Y(n_18003)
);

INVx2_ASAP7_75t_L g18004 ( 
.A(n_17871),
.Y(n_18004)
);

NOR2xp67_ASAP7_75t_L g18005 ( 
.A(n_17841),
.B(n_2691),
.Y(n_18005)
);

OAI21xp33_ASAP7_75t_L g18006 ( 
.A1(n_17868),
.A2(n_2691),
.B(n_2692),
.Y(n_18006)
);

INVxp67_ASAP7_75t_SL g18007 ( 
.A(n_17842),
.Y(n_18007)
);

INVx1_ASAP7_75t_L g18008 ( 
.A(n_17817),
.Y(n_18008)
);

BUFx3_ASAP7_75t_L g18009 ( 
.A(n_17870),
.Y(n_18009)
);

NAND2x1p5_ASAP7_75t_L g18010 ( 
.A(n_17859),
.B(n_2692),
.Y(n_18010)
);

HB1xp67_ASAP7_75t_L g18011 ( 
.A(n_17839),
.Y(n_18011)
);

INVx4_ASAP7_75t_L g18012 ( 
.A(n_17885),
.Y(n_18012)
);

AND2x2_ASAP7_75t_L g18013 ( 
.A(n_17890),
.B(n_2693),
.Y(n_18013)
);

NAND2xp5_ASAP7_75t_L g18014 ( 
.A(n_17881),
.B(n_2693),
.Y(n_18014)
);

BUFx2_ASAP7_75t_L g18015 ( 
.A(n_17828),
.Y(n_18015)
);

INVx1_ASAP7_75t_L g18016 ( 
.A(n_17827),
.Y(n_18016)
);

OR2x2_ASAP7_75t_L g18017 ( 
.A(n_17832),
.B(n_2694),
.Y(n_18017)
);

NAND2xp5_ASAP7_75t_L g18018 ( 
.A(n_17856),
.B(n_2694),
.Y(n_18018)
);

OR2x2_ASAP7_75t_L g18019 ( 
.A(n_17863),
.B(n_2695),
.Y(n_18019)
);

AND2x2_ASAP7_75t_L g18020 ( 
.A(n_17874),
.B(n_17852),
.Y(n_18020)
);

INVx1_ASAP7_75t_L g18021 ( 
.A(n_17843),
.Y(n_18021)
);

NAND4xp25_ASAP7_75t_L g18022 ( 
.A(n_17879),
.B(n_2697),
.C(n_2695),
.D(n_2696),
.Y(n_18022)
);

INVx2_ASAP7_75t_L g18023 ( 
.A(n_17845),
.Y(n_18023)
);

AND2x2_ASAP7_75t_L g18024 ( 
.A(n_17851),
.B(n_2696),
.Y(n_18024)
);

OR2x2_ASAP7_75t_L g18025 ( 
.A(n_17878),
.B(n_2698),
.Y(n_18025)
);

AND2x2_ASAP7_75t_L g18026 ( 
.A(n_17788),
.B(n_2698),
.Y(n_18026)
);

BUFx2_ASAP7_75t_L g18027 ( 
.A(n_17783),
.Y(n_18027)
);

INVx2_ASAP7_75t_L g18028 ( 
.A(n_17783),
.Y(n_18028)
);

NAND2xp5_ASAP7_75t_L g18029 ( 
.A(n_17783),
.B(n_2699),
.Y(n_18029)
);

AOI22xp33_ASAP7_75t_L g18030 ( 
.A1(n_17896),
.A2(n_2701),
.B1(n_2699),
.B2(n_2700),
.Y(n_18030)
);

NAND2xp5_ASAP7_75t_L g18031 ( 
.A(n_17783),
.B(n_2700),
.Y(n_18031)
);

NAND2xp5_ASAP7_75t_L g18032 ( 
.A(n_17783),
.B(n_2701),
.Y(n_18032)
);

NAND2xp5_ASAP7_75t_L g18033 ( 
.A(n_17783),
.B(n_2702),
.Y(n_18033)
);

NAND2xp5_ASAP7_75t_L g18034 ( 
.A(n_17783),
.B(n_2702),
.Y(n_18034)
);

AND2x2_ASAP7_75t_L g18035 ( 
.A(n_17788),
.B(n_2703),
.Y(n_18035)
);

INVx1_ASAP7_75t_L g18036 ( 
.A(n_17783),
.Y(n_18036)
);

AND2x2_ASAP7_75t_L g18037 ( 
.A(n_17788),
.B(n_2703),
.Y(n_18037)
);

AND2x2_ASAP7_75t_L g18038 ( 
.A(n_17788),
.B(n_2704),
.Y(n_18038)
);

AND2x4_ASAP7_75t_L g18039 ( 
.A(n_17896),
.B(n_2705),
.Y(n_18039)
);

AND2x2_ASAP7_75t_L g18040 ( 
.A(n_17788),
.B(n_2705),
.Y(n_18040)
);

INVx1_ASAP7_75t_L g18041 ( 
.A(n_17783),
.Y(n_18041)
);

INVx3_ASAP7_75t_L g18042 ( 
.A(n_17896),
.Y(n_18042)
);

INVx1_ASAP7_75t_SL g18043 ( 
.A(n_17783),
.Y(n_18043)
);

INVxp67_ASAP7_75t_L g18044 ( 
.A(n_17783),
.Y(n_18044)
);

INVx2_ASAP7_75t_SL g18045 ( 
.A(n_17783),
.Y(n_18045)
);

AND2x2_ASAP7_75t_L g18046 ( 
.A(n_17788),
.B(n_2706),
.Y(n_18046)
);

AND2x2_ASAP7_75t_L g18047 ( 
.A(n_17788),
.B(n_2706),
.Y(n_18047)
);

NAND2xp5_ASAP7_75t_L g18048 ( 
.A(n_17783),
.B(n_2707),
.Y(n_18048)
);

NAND2xp5_ASAP7_75t_L g18049 ( 
.A(n_17783),
.B(n_2707),
.Y(n_18049)
);

AND2x2_ASAP7_75t_L g18050 ( 
.A(n_17788),
.B(n_2708),
.Y(n_18050)
);

INVx1_ASAP7_75t_SL g18051 ( 
.A(n_17783),
.Y(n_18051)
);

AND2x2_ASAP7_75t_L g18052 ( 
.A(n_17788),
.B(n_2709),
.Y(n_18052)
);

AND2x2_ASAP7_75t_L g18053 ( 
.A(n_17788),
.B(n_2709),
.Y(n_18053)
);

INVx1_ASAP7_75t_L g18054 ( 
.A(n_17783),
.Y(n_18054)
);

OR2x2_ASAP7_75t_L g18055 ( 
.A(n_17791),
.B(n_2710),
.Y(n_18055)
);

NAND2xp5_ASAP7_75t_L g18056 ( 
.A(n_17783),
.B(n_2710),
.Y(n_18056)
);

INVx2_ASAP7_75t_SL g18057 ( 
.A(n_17783),
.Y(n_18057)
);

INVxp67_ASAP7_75t_SL g18058 ( 
.A(n_17906),
.Y(n_18058)
);

INVx1_ASAP7_75t_L g18059 ( 
.A(n_17783),
.Y(n_18059)
);

INVx4_ASAP7_75t_L g18060 ( 
.A(n_18042),
.Y(n_18060)
);

OR2x2_ASAP7_75t_L g18061 ( 
.A(n_18043),
.B(n_2711),
.Y(n_18061)
);

INVx1_ASAP7_75t_L g18062 ( 
.A(n_17947),
.Y(n_18062)
);

OR2x2_ASAP7_75t_L g18063 ( 
.A(n_18051),
.B(n_2711),
.Y(n_18063)
);

HB1xp67_ASAP7_75t_L g18064 ( 
.A(n_17957),
.Y(n_18064)
);

BUFx2_ASAP7_75t_L g18065 ( 
.A(n_17959),
.Y(n_18065)
);

INVx1_ASAP7_75t_L g18066 ( 
.A(n_18027),
.Y(n_18066)
);

INVx1_ASAP7_75t_L g18067 ( 
.A(n_17961),
.Y(n_18067)
);

AND2x2_ASAP7_75t_L g18068 ( 
.A(n_17914),
.B(n_2712),
.Y(n_18068)
);

OA21x2_ASAP7_75t_L g18069 ( 
.A1(n_17969),
.A2(n_2712),
.B(n_2713),
.Y(n_18069)
);

OA21x2_ASAP7_75t_L g18070 ( 
.A1(n_17974),
.A2(n_2713),
.B(n_2714),
.Y(n_18070)
);

INVx2_ASAP7_75t_SL g18071 ( 
.A(n_17920),
.Y(n_18071)
);

INVx4_ASAP7_75t_L g18072 ( 
.A(n_17918),
.Y(n_18072)
);

INVx1_ASAP7_75t_L g18073 ( 
.A(n_17933),
.Y(n_18073)
);

AND2x2_ASAP7_75t_L g18074 ( 
.A(n_17909),
.B(n_2714),
.Y(n_18074)
);

AO21x2_ASAP7_75t_L g18075 ( 
.A1(n_18029),
.A2(n_2715),
.B(n_2716),
.Y(n_18075)
);

BUFx2_ASAP7_75t_L g18076 ( 
.A(n_17937),
.Y(n_18076)
);

INVx1_ASAP7_75t_L g18077 ( 
.A(n_18036),
.Y(n_18077)
);

INVx3_ASAP7_75t_L g18078 ( 
.A(n_17915),
.Y(n_18078)
);

INVx2_ASAP7_75t_L g18079 ( 
.A(n_18045),
.Y(n_18079)
);

NAND2xp5_ASAP7_75t_L g18080 ( 
.A(n_18057),
.B(n_2715),
.Y(n_18080)
);

NAND2xp5_ASAP7_75t_L g18081 ( 
.A(n_18041),
.B(n_2716),
.Y(n_18081)
);

AND2x2_ASAP7_75t_L g18082 ( 
.A(n_17922),
.B(n_2717),
.Y(n_18082)
);

INVx5_ASAP7_75t_L g18083 ( 
.A(n_17910),
.Y(n_18083)
);

INVx3_ASAP7_75t_L g18084 ( 
.A(n_17950),
.Y(n_18084)
);

INVx1_ASAP7_75t_L g18085 ( 
.A(n_18054),
.Y(n_18085)
);

NOR4xp25_ASAP7_75t_L g18086 ( 
.A(n_18044),
.B(n_2719),
.C(n_2717),
.D(n_2718),
.Y(n_18086)
);

BUFx2_ASAP7_75t_L g18087 ( 
.A(n_17979),
.Y(n_18087)
);

OR2x2_ASAP7_75t_L g18088 ( 
.A(n_18028),
.B(n_2718),
.Y(n_18088)
);

INVxp67_ASAP7_75t_L g18089 ( 
.A(n_18011),
.Y(n_18089)
);

INVx1_ASAP7_75t_L g18090 ( 
.A(n_18059),
.Y(n_18090)
);

BUFx3_ASAP7_75t_L g18091 ( 
.A(n_18039),
.Y(n_18091)
);

BUFx2_ASAP7_75t_L g18092 ( 
.A(n_17979),
.Y(n_18092)
);

HB1xp67_ASAP7_75t_L g18093 ( 
.A(n_17911),
.Y(n_18093)
);

INVx1_ASAP7_75t_L g18094 ( 
.A(n_18026),
.Y(n_18094)
);

AO21x2_ASAP7_75t_L g18095 ( 
.A1(n_18031),
.A2(n_2719),
.B(n_2720),
.Y(n_18095)
);

INVx1_ASAP7_75t_L g18096 ( 
.A(n_18035),
.Y(n_18096)
);

INVx2_ASAP7_75t_SL g18097 ( 
.A(n_17916),
.Y(n_18097)
);

OR2x6_ASAP7_75t_L g18098 ( 
.A(n_17923),
.B(n_2720),
.Y(n_18098)
);

AND2x2_ASAP7_75t_L g18099 ( 
.A(n_17944),
.B(n_2721),
.Y(n_18099)
);

AOI22xp5_ASAP7_75t_L g18100 ( 
.A1(n_17917),
.A2(n_2723),
.B1(n_2721),
.B2(n_2722),
.Y(n_18100)
);

INVx1_ASAP7_75t_L g18101 ( 
.A(n_18037),
.Y(n_18101)
);

INVx1_ASAP7_75t_L g18102 ( 
.A(n_18038),
.Y(n_18102)
);

BUFx3_ASAP7_75t_L g18103 ( 
.A(n_18040),
.Y(n_18103)
);

INVx1_ASAP7_75t_L g18104 ( 
.A(n_18046),
.Y(n_18104)
);

OR2x2_ASAP7_75t_L g18105 ( 
.A(n_17919),
.B(n_2722),
.Y(n_18105)
);

INVx1_ASAP7_75t_L g18106 ( 
.A(n_18047),
.Y(n_18106)
);

INVx1_ASAP7_75t_L g18107 ( 
.A(n_18050),
.Y(n_18107)
);

NAND4xp25_ASAP7_75t_L g18108 ( 
.A(n_17981),
.B(n_2726),
.C(n_2724),
.D(n_2725),
.Y(n_18108)
);

AO21x2_ASAP7_75t_L g18109 ( 
.A1(n_18032),
.A2(n_2727),
.B(n_2728),
.Y(n_18109)
);

INVx2_ASAP7_75t_SL g18110 ( 
.A(n_17928),
.Y(n_18110)
);

AND2x2_ASAP7_75t_L g18111 ( 
.A(n_18052),
.B(n_18053),
.Y(n_18111)
);

OAI31xp33_ASAP7_75t_L g18112 ( 
.A1(n_17929),
.A2(n_2730),
.A3(n_2728),
.B(n_2729),
.Y(n_18112)
);

INVx1_ASAP7_75t_L g18113 ( 
.A(n_17924),
.Y(n_18113)
);

INVx1_ASAP7_75t_L g18114 ( 
.A(n_18033),
.Y(n_18114)
);

INVx3_ASAP7_75t_L g18115 ( 
.A(n_17956),
.Y(n_18115)
);

INVx1_ASAP7_75t_L g18116 ( 
.A(n_18034),
.Y(n_18116)
);

AND2x4_ASAP7_75t_L g18117 ( 
.A(n_17960),
.B(n_2730),
.Y(n_18117)
);

INVx2_ASAP7_75t_SL g18118 ( 
.A(n_17927),
.Y(n_18118)
);

INVx2_ASAP7_75t_L g18119 ( 
.A(n_18055),
.Y(n_18119)
);

INVx2_ASAP7_75t_L g18120 ( 
.A(n_17946),
.Y(n_18120)
);

OAI21xp5_ASAP7_75t_L g18121 ( 
.A1(n_17948),
.A2(n_2731),
.B(n_2732),
.Y(n_18121)
);

INVx1_ASAP7_75t_L g18122 ( 
.A(n_18048),
.Y(n_18122)
);

INVx2_ASAP7_75t_L g18123 ( 
.A(n_17949),
.Y(n_18123)
);

INVx1_ASAP7_75t_SL g18124 ( 
.A(n_17987),
.Y(n_18124)
);

AND2x2_ASAP7_75t_L g18125 ( 
.A(n_17966),
.B(n_17985),
.Y(n_18125)
);

INVx1_ASAP7_75t_L g18126 ( 
.A(n_18049),
.Y(n_18126)
);

INVx1_ASAP7_75t_L g18127 ( 
.A(n_18056),
.Y(n_18127)
);

INVx1_ASAP7_75t_L g18128 ( 
.A(n_17913),
.Y(n_18128)
);

AOI31xp33_ASAP7_75t_L g18129 ( 
.A1(n_18010),
.A2(n_2733),
.A3(n_2731),
.B(n_2732),
.Y(n_18129)
);

AND2x2_ASAP7_75t_L g18130 ( 
.A(n_17965),
.B(n_2733),
.Y(n_18130)
);

INVx2_ASAP7_75t_L g18131 ( 
.A(n_17925),
.Y(n_18131)
);

INVx1_ASAP7_75t_SL g18132 ( 
.A(n_17930),
.Y(n_18132)
);

HB1xp67_ASAP7_75t_L g18133 ( 
.A(n_18005),
.Y(n_18133)
);

BUFx2_ASAP7_75t_L g18134 ( 
.A(n_18058),
.Y(n_18134)
);

OAI21x1_ASAP7_75t_L g18135 ( 
.A1(n_17991),
.A2(n_2734),
.B(n_2735),
.Y(n_18135)
);

OR2x2_ASAP7_75t_L g18136 ( 
.A(n_17955),
.B(n_2735),
.Y(n_18136)
);

AND2x2_ASAP7_75t_L g18137 ( 
.A(n_17970),
.B(n_2736),
.Y(n_18137)
);

INVx1_ASAP7_75t_L g18138 ( 
.A(n_17945),
.Y(n_18138)
);

INVx1_ASAP7_75t_SL g18139 ( 
.A(n_17998),
.Y(n_18139)
);

AND2x2_ASAP7_75t_L g18140 ( 
.A(n_17938),
.B(n_2736),
.Y(n_18140)
);

INVx2_ASAP7_75t_SL g18141 ( 
.A(n_17967),
.Y(n_18141)
);

NAND2xp5_ASAP7_75t_L g18142 ( 
.A(n_17977),
.B(n_2737),
.Y(n_18142)
);

HB1xp67_ASAP7_75t_L g18143 ( 
.A(n_17984),
.Y(n_18143)
);

INVx2_ASAP7_75t_SL g18144 ( 
.A(n_18001),
.Y(n_18144)
);

INVx1_ASAP7_75t_L g18145 ( 
.A(n_17976),
.Y(n_18145)
);

OR2x2_ASAP7_75t_L g18146 ( 
.A(n_17990),
.B(n_17973),
.Y(n_18146)
);

OAI21xp5_ASAP7_75t_L g18147 ( 
.A1(n_17941),
.A2(n_2737),
.B(n_2738),
.Y(n_18147)
);

INVx2_ASAP7_75t_L g18148 ( 
.A(n_17968),
.Y(n_18148)
);

INVx1_ASAP7_75t_L g18149 ( 
.A(n_17926),
.Y(n_18149)
);

OR2x2_ASAP7_75t_L g18150 ( 
.A(n_17995),
.B(n_2738),
.Y(n_18150)
);

INVx1_ASAP7_75t_L g18151 ( 
.A(n_17939),
.Y(n_18151)
);

INVx1_ASAP7_75t_L g18152 ( 
.A(n_17912),
.Y(n_18152)
);

OR2x2_ASAP7_75t_L g18153 ( 
.A(n_17954),
.B(n_2739),
.Y(n_18153)
);

AND2x2_ASAP7_75t_L g18154 ( 
.A(n_17940),
.B(n_2740),
.Y(n_18154)
);

OR2x2_ASAP7_75t_L g18155 ( 
.A(n_17942),
.B(n_2740),
.Y(n_18155)
);

INVx2_ASAP7_75t_L g18156 ( 
.A(n_17992),
.Y(n_18156)
);

HB1xp67_ASAP7_75t_L g18157 ( 
.A(n_17934),
.Y(n_18157)
);

INVx3_ASAP7_75t_L g18158 ( 
.A(n_17971),
.Y(n_18158)
);

AND2x2_ASAP7_75t_L g18159 ( 
.A(n_17951),
.B(n_2741),
.Y(n_18159)
);

BUFx3_ASAP7_75t_L g18160 ( 
.A(n_17952),
.Y(n_18160)
);

INVx1_ASAP7_75t_L g18161 ( 
.A(n_17953),
.Y(n_18161)
);

BUFx3_ASAP7_75t_L g18162 ( 
.A(n_17936),
.Y(n_18162)
);

INVx1_ASAP7_75t_L g18163 ( 
.A(n_17975),
.Y(n_18163)
);

INVx2_ASAP7_75t_L g18164 ( 
.A(n_17999),
.Y(n_18164)
);

INVx1_ASAP7_75t_L g18165 ( 
.A(n_17962),
.Y(n_18165)
);

INVx1_ASAP7_75t_L g18166 ( 
.A(n_17972),
.Y(n_18166)
);

INVx1_ASAP7_75t_L g18167 ( 
.A(n_17996),
.Y(n_18167)
);

INVx1_ASAP7_75t_L g18168 ( 
.A(n_17932),
.Y(n_18168)
);

INVx1_ASAP7_75t_L g18169 ( 
.A(n_17993),
.Y(n_18169)
);

INVx2_ASAP7_75t_SL g18170 ( 
.A(n_17963),
.Y(n_18170)
);

INVx1_ASAP7_75t_L g18171 ( 
.A(n_17943),
.Y(n_18171)
);

INVx1_ASAP7_75t_L g18172 ( 
.A(n_18017),
.Y(n_18172)
);

NOR3xp33_ASAP7_75t_SL g18173 ( 
.A(n_17935),
.B(n_2741),
.C(n_2742),
.Y(n_18173)
);

AOI22xp33_ASAP7_75t_L g18174 ( 
.A1(n_17982),
.A2(n_2744),
.B1(n_2742),
.B2(n_2743),
.Y(n_18174)
);

NAND4xp25_ASAP7_75t_L g18175 ( 
.A(n_18015),
.B(n_18016),
.C(n_17983),
.D(n_18009),
.Y(n_18175)
);

NAND3xp33_ASAP7_75t_L g18176 ( 
.A(n_18006),
.B(n_2743),
.C(n_2744),
.Y(n_18176)
);

AO21x1_ASAP7_75t_L g18177 ( 
.A1(n_18014),
.A2(n_2745),
.B(n_2746),
.Y(n_18177)
);

INVx2_ASAP7_75t_L g18178 ( 
.A(n_17988),
.Y(n_18178)
);

OA21x2_ASAP7_75t_L g18179 ( 
.A1(n_17931),
.A2(n_2745),
.B(n_2746),
.Y(n_18179)
);

NAND2xp5_ASAP7_75t_L g18180 ( 
.A(n_17964),
.B(n_2747),
.Y(n_18180)
);

OA21x2_ASAP7_75t_L g18181 ( 
.A1(n_17980),
.A2(n_2747),
.B(n_2748),
.Y(n_18181)
);

AND2x2_ASAP7_75t_L g18182 ( 
.A(n_18013),
.B(n_2749),
.Y(n_18182)
);

OR2x2_ASAP7_75t_L g18183 ( 
.A(n_18022),
.B(n_2749),
.Y(n_18183)
);

INVx1_ASAP7_75t_L g18184 ( 
.A(n_18019),
.Y(n_18184)
);

INVx2_ASAP7_75t_SL g18185 ( 
.A(n_17994),
.Y(n_18185)
);

INVx1_ASAP7_75t_SL g18186 ( 
.A(n_18000),
.Y(n_18186)
);

OR2x2_ASAP7_75t_L g18187 ( 
.A(n_18025),
.B(n_17986),
.Y(n_18187)
);

INVx1_ASAP7_75t_L g18188 ( 
.A(n_17978),
.Y(n_18188)
);

BUFx2_ASAP7_75t_L g18189 ( 
.A(n_17921),
.Y(n_18189)
);

INVx2_ASAP7_75t_L g18190 ( 
.A(n_18004),
.Y(n_18190)
);

INVx1_ASAP7_75t_L g18191 ( 
.A(n_17997),
.Y(n_18191)
);

AND2x4_ASAP7_75t_SL g18192 ( 
.A(n_17989),
.B(n_2750),
.Y(n_18192)
);

INVx4_ASAP7_75t_L g18193 ( 
.A(n_18012),
.Y(n_18193)
);

OA21x2_ASAP7_75t_L g18194 ( 
.A1(n_18018),
.A2(n_2750),
.B(n_2751),
.Y(n_18194)
);

INVx1_ASAP7_75t_L g18195 ( 
.A(n_18007),
.Y(n_18195)
);

OR2x2_ASAP7_75t_L g18196 ( 
.A(n_18003),
.B(n_2751),
.Y(n_18196)
);

INVx2_ASAP7_75t_L g18197 ( 
.A(n_17958),
.Y(n_18197)
);

INVx1_ASAP7_75t_L g18198 ( 
.A(n_18008),
.Y(n_18198)
);

INVx2_ASAP7_75t_SL g18199 ( 
.A(n_18002),
.Y(n_18199)
);

BUFx2_ASAP7_75t_L g18200 ( 
.A(n_18023),
.Y(n_18200)
);

INVx2_ASAP7_75t_SL g18201 ( 
.A(n_18024),
.Y(n_18201)
);

NAND2xp5_ASAP7_75t_SL g18202 ( 
.A(n_18021),
.B(n_2753),
.Y(n_18202)
);

AND2x2_ASAP7_75t_L g18203 ( 
.A(n_18111),
.B(n_18020),
.Y(n_18203)
);

OR2x2_ASAP7_75t_L g18204 ( 
.A(n_18086),
.B(n_18030),
.Y(n_18204)
);

OR2x2_ASAP7_75t_L g18205 ( 
.A(n_18062),
.B(n_18071),
.Y(n_18205)
);

INVx2_ASAP7_75t_L g18206 ( 
.A(n_18069),
.Y(n_18206)
);

NAND2xp5_ASAP7_75t_L g18207 ( 
.A(n_18083),
.B(n_2753),
.Y(n_18207)
);

BUFx2_ASAP7_75t_L g18208 ( 
.A(n_18098),
.Y(n_18208)
);

INVx1_ASAP7_75t_L g18209 ( 
.A(n_18064),
.Y(n_18209)
);

OR2x2_ASAP7_75t_L g18210 ( 
.A(n_18061),
.B(n_2754),
.Y(n_18210)
);

NOR2xp33_ASAP7_75t_L g18211 ( 
.A(n_18072),
.B(n_2754),
.Y(n_18211)
);

INVx1_ASAP7_75t_L g18212 ( 
.A(n_18074),
.Y(n_18212)
);

INVx1_ASAP7_75t_SL g18213 ( 
.A(n_18076),
.Y(n_18213)
);

XNOR2xp5_ASAP7_75t_L g18214 ( 
.A(n_18143),
.B(n_2755),
.Y(n_18214)
);

NAND2xp5_ASAP7_75t_L g18215 ( 
.A(n_18083),
.B(n_18099),
.Y(n_18215)
);

INVx1_ASAP7_75t_L g18216 ( 
.A(n_18068),
.Y(n_18216)
);

AND2x2_ASAP7_75t_L g18217 ( 
.A(n_18125),
.B(n_2755),
.Y(n_18217)
);

INVx1_ASAP7_75t_SL g18218 ( 
.A(n_18065),
.Y(n_18218)
);

OR2x2_ASAP7_75t_L g18219 ( 
.A(n_18063),
.B(n_2756),
.Y(n_18219)
);

INVx1_ASAP7_75t_L g18220 ( 
.A(n_18134),
.Y(n_18220)
);

INVx1_ASAP7_75t_L g18221 ( 
.A(n_18066),
.Y(n_18221)
);

INVx1_ASAP7_75t_L g18222 ( 
.A(n_18082),
.Y(n_18222)
);

INVx1_ASAP7_75t_L g18223 ( 
.A(n_18103),
.Y(n_18223)
);

INVx1_ASAP7_75t_L g18224 ( 
.A(n_18157),
.Y(n_18224)
);

INVx1_ASAP7_75t_SL g18225 ( 
.A(n_18192),
.Y(n_18225)
);

BUFx2_ASAP7_75t_L g18226 ( 
.A(n_18098),
.Y(n_18226)
);

AND2x2_ASAP7_75t_L g18227 ( 
.A(n_18078),
.B(n_2757),
.Y(n_18227)
);

OR2x2_ASAP7_75t_L g18228 ( 
.A(n_18097),
.B(n_2757),
.Y(n_18228)
);

AND2x4_ASAP7_75t_L g18229 ( 
.A(n_18079),
.B(n_2758),
.Y(n_18229)
);

AND2x2_ASAP7_75t_L g18230 ( 
.A(n_18084),
.B(n_2758),
.Y(n_18230)
);

AND2x2_ASAP7_75t_L g18231 ( 
.A(n_18115),
.B(n_2759),
.Y(n_18231)
);

AND2x2_ASAP7_75t_L g18232 ( 
.A(n_18060),
.B(n_2759),
.Y(n_18232)
);

INVx1_ASAP7_75t_L g18233 ( 
.A(n_18093),
.Y(n_18233)
);

INVx2_ASAP7_75t_L g18234 ( 
.A(n_18091),
.Y(n_18234)
);

INVx1_ASAP7_75t_L g18235 ( 
.A(n_18130),
.Y(n_18235)
);

AND2x2_ASAP7_75t_L g18236 ( 
.A(n_18089),
.B(n_2760),
.Y(n_18236)
);

HB1xp67_ASAP7_75t_L g18237 ( 
.A(n_18075),
.Y(n_18237)
);

AND2x2_ASAP7_75t_L g18238 ( 
.A(n_18189),
.B(n_2760),
.Y(n_18238)
);

INVx1_ASAP7_75t_L g18239 ( 
.A(n_18137),
.Y(n_18239)
);

INVxp67_ASAP7_75t_SL g18240 ( 
.A(n_18177),
.Y(n_18240)
);

AND2x4_ASAP7_75t_L g18241 ( 
.A(n_18118),
.B(n_2761),
.Y(n_18241)
);

AND2x2_ASAP7_75t_L g18242 ( 
.A(n_18094),
.B(n_2761),
.Y(n_18242)
);

INVx2_ASAP7_75t_L g18243 ( 
.A(n_18095),
.Y(n_18243)
);

OR2x2_ASAP7_75t_L g18244 ( 
.A(n_18110),
.B(n_2762),
.Y(n_18244)
);

INVx2_ASAP7_75t_L g18245 ( 
.A(n_18109),
.Y(n_18245)
);

NAND2x1p5_ASAP7_75t_L g18246 ( 
.A(n_18132),
.B(n_18158),
.Y(n_18246)
);

INVx2_ASAP7_75t_L g18247 ( 
.A(n_18160),
.Y(n_18247)
);

AND2x4_ASAP7_75t_SL g18248 ( 
.A(n_18131),
.B(n_2762),
.Y(n_18248)
);

INVx2_ASAP7_75t_L g18249 ( 
.A(n_18162),
.Y(n_18249)
);

INVx1_ASAP7_75t_SL g18250 ( 
.A(n_18087),
.Y(n_18250)
);

AND2x2_ASAP7_75t_L g18251 ( 
.A(n_18096),
.B(n_2763),
.Y(n_18251)
);

INVx2_ASAP7_75t_L g18252 ( 
.A(n_18117),
.Y(n_18252)
);

OR2x2_ASAP7_75t_L g18253 ( 
.A(n_18080),
.B(n_2763),
.Y(n_18253)
);

INVxp33_ASAP7_75t_L g18254 ( 
.A(n_18108),
.Y(n_18254)
);

AOI22xp5_ASAP7_75t_L g18255 ( 
.A1(n_18144),
.A2(n_2766),
.B1(n_2764),
.B2(n_2765),
.Y(n_18255)
);

AND2x2_ASAP7_75t_L g18256 ( 
.A(n_18101),
.B(n_2764),
.Y(n_18256)
);

AND2x2_ASAP7_75t_L g18257 ( 
.A(n_18102),
.B(n_2765),
.Y(n_18257)
);

INVx1_ASAP7_75t_L g18258 ( 
.A(n_18159),
.Y(n_18258)
);

NAND2xp5_ASAP7_75t_L g18259 ( 
.A(n_18104),
.B(n_18106),
.Y(n_18259)
);

INVx2_ASAP7_75t_SL g18260 ( 
.A(n_18088),
.Y(n_18260)
);

OR2x2_ASAP7_75t_L g18261 ( 
.A(n_18107),
.B(n_2766),
.Y(n_18261)
);

NAND2xp5_ASAP7_75t_L g18262 ( 
.A(n_18140),
.B(n_2767),
.Y(n_18262)
);

INVx1_ASAP7_75t_L g18263 ( 
.A(n_18155),
.Y(n_18263)
);

HB1xp67_ASAP7_75t_L g18264 ( 
.A(n_18194),
.Y(n_18264)
);

OR2x2_ASAP7_75t_L g18265 ( 
.A(n_18136),
.B(n_2767),
.Y(n_18265)
);

NAND2xp5_ASAP7_75t_L g18266 ( 
.A(n_18154),
.B(n_2768),
.Y(n_18266)
);

NAND2xp5_ASAP7_75t_L g18267 ( 
.A(n_18077),
.B(n_2768),
.Y(n_18267)
);

NAND2xp5_ASAP7_75t_L g18268 ( 
.A(n_18085),
.B(n_2769),
.Y(n_18268)
);

INVx2_ASAP7_75t_L g18269 ( 
.A(n_18150),
.Y(n_18269)
);

NAND2xp5_ASAP7_75t_L g18270 ( 
.A(n_18090),
.B(n_2769),
.Y(n_18270)
);

INVx2_ASAP7_75t_L g18271 ( 
.A(n_18070),
.Y(n_18271)
);

AND2x2_ASAP7_75t_L g18272 ( 
.A(n_18120),
.B(n_2770),
.Y(n_18272)
);

INVx1_ASAP7_75t_L g18273 ( 
.A(n_18092),
.Y(n_18273)
);

NOR3xp33_ASAP7_75t_L g18274 ( 
.A(n_18175),
.B(n_2770),
.C(n_2771),
.Y(n_18274)
);

INVx1_ASAP7_75t_L g18275 ( 
.A(n_18129),
.Y(n_18275)
);

AND2x2_ASAP7_75t_L g18276 ( 
.A(n_18123),
.B(n_2771),
.Y(n_18276)
);

NAND2xp5_ASAP7_75t_L g18277 ( 
.A(n_18170),
.B(n_2772),
.Y(n_18277)
);

NOR2xp33_ASAP7_75t_L g18278 ( 
.A(n_18124),
.B(n_2773),
.Y(n_18278)
);

NAND2xp5_ASAP7_75t_L g18279 ( 
.A(n_18141),
.B(n_2773),
.Y(n_18279)
);

INVx2_ASAP7_75t_SL g18280 ( 
.A(n_18148),
.Y(n_18280)
);

AND2x2_ASAP7_75t_L g18281 ( 
.A(n_18200),
.B(n_2774),
.Y(n_18281)
);

NAND2xp5_ASAP7_75t_L g18282 ( 
.A(n_18167),
.B(n_2775),
.Y(n_18282)
);

OR2x2_ASAP7_75t_L g18283 ( 
.A(n_18105),
.B(n_2775),
.Y(n_18283)
);

OR2x2_ASAP7_75t_L g18284 ( 
.A(n_18196),
.B(n_18081),
.Y(n_18284)
);

NAND2xp5_ASAP7_75t_L g18285 ( 
.A(n_18182),
.B(n_2776),
.Y(n_18285)
);

NOR2xp33_ASAP7_75t_L g18286 ( 
.A(n_18073),
.B(n_2776),
.Y(n_18286)
);

NAND2xp5_ASAP7_75t_L g18287 ( 
.A(n_18138),
.B(n_2777),
.Y(n_18287)
);

AND2x2_ASAP7_75t_L g18288 ( 
.A(n_18173),
.B(n_18156),
.Y(n_18288)
);

OR2x2_ASAP7_75t_L g18289 ( 
.A(n_18183),
.B(n_2777),
.Y(n_18289)
);

OR2x2_ASAP7_75t_L g18290 ( 
.A(n_18153),
.B(n_2778),
.Y(n_18290)
);

INVx1_ASAP7_75t_L g18291 ( 
.A(n_18142),
.Y(n_18291)
);

INVx1_ASAP7_75t_SL g18292 ( 
.A(n_18181),
.Y(n_18292)
);

INVx1_ASAP7_75t_L g18293 ( 
.A(n_18133),
.Y(n_18293)
);

AND2x2_ASAP7_75t_L g18294 ( 
.A(n_18178),
.B(n_2778),
.Y(n_18294)
);

INVx1_ASAP7_75t_L g18295 ( 
.A(n_18067),
.Y(n_18295)
);

NAND2xp5_ASAP7_75t_L g18296 ( 
.A(n_18174),
.B(n_2779),
.Y(n_18296)
);

NAND2xp5_ASAP7_75t_L g18297 ( 
.A(n_18112),
.B(n_2779),
.Y(n_18297)
);

AND2x2_ASAP7_75t_L g18298 ( 
.A(n_18113),
.B(n_2780),
.Y(n_18298)
);

NAND2x1p5_ASAP7_75t_L g18299 ( 
.A(n_18139),
.B(n_2780),
.Y(n_18299)
);

OR2x2_ASAP7_75t_L g18300 ( 
.A(n_18180),
.B(n_2781),
.Y(n_18300)
);

INVx2_ASAP7_75t_L g18301 ( 
.A(n_18135),
.Y(n_18301)
);

AOI22xp5_ASAP7_75t_L g18302 ( 
.A1(n_18165),
.A2(n_2783),
.B1(n_2781),
.B2(n_2782),
.Y(n_18302)
);

AND2x2_ASAP7_75t_L g18303 ( 
.A(n_18119),
.B(n_2783),
.Y(n_18303)
);

INVx1_ASAP7_75t_L g18304 ( 
.A(n_18179),
.Y(n_18304)
);

NAND2xp5_ASAP7_75t_L g18305 ( 
.A(n_18201),
.B(n_2784),
.Y(n_18305)
);

NAND2xp5_ASAP7_75t_L g18306 ( 
.A(n_18185),
.B(n_2785),
.Y(n_18306)
);

NAND2xp5_ASAP7_75t_L g18307 ( 
.A(n_18100),
.B(n_2785),
.Y(n_18307)
);

OR2x2_ASAP7_75t_L g18308 ( 
.A(n_18146),
.B(n_2786),
.Y(n_18308)
);

OR2x2_ASAP7_75t_L g18309 ( 
.A(n_18168),
.B(n_2786),
.Y(n_18309)
);

AND2x2_ASAP7_75t_L g18310 ( 
.A(n_18195),
.B(n_2787),
.Y(n_18310)
);

INVx1_ASAP7_75t_L g18311 ( 
.A(n_18176),
.Y(n_18311)
);

AND2x2_ASAP7_75t_L g18312 ( 
.A(n_18145),
.B(n_18166),
.Y(n_18312)
);

OAI22xp33_ASAP7_75t_L g18313 ( 
.A1(n_18199),
.A2(n_2789),
.B1(n_2787),
.B2(n_2788),
.Y(n_18313)
);

INVx2_ASAP7_75t_L g18314 ( 
.A(n_18187),
.Y(n_18314)
);

OAI33xp33_ASAP7_75t_L g18315 ( 
.A1(n_18198),
.A2(n_2790),
.A3(n_2792),
.B1(n_2788),
.B2(n_2789),
.B3(n_2791),
.Y(n_18315)
);

NOR2xp33_ASAP7_75t_L g18316 ( 
.A(n_18193),
.B(n_2790),
.Y(n_18316)
);

AND2x2_ASAP7_75t_L g18317 ( 
.A(n_18190),
.B(n_2791),
.Y(n_18317)
);

INVx1_ASAP7_75t_L g18318 ( 
.A(n_18202),
.Y(n_18318)
);

OR2x2_ASAP7_75t_L g18319 ( 
.A(n_18186),
.B(n_2792),
.Y(n_18319)
);

NAND2xp5_ASAP7_75t_L g18320 ( 
.A(n_18191),
.B(n_2793),
.Y(n_18320)
);

NAND2xp5_ASAP7_75t_L g18321 ( 
.A(n_18149),
.B(n_2793),
.Y(n_18321)
);

HB1xp67_ASAP7_75t_L g18322 ( 
.A(n_18121),
.Y(n_18322)
);

AND2x2_ASAP7_75t_L g18323 ( 
.A(n_18164),
.B(n_2794),
.Y(n_18323)
);

NOR2xp33_ASAP7_75t_L g18324 ( 
.A(n_18171),
.B(n_2794),
.Y(n_18324)
);

INVx1_ASAP7_75t_SL g18325 ( 
.A(n_18169),
.Y(n_18325)
);

NOR2xp67_ASAP7_75t_SL g18326 ( 
.A(n_18172),
.B(n_2795),
.Y(n_18326)
);

INVx1_ASAP7_75t_L g18327 ( 
.A(n_18147),
.Y(n_18327)
);

AND2x2_ASAP7_75t_L g18328 ( 
.A(n_18184),
.B(n_2796),
.Y(n_18328)
);

INVx2_ASAP7_75t_L g18329 ( 
.A(n_18161),
.Y(n_18329)
);

AND2x4_ASAP7_75t_L g18330 ( 
.A(n_18197),
.B(n_2796),
.Y(n_18330)
);

NAND2xp5_ASAP7_75t_L g18331 ( 
.A(n_18163),
.B(n_18114),
.Y(n_18331)
);

OR2x2_ASAP7_75t_L g18332 ( 
.A(n_18116),
.B(n_2797),
.Y(n_18332)
);

NAND2xp5_ASAP7_75t_L g18333 ( 
.A(n_18122),
.B(n_2797),
.Y(n_18333)
);

INVx1_ASAP7_75t_L g18334 ( 
.A(n_18126),
.Y(n_18334)
);

INVx2_ASAP7_75t_L g18335 ( 
.A(n_18151),
.Y(n_18335)
);

AND2x2_ASAP7_75t_L g18336 ( 
.A(n_18127),
.B(n_2798),
.Y(n_18336)
);

OR2x2_ASAP7_75t_L g18337 ( 
.A(n_18152),
.B(n_2799),
.Y(n_18337)
);

INVxp67_ASAP7_75t_SL g18338 ( 
.A(n_18128),
.Y(n_18338)
);

OR2x2_ASAP7_75t_L g18339 ( 
.A(n_18299),
.B(n_18246),
.Y(n_18339)
);

OR2x2_ASAP7_75t_L g18340 ( 
.A(n_18228),
.B(n_18188),
.Y(n_18340)
);

INVx1_ASAP7_75t_L g18341 ( 
.A(n_18237),
.Y(n_18341)
);

BUFx3_ASAP7_75t_L g18342 ( 
.A(n_18208),
.Y(n_18342)
);

AND2x2_ASAP7_75t_L g18343 ( 
.A(n_18203),
.B(n_2800),
.Y(n_18343)
);

INVx1_ASAP7_75t_L g18344 ( 
.A(n_18264),
.Y(n_18344)
);

NAND2xp5_ASAP7_75t_L g18345 ( 
.A(n_18241),
.B(n_2800),
.Y(n_18345)
);

AND2x2_ASAP7_75t_L g18346 ( 
.A(n_18217),
.B(n_2801),
.Y(n_18346)
);

INVx1_ASAP7_75t_L g18347 ( 
.A(n_18214),
.Y(n_18347)
);

AND2x2_ASAP7_75t_L g18348 ( 
.A(n_18213),
.B(n_2801),
.Y(n_18348)
);

AND2x2_ASAP7_75t_L g18349 ( 
.A(n_18238),
.B(n_2802),
.Y(n_18349)
);

AND2x4_ASAP7_75t_L g18350 ( 
.A(n_18234),
.B(n_2802),
.Y(n_18350)
);

INVx1_ASAP7_75t_L g18351 ( 
.A(n_18207),
.Y(n_18351)
);

AND2x2_ASAP7_75t_L g18352 ( 
.A(n_18225),
.B(n_2803),
.Y(n_18352)
);

INVx1_ASAP7_75t_L g18353 ( 
.A(n_18281),
.Y(n_18353)
);

NOR3xp33_ASAP7_75t_L g18354 ( 
.A(n_18273),
.B(n_2803),
.C(n_2805),
.Y(n_18354)
);

INVx2_ASAP7_75t_L g18355 ( 
.A(n_18205),
.Y(n_18355)
);

INVx1_ASAP7_75t_L g18356 ( 
.A(n_18231),
.Y(n_18356)
);

O2A1O1Ixp33_ASAP7_75t_L g18357 ( 
.A1(n_18206),
.A2(n_2807),
.B(n_2805),
.C(n_2806),
.Y(n_18357)
);

OR2x2_ASAP7_75t_L g18358 ( 
.A(n_18244),
.B(n_2806),
.Y(n_18358)
);

AND2x2_ASAP7_75t_L g18359 ( 
.A(n_18272),
.B(n_2807),
.Y(n_18359)
);

INVx1_ASAP7_75t_L g18360 ( 
.A(n_18248),
.Y(n_18360)
);

OR2x2_ASAP7_75t_L g18361 ( 
.A(n_18215),
.B(n_2808),
.Y(n_18361)
);

INVx2_ASAP7_75t_L g18362 ( 
.A(n_18232),
.Y(n_18362)
);

INVx2_ASAP7_75t_SL g18363 ( 
.A(n_18227),
.Y(n_18363)
);

AND2x4_ASAP7_75t_L g18364 ( 
.A(n_18216),
.B(n_18276),
.Y(n_18364)
);

INVx1_ASAP7_75t_L g18365 ( 
.A(n_18230),
.Y(n_18365)
);

AND2x2_ASAP7_75t_L g18366 ( 
.A(n_18218),
.B(n_2808),
.Y(n_18366)
);

AND2x2_ASAP7_75t_L g18367 ( 
.A(n_18250),
.B(n_2809),
.Y(n_18367)
);

INVx1_ASAP7_75t_L g18368 ( 
.A(n_18236),
.Y(n_18368)
);

AND2x2_ASAP7_75t_L g18369 ( 
.A(n_18252),
.B(n_2810),
.Y(n_18369)
);

INVx1_ASAP7_75t_L g18370 ( 
.A(n_18226),
.Y(n_18370)
);

INVxp67_ASAP7_75t_L g18371 ( 
.A(n_18326),
.Y(n_18371)
);

INVx2_ASAP7_75t_SL g18372 ( 
.A(n_18229),
.Y(n_18372)
);

INVx2_ASAP7_75t_L g18373 ( 
.A(n_18261),
.Y(n_18373)
);

NAND2xp5_ASAP7_75t_L g18374 ( 
.A(n_18240),
.B(n_2810),
.Y(n_18374)
);

INVx1_ASAP7_75t_L g18375 ( 
.A(n_18242),
.Y(n_18375)
);

INVx1_ASAP7_75t_L g18376 ( 
.A(n_18251),
.Y(n_18376)
);

INVx1_ASAP7_75t_L g18377 ( 
.A(n_18256),
.Y(n_18377)
);

AND2x2_ASAP7_75t_L g18378 ( 
.A(n_18212),
.B(n_2811),
.Y(n_18378)
);

NAND2xp5_ASAP7_75t_L g18379 ( 
.A(n_18257),
.B(n_2811),
.Y(n_18379)
);

NAND2x1p5_ASAP7_75t_L g18380 ( 
.A(n_18224),
.B(n_2812),
.Y(n_18380)
);

INVxp67_ASAP7_75t_L g18381 ( 
.A(n_18211),
.Y(n_18381)
);

INVx1_ASAP7_75t_L g18382 ( 
.A(n_18298),
.Y(n_18382)
);

INVx2_ASAP7_75t_L g18383 ( 
.A(n_18290),
.Y(n_18383)
);

INVx2_ASAP7_75t_L g18384 ( 
.A(n_18210),
.Y(n_18384)
);

INVx1_ASAP7_75t_SL g18385 ( 
.A(n_18292),
.Y(n_18385)
);

NAND2xp5_ASAP7_75t_L g18386 ( 
.A(n_18330),
.B(n_2812),
.Y(n_18386)
);

INVx1_ASAP7_75t_L g18387 ( 
.A(n_18309),
.Y(n_18387)
);

OR2x2_ASAP7_75t_L g18388 ( 
.A(n_18204),
.B(n_2813),
.Y(n_18388)
);

INVx1_ASAP7_75t_L g18389 ( 
.A(n_18310),
.Y(n_18389)
);

AOI22xp5_ASAP7_75t_L g18390 ( 
.A1(n_18233),
.A2(n_2815),
.B1(n_2813),
.B2(n_2814),
.Y(n_18390)
);

NOR2x1_ASAP7_75t_L g18391 ( 
.A(n_18243),
.B(n_2814),
.Y(n_18391)
);

NAND2xp5_ASAP7_75t_SL g18392 ( 
.A(n_18245),
.B(n_2815),
.Y(n_18392)
);

OR2x2_ASAP7_75t_L g18393 ( 
.A(n_18219),
.B(n_2816),
.Y(n_18393)
);

INVx1_ASAP7_75t_L g18394 ( 
.A(n_18294),
.Y(n_18394)
);

INVx1_ASAP7_75t_L g18395 ( 
.A(n_18328),
.Y(n_18395)
);

OR2x2_ASAP7_75t_L g18396 ( 
.A(n_18308),
.B(n_18319),
.Y(n_18396)
);

AND2x2_ASAP7_75t_L g18397 ( 
.A(n_18220),
.B(n_2816),
.Y(n_18397)
);

AOI22xp5_ASAP7_75t_L g18398 ( 
.A1(n_18221),
.A2(n_2819),
.B1(n_2817),
.B2(n_2818),
.Y(n_18398)
);

NAND2xp5_ASAP7_75t_L g18399 ( 
.A(n_18209),
.B(n_2817),
.Y(n_18399)
);

AND2x2_ASAP7_75t_L g18400 ( 
.A(n_18288),
.B(n_2818),
.Y(n_18400)
);

OR2x2_ASAP7_75t_L g18401 ( 
.A(n_18304),
.B(n_2819),
.Y(n_18401)
);

INVx1_ASAP7_75t_L g18402 ( 
.A(n_18332),
.Y(n_18402)
);

OR2x2_ASAP7_75t_L g18403 ( 
.A(n_18277),
.B(n_18265),
.Y(n_18403)
);

AND3x2_ASAP7_75t_L g18404 ( 
.A(n_18271),
.B(n_18274),
.C(n_18278),
.Y(n_18404)
);

AND2x2_ASAP7_75t_L g18405 ( 
.A(n_18249),
.B(n_2820),
.Y(n_18405)
);

AND2x2_ASAP7_75t_L g18406 ( 
.A(n_18247),
.B(n_2820),
.Y(n_18406)
);

OR2x2_ASAP7_75t_L g18407 ( 
.A(n_18306),
.B(n_18283),
.Y(n_18407)
);

AOI31xp33_ASAP7_75t_L g18408 ( 
.A1(n_18275),
.A2(n_2823),
.A3(n_2821),
.B(n_2822),
.Y(n_18408)
);

INVx1_ASAP7_75t_L g18409 ( 
.A(n_18303),
.Y(n_18409)
);

NAND2xp5_ASAP7_75t_L g18410 ( 
.A(n_18317),
.B(n_2821),
.Y(n_18410)
);

INVx2_ASAP7_75t_SL g18411 ( 
.A(n_18323),
.Y(n_18411)
);

AND2x2_ASAP7_75t_L g18412 ( 
.A(n_18222),
.B(n_2822),
.Y(n_18412)
);

NAND2xp5_ASAP7_75t_L g18413 ( 
.A(n_18280),
.B(n_18313),
.Y(n_18413)
);

AND4x1_ASAP7_75t_L g18414 ( 
.A(n_18316),
.B(n_2826),
.C(n_2824),
.D(n_2825),
.Y(n_18414)
);

BUFx2_ASAP7_75t_L g18415 ( 
.A(n_18336),
.Y(n_18415)
);

NAND2xp5_ASAP7_75t_L g18416 ( 
.A(n_18286),
.B(n_2824),
.Y(n_18416)
);

INVx1_ASAP7_75t_L g18417 ( 
.A(n_18337),
.Y(n_18417)
);

AND2x2_ASAP7_75t_L g18418 ( 
.A(n_18223),
.B(n_18312),
.Y(n_18418)
);

NAND2xp5_ASAP7_75t_L g18419 ( 
.A(n_18235),
.B(n_2825),
.Y(n_18419)
);

NAND2xp5_ASAP7_75t_L g18420 ( 
.A(n_18239),
.B(n_2826),
.Y(n_18420)
);

INVx1_ASAP7_75t_L g18421 ( 
.A(n_18285),
.Y(n_18421)
);

INVx2_ASAP7_75t_L g18422 ( 
.A(n_18253),
.Y(n_18422)
);

INVx1_ASAP7_75t_L g18423 ( 
.A(n_18262),
.Y(n_18423)
);

NAND2xp5_ASAP7_75t_L g18424 ( 
.A(n_18258),
.B(n_2827),
.Y(n_18424)
);

NOR2xp33_ASAP7_75t_SL g18425 ( 
.A(n_18315),
.B(n_2827),
.Y(n_18425)
);

AOI22xp33_ASAP7_75t_L g18426 ( 
.A1(n_18293),
.A2(n_18314),
.B1(n_18325),
.B2(n_18311),
.Y(n_18426)
);

INVx1_ASAP7_75t_L g18427 ( 
.A(n_18266),
.Y(n_18427)
);

NOR2x1_ASAP7_75t_L g18428 ( 
.A(n_18305),
.B(n_2828),
.Y(n_18428)
);

INVx1_ASAP7_75t_L g18429 ( 
.A(n_18279),
.Y(n_18429)
);

AND2x2_ASAP7_75t_L g18430 ( 
.A(n_18269),
.B(n_2828),
.Y(n_18430)
);

AND2x2_ASAP7_75t_L g18431 ( 
.A(n_18260),
.B(n_2829),
.Y(n_18431)
);

AND2x2_ASAP7_75t_L g18432 ( 
.A(n_18322),
.B(n_2829),
.Y(n_18432)
);

AND2x2_ASAP7_75t_L g18433 ( 
.A(n_18263),
.B(n_2830),
.Y(n_18433)
);

AOI22xp5_ASAP7_75t_L g18434 ( 
.A1(n_18259),
.A2(n_2832),
.B1(n_2830),
.B2(n_2831),
.Y(n_18434)
);

HB1xp67_ASAP7_75t_L g18435 ( 
.A(n_18301),
.Y(n_18435)
);

NAND2xp5_ASAP7_75t_L g18436 ( 
.A(n_18255),
.B(n_2831),
.Y(n_18436)
);

NOR2xp33_ASAP7_75t_L g18437 ( 
.A(n_18254),
.B(n_2832),
.Y(n_18437)
);

NAND2xp5_ASAP7_75t_L g18438 ( 
.A(n_18324),
.B(n_2833),
.Y(n_18438)
);

OAI21xp5_ASAP7_75t_SL g18439 ( 
.A1(n_18297),
.A2(n_2833),
.B(n_2834),
.Y(n_18439)
);

OR2x2_ASAP7_75t_L g18440 ( 
.A(n_18289),
.B(n_2834),
.Y(n_18440)
);

NAND2xp5_ASAP7_75t_L g18441 ( 
.A(n_18295),
.B(n_2835),
.Y(n_18441)
);

INVx1_ASAP7_75t_L g18442 ( 
.A(n_18267),
.Y(n_18442)
);

HB1xp67_ASAP7_75t_L g18443 ( 
.A(n_18287),
.Y(n_18443)
);

INVx1_ASAP7_75t_SL g18444 ( 
.A(n_18300),
.Y(n_18444)
);

OR2x2_ASAP7_75t_L g18445 ( 
.A(n_18282),
.B(n_2835),
.Y(n_18445)
);

NAND2xp5_ASAP7_75t_L g18446 ( 
.A(n_18302),
.B(n_2836),
.Y(n_18446)
);

INVx1_ASAP7_75t_SL g18447 ( 
.A(n_18268),
.Y(n_18447)
);

OR2x2_ASAP7_75t_L g18448 ( 
.A(n_18270),
.B(n_2836),
.Y(n_18448)
);

INVx1_ASAP7_75t_L g18449 ( 
.A(n_18320),
.Y(n_18449)
);

INVx1_ASAP7_75t_L g18450 ( 
.A(n_18296),
.Y(n_18450)
);

INVx2_ASAP7_75t_L g18451 ( 
.A(n_18284),
.Y(n_18451)
);

OR2x2_ASAP7_75t_L g18452 ( 
.A(n_18307),
.B(n_2837),
.Y(n_18452)
);

INVx2_ASAP7_75t_L g18453 ( 
.A(n_18291),
.Y(n_18453)
);

NOR2xp33_ASAP7_75t_L g18454 ( 
.A(n_18318),
.B(n_2837),
.Y(n_18454)
);

OR2x2_ASAP7_75t_L g18455 ( 
.A(n_18333),
.B(n_2838),
.Y(n_18455)
);

AND2x2_ASAP7_75t_L g18456 ( 
.A(n_18329),
.B(n_2838),
.Y(n_18456)
);

OAI21xp33_ASAP7_75t_L g18457 ( 
.A1(n_18327),
.A2(n_18338),
.B(n_18331),
.Y(n_18457)
);

NOR2xp33_ASAP7_75t_L g18458 ( 
.A(n_18321),
.B(n_2839),
.Y(n_18458)
);

NAND2xp5_ASAP7_75t_L g18459 ( 
.A(n_18335),
.B(n_2839),
.Y(n_18459)
);

AND2x4_ASAP7_75t_L g18460 ( 
.A(n_18334),
.B(n_2840),
.Y(n_18460)
);

INVx1_ASAP7_75t_SL g18461 ( 
.A(n_18248),
.Y(n_18461)
);

AOI211xp5_ASAP7_75t_L g18462 ( 
.A1(n_18213),
.A2(n_2843),
.B(n_2841),
.C(n_2842),
.Y(n_18462)
);

OR2x2_ASAP7_75t_L g18463 ( 
.A(n_18299),
.B(n_2841),
.Y(n_18463)
);

AND2x2_ASAP7_75t_L g18464 ( 
.A(n_18203),
.B(n_2842),
.Y(n_18464)
);

AND2x2_ASAP7_75t_L g18465 ( 
.A(n_18352),
.B(n_2843),
.Y(n_18465)
);

AOI22xp5_ASAP7_75t_L g18466 ( 
.A1(n_18355),
.A2(n_2846),
.B1(n_2844),
.B2(n_2845),
.Y(n_18466)
);

CKINVDCx20_ASAP7_75t_R g18467 ( 
.A(n_18342),
.Y(n_18467)
);

INVx2_ASAP7_75t_SL g18468 ( 
.A(n_18339),
.Y(n_18468)
);

AND2x2_ASAP7_75t_L g18469 ( 
.A(n_18367),
.B(n_2845),
.Y(n_18469)
);

AND2x2_ASAP7_75t_L g18470 ( 
.A(n_18348),
.B(n_2847),
.Y(n_18470)
);

INVx3_ASAP7_75t_L g18471 ( 
.A(n_18350),
.Y(n_18471)
);

INVx1_ASAP7_75t_L g18472 ( 
.A(n_18343),
.Y(n_18472)
);

INVx1_ASAP7_75t_L g18473 ( 
.A(n_18464),
.Y(n_18473)
);

INVx2_ASAP7_75t_L g18474 ( 
.A(n_18463),
.Y(n_18474)
);

CKINVDCx16_ASAP7_75t_R g18475 ( 
.A(n_18418),
.Y(n_18475)
);

INVxp67_ASAP7_75t_L g18476 ( 
.A(n_18425),
.Y(n_18476)
);

AND2x2_ASAP7_75t_L g18477 ( 
.A(n_18366),
.B(n_2848),
.Y(n_18477)
);

INVx1_ASAP7_75t_L g18478 ( 
.A(n_18349),
.Y(n_18478)
);

HB1xp67_ASAP7_75t_L g18479 ( 
.A(n_18391),
.Y(n_18479)
);

AOI22xp33_ASAP7_75t_L g18480 ( 
.A1(n_18370),
.A2(n_2851),
.B1(n_2849),
.B2(n_2850),
.Y(n_18480)
);

NOR2x1_ASAP7_75t_R g18481 ( 
.A(n_18415),
.B(n_2851),
.Y(n_18481)
);

AND2x2_ASAP7_75t_L g18482 ( 
.A(n_18400),
.B(n_2852),
.Y(n_18482)
);

INVx1_ASAP7_75t_SL g18483 ( 
.A(n_18346),
.Y(n_18483)
);

INVx1_ASAP7_75t_L g18484 ( 
.A(n_18401),
.Y(n_18484)
);

INVx1_ASAP7_75t_L g18485 ( 
.A(n_18378),
.Y(n_18485)
);

NAND2xp5_ASAP7_75t_L g18486 ( 
.A(n_18412),
.B(n_2852),
.Y(n_18486)
);

NAND2xp5_ASAP7_75t_L g18487 ( 
.A(n_18397),
.B(n_2853),
.Y(n_18487)
);

INVx1_ASAP7_75t_SL g18488 ( 
.A(n_18461),
.Y(n_18488)
);

INVx1_ASAP7_75t_L g18489 ( 
.A(n_18380),
.Y(n_18489)
);

INVx1_ASAP7_75t_L g18490 ( 
.A(n_18369),
.Y(n_18490)
);

INVx1_ASAP7_75t_L g18491 ( 
.A(n_18433),
.Y(n_18491)
);

AOI22xp33_ASAP7_75t_L g18492 ( 
.A1(n_18385),
.A2(n_2856),
.B1(n_2854),
.B2(n_2855),
.Y(n_18492)
);

OAI21xp33_ASAP7_75t_SL g18493 ( 
.A1(n_18392),
.A2(n_2855),
.B(n_2856),
.Y(n_18493)
);

OR2x2_ASAP7_75t_L g18494 ( 
.A(n_18388),
.B(n_2857),
.Y(n_18494)
);

INVx1_ASAP7_75t_SL g18495 ( 
.A(n_18358),
.Y(n_18495)
);

AND2x2_ASAP7_75t_L g18496 ( 
.A(n_18362),
.B(n_2857),
.Y(n_18496)
);

OAI22xp5_ASAP7_75t_L g18497 ( 
.A1(n_18426),
.A2(n_2860),
.B1(n_2858),
.B2(n_2859),
.Y(n_18497)
);

AND2x4_ASAP7_75t_L g18498 ( 
.A(n_18364),
.B(n_18360),
.Y(n_18498)
);

AND2x2_ASAP7_75t_L g18499 ( 
.A(n_18359),
.B(n_18405),
.Y(n_18499)
);

AND2x2_ASAP7_75t_L g18500 ( 
.A(n_18406),
.B(n_2859),
.Y(n_18500)
);

AOI21xp5_ASAP7_75t_L g18501 ( 
.A1(n_18344),
.A2(n_2860),
.B(n_2861),
.Y(n_18501)
);

NOR2x1_ASAP7_75t_R g18502 ( 
.A(n_18413),
.B(n_2861),
.Y(n_18502)
);

INVx1_ASAP7_75t_SL g18503 ( 
.A(n_18393),
.Y(n_18503)
);

CKINVDCx16_ASAP7_75t_R g18504 ( 
.A(n_18396),
.Y(n_18504)
);

OAI221xp5_ASAP7_75t_L g18505 ( 
.A1(n_18457),
.A2(n_2864),
.B1(n_2862),
.B2(n_2863),
.C(n_2865),
.Y(n_18505)
);

NAND2xp5_ASAP7_75t_L g18506 ( 
.A(n_18430),
.B(n_2862),
.Y(n_18506)
);

AND2x2_ASAP7_75t_L g18507 ( 
.A(n_18431),
.B(n_2863),
.Y(n_18507)
);

BUFx3_ASAP7_75t_L g18508 ( 
.A(n_18353),
.Y(n_18508)
);

INVx1_ASAP7_75t_SL g18509 ( 
.A(n_18432),
.Y(n_18509)
);

INVx1_ASAP7_75t_L g18510 ( 
.A(n_18460),
.Y(n_18510)
);

BUFx3_ASAP7_75t_L g18511 ( 
.A(n_18356),
.Y(n_18511)
);

HB1xp67_ASAP7_75t_L g18512 ( 
.A(n_18414),
.Y(n_18512)
);

NAND2xp5_ASAP7_75t_L g18513 ( 
.A(n_18408),
.B(n_2865),
.Y(n_18513)
);

AND2x2_ASAP7_75t_L g18514 ( 
.A(n_18371),
.B(n_2866),
.Y(n_18514)
);

NOR2x1p5_ASAP7_75t_L g18515 ( 
.A(n_18379),
.B(n_2866),
.Y(n_18515)
);

AND2x2_ASAP7_75t_L g18516 ( 
.A(n_18372),
.B(n_2867),
.Y(n_18516)
);

INVx1_ASAP7_75t_L g18517 ( 
.A(n_18460),
.Y(n_18517)
);

CKINVDCx16_ASAP7_75t_R g18518 ( 
.A(n_18428),
.Y(n_18518)
);

INVx2_ASAP7_75t_L g18519 ( 
.A(n_18440),
.Y(n_18519)
);

AND2x2_ASAP7_75t_L g18520 ( 
.A(n_18363),
.B(n_2867),
.Y(n_18520)
);

INVx2_ASAP7_75t_L g18521 ( 
.A(n_18361),
.Y(n_18521)
);

INVx1_ASAP7_75t_L g18522 ( 
.A(n_18374),
.Y(n_18522)
);

INVx2_ASAP7_75t_L g18523 ( 
.A(n_18456),
.Y(n_18523)
);

INVx1_ASAP7_75t_SL g18524 ( 
.A(n_18345),
.Y(n_18524)
);

INVx1_ASAP7_75t_L g18525 ( 
.A(n_18435),
.Y(n_18525)
);

NAND2xp5_ASAP7_75t_L g18526 ( 
.A(n_18404),
.B(n_2868),
.Y(n_18526)
);

AND2x4_ASAP7_75t_L g18527 ( 
.A(n_18365),
.B(n_2868),
.Y(n_18527)
);

INVx2_ASAP7_75t_L g18528 ( 
.A(n_18445),
.Y(n_18528)
);

OAI21x1_ASAP7_75t_L g18529 ( 
.A1(n_18357),
.A2(n_18341),
.B(n_18386),
.Y(n_18529)
);

NAND2xp5_ASAP7_75t_L g18530 ( 
.A(n_18462),
.B(n_2869),
.Y(n_18530)
);

AND2x2_ASAP7_75t_L g18531 ( 
.A(n_18383),
.B(n_2869),
.Y(n_18531)
);

NAND3x1_ASAP7_75t_L g18532 ( 
.A(n_18441),
.B(n_2870),
.C(n_2871),
.Y(n_18532)
);

AND2x2_ASAP7_75t_L g18533 ( 
.A(n_18375),
.B(n_2870),
.Y(n_18533)
);

NAND2xp5_ASAP7_75t_L g18534 ( 
.A(n_18354),
.B(n_2871),
.Y(n_18534)
);

OR2x2_ASAP7_75t_L g18535 ( 
.A(n_18399),
.B(n_2872),
.Y(n_18535)
);

NOR2x1_ASAP7_75t_L g18536 ( 
.A(n_18439),
.B(n_2872),
.Y(n_18536)
);

INVx1_ASAP7_75t_L g18537 ( 
.A(n_18410),
.Y(n_18537)
);

INVx1_ASAP7_75t_L g18538 ( 
.A(n_18419),
.Y(n_18538)
);

INVx1_ASAP7_75t_SL g18539 ( 
.A(n_18340),
.Y(n_18539)
);

INVx1_ASAP7_75t_L g18540 ( 
.A(n_18420),
.Y(n_18540)
);

INVx1_ASAP7_75t_L g18541 ( 
.A(n_18424),
.Y(n_18541)
);

INVx1_ASAP7_75t_L g18542 ( 
.A(n_18459),
.Y(n_18542)
);

OR2x2_ASAP7_75t_L g18543 ( 
.A(n_18448),
.B(n_2873),
.Y(n_18543)
);

NAND3xp33_ASAP7_75t_L g18544 ( 
.A(n_18437),
.B(n_2873),
.C(n_2874),
.Y(n_18544)
);

INVxp67_ASAP7_75t_L g18545 ( 
.A(n_18454),
.Y(n_18545)
);

AND2x2_ASAP7_75t_L g18546 ( 
.A(n_18376),
.B(n_2874),
.Y(n_18546)
);

INVx2_ASAP7_75t_SL g18547 ( 
.A(n_18384),
.Y(n_18547)
);

INVx2_ASAP7_75t_SL g18548 ( 
.A(n_18373),
.Y(n_18548)
);

INVx2_ASAP7_75t_L g18549 ( 
.A(n_18455),
.Y(n_18549)
);

INVx2_ASAP7_75t_SL g18550 ( 
.A(n_18411),
.Y(n_18550)
);

INVx1_ASAP7_75t_L g18551 ( 
.A(n_18416),
.Y(n_18551)
);

INVx1_ASAP7_75t_L g18552 ( 
.A(n_18438),
.Y(n_18552)
);

NOR2x1_ASAP7_75t_L g18553 ( 
.A(n_18387),
.B(n_2875),
.Y(n_18553)
);

NOR2xp67_ASAP7_75t_L g18554 ( 
.A(n_18377),
.B(n_2875),
.Y(n_18554)
);

XNOR2xp5_ASAP7_75t_L g18555 ( 
.A(n_18347),
.B(n_2876),
.Y(n_18555)
);

NAND3xp33_ASAP7_75t_L g18556 ( 
.A(n_18458),
.B(n_2877),
.C(n_2878),
.Y(n_18556)
);

INVx1_ASAP7_75t_L g18557 ( 
.A(n_18436),
.Y(n_18557)
);

INVx1_ASAP7_75t_L g18558 ( 
.A(n_18452),
.Y(n_18558)
);

INVx1_ASAP7_75t_L g18559 ( 
.A(n_18382),
.Y(n_18559)
);

NAND2xp5_ASAP7_75t_L g18560 ( 
.A(n_18395),
.B(n_2877),
.Y(n_18560)
);

NAND3xp33_ASAP7_75t_L g18561 ( 
.A(n_18451),
.B(n_2878),
.C(n_2879),
.Y(n_18561)
);

NAND2xp33_ASAP7_75t_SL g18562 ( 
.A(n_18402),
.B(n_2879),
.Y(n_18562)
);

AND2x4_ASAP7_75t_L g18563 ( 
.A(n_18389),
.B(n_2880),
.Y(n_18563)
);

AND2x2_ASAP7_75t_L g18564 ( 
.A(n_18368),
.B(n_2880),
.Y(n_18564)
);

AND2x4_ASAP7_75t_L g18565 ( 
.A(n_18409),
.B(n_18394),
.Y(n_18565)
);

NAND2xp5_ASAP7_75t_L g18566 ( 
.A(n_18417),
.B(n_2881),
.Y(n_18566)
);

INVx2_ASAP7_75t_L g18567 ( 
.A(n_18403),
.Y(n_18567)
);

AND2x2_ASAP7_75t_L g18568 ( 
.A(n_18453),
.B(n_2881),
.Y(n_18568)
);

INVx1_ASAP7_75t_L g18569 ( 
.A(n_18446),
.Y(n_18569)
);

INVx2_ASAP7_75t_L g18570 ( 
.A(n_18407),
.Y(n_18570)
);

INVx1_ASAP7_75t_L g18571 ( 
.A(n_18351),
.Y(n_18571)
);

OR2x2_ASAP7_75t_L g18572 ( 
.A(n_18444),
.B(n_2882),
.Y(n_18572)
);

BUFx2_ASAP7_75t_L g18573 ( 
.A(n_18422),
.Y(n_18573)
);

INVx1_ASAP7_75t_L g18574 ( 
.A(n_18443),
.Y(n_18574)
);

NAND2xp5_ASAP7_75t_L g18575 ( 
.A(n_18434),
.B(n_2882),
.Y(n_18575)
);

INVx2_ASAP7_75t_L g18576 ( 
.A(n_18421),
.Y(n_18576)
);

INVx1_ASAP7_75t_SL g18577 ( 
.A(n_18447),
.Y(n_18577)
);

OR2x2_ASAP7_75t_L g18578 ( 
.A(n_18423),
.B(n_2883),
.Y(n_18578)
);

AND2x2_ASAP7_75t_L g18579 ( 
.A(n_18381),
.B(n_2883),
.Y(n_18579)
);

INVx2_ASAP7_75t_L g18580 ( 
.A(n_18427),
.Y(n_18580)
);

NOR3xp33_ASAP7_75t_L g18581 ( 
.A(n_18450),
.B(n_2884),
.C(n_2885),
.Y(n_18581)
);

BUFx3_ASAP7_75t_L g18582 ( 
.A(n_18429),
.Y(n_18582)
);

NOR2xp33_ASAP7_75t_L g18583 ( 
.A(n_18442),
.B(n_2884),
.Y(n_18583)
);

AO21x1_ASAP7_75t_L g18584 ( 
.A1(n_18449),
.A2(n_2885),
.B(n_2886),
.Y(n_18584)
);

OR2x2_ASAP7_75t_L g18585 ( 
.A(n_18390),
.B(n_2886),
.Y(n_18585)
);

NAND2xp5_ASAP7_75t_L g18586 ( 
.A(n_18398),
.B(n_2887),
.Y(n_18586)
);

BUFx3_ASAP7_75t_L g18587 ( 
.A(n_18342),
.Y(n_18587)
);

INVx1_ASAP7_75t_L g18588 ( 
.A(n_18343),
.Y(n_18588)
);

INVx1_ASAP7_75t_L g18589 ( 
.A(n_18343),
.Y(n_18589)
);

INVx3_ASAP7_75t_L g18590 ( 
.A(n_18339),
.Y(n_18590)
);

AND2x2_ASAP7_75t_L g18591 ( 
.A(n_18352),
.B(n_2888),
.Y(n_18591)
);

AOI22xp5_ASAP7_75t_L g18592 ( 
.A1(n_18355),
.A2(n_2890),
.B1(n_2888),
.B2(n_2889),
.Y(n_18592)
);

AND2x4_ASAP7_75t_L g18593 ( 
.A(n_18355),
.B(n_2889),
.Y(n_18593)
);

NOR2x1_ASAP7_75t_L g18594 ( 
.A(n_18339),
.B(n_2891),
.Y(n_18594)
);

OR2x2_ASAP7_75t_L g18595 ( 
.A(n_18463),
.B(n_2891),
.Y(n_18595)
);

NOR2xp33_ASAP7_75t_L g18596 ( 
.A(n_18475),
.B(n_2892),
.Y(n_18596)
);

INVx1_ASAP7_75t_L g18597 ( 
.A(n_18584),
.Y(n_18597)
);

INVx1_ASAP7_75t_L g18598 ( 
.A(n_18482),
.Y(n_18598)
);

INVx1_ASAP7_75t_L g18599 ( 
.A(n_18555),
.Y(n_18599)
);

AND2x2_ASAP7_75t_SL g18600 ( 
.A(n_18504),
.B(n_2892),
.Y(n_18600)
);

BUFx3_ASAP7_75t_L g18601 ( 
.A(n_18467),
.Y(n_18601)
);

INVx1_ASAP7_75t_SL g18602 ( 
.A(n_18562),
.Y(n_18602)
);

NAND3xp33_ASAP7_75t_SL g18603 ( 
.A(n_18539),
.B(n_2893),
.C(n_2894),
.Y(n_18603)
);

INVxp33_ASAP7_75t_SL g18604 ( 
.A(n_18502),
.Y(n_18604)
);

AOI22xp33_ASAP7_75t_L g18605 ( 
.A1(n_18587),
.A2(n_2896),
.B1(n_2893),
.B2(n_2895),
.Y(n_18605)
);

INVx1_ASAP7_75t_L g18606 ( 
.A(n_18553),
.Y(n_18606)
);

INVx1_ASAP7_75t_L g18607 ( 
.A(n_18533),
.Y(n_18607)
);

INVx1_ASAP7_75t_SL g18608 ( 
.A(n_18465),
.Y(n_18608)
);

NAND3xp33_ASAP7_75t_L g18609 ( 
.A(n_18594),
.B(n_2895),
.C(n_2896),
.Y(n_18609)
);

INVx1_ASAP7_75t_SL g18610 ( 
.A(n_18591),
.Y(n_18610)
);

INVxp67_ASAP7_75t_L g18611 ( 
.A(n_18481),
.Y(n_18611)
);

INVx1_ASAP7_75t_L g18612 ( 
.A(n_18546),
.Y(n_18612)
);

OAI211xp5_ASAP7_75t_SL g18613 ( 
.A1(n_18476),
.A2(n_2899),
.B(n_2897),
.C(n_2898),
.Y(n_18613)
);

OAI221xp5_ASAP7_75t_L g18614 ( 
.A1(n_18488),
.A2(n_18493),
.B1(n_18468),
.B2(n_18525),
.C(n_18526),
.Y(n_18614)
);

OAI21xp33_ASAP7_75t_L g18615 ( 
.A1(n_18511),
.A2(n_2897),
.B(n_2898),
.Y(n_18615)
);

AOI22xp5_ASAP7_75t_L g18616 ( 
.A1(n_18547),
.A2(n_2901),
.B1(n_2899),
.B2(n_2900),
.Y(n_18616)
);

AOI22xp5_ASAP7_75t_L g18617 ( 
.A1(n_18498),
.A2(n_18548),
.B1(n_18550),
.B2(n_18590),
.Y(n_18617)
);

NAND2xp5_ASAP7_75t_L g18618 ( 
.A(n_18554),
.B(n_18593),
.Y(n_18618)
);

AOI21xp33_ASAP7_75t_L g18619 ( 
.A1(n_18479),
.A2(n_2901),
.B(n_2902),
.Y(n_18619)
);

AOI21xp33_ASAP7_75t_L g18620 ( 
.A1(n_18572),
.A2(n_2902),
.B(n_2904),
.Y(n_18620)
);

NOR2xp67_ASAP7_75t_L g18621 ( 
.A(n_18561),
.B(n_2904),
.Y(n_18621)
);

INVx1_ASAP7_75t_SL g18622 ( 
.A(n_18507),
.Y(n_18622)
);

INVx1_ASAP7_75t_L g18623 ( 
.A(n_18564),
.Y(n_18623)
);

INVx1_ASAP7_75t_L g18624 ( 
.A(n_18496),
.Y(n_18624)
);

HB1xp67_ASAP7_75t_L g18625 ( 
.A(n_18518),
.Y(n_18625)
);

AOI22xp5_ASAP7_75t_L g18626 ( 
.A1(n_18559),
.A2(n_2907),
.B1(n_2905),
.B2(n_2906),
.Y(n_18626)
);

INVx1_ASAP7_75t_L g18627 ( 
.A(n_18531),
.Y(n_18627)
);

AND2x2_ASAP7_75t_L g18628 ( 
.A(n_18516),
.B(n_2905),
.Y(n_18628)
);

OAI31xp33_ASAP7_75t_L g18629 ( 
.A1(n_18489),
.A2(n_2909),
.A3(n_2907),
.B(n_2908),
.Y(n_18629)
);

NAND2xp5_ASAP7_75t_L g18630 ( 
.A(n_18469),
.B(n_2908),
.Y(n_18630)
);

NOR2xp33_ASAP7_75t_L g18631 ( 
.A(n_18510),
.B(n_2910),
.Y(n_18631)
);

NAND3xp33_ASAP7_75t_L g18632 ( 
.A(n_18492),
.B(n_2910),
.C(n_2911),
.Y(n_18632)
);

OAI32xp33_ASAP7_75t_L g18633 ( 
.A1(n_18513),
.A2(n_2913),
.A3(n_2911),
.B1(n_2912),
.B2(n_2914),
.Y(n_18633)
);

NAND2xp5_ASAP7_75t_L g18634 ( 
.A(n_18470),
.B(n_18477),
.Y(n_18634)
);

OAI22xp5_ASAP7_75t_L g18635 ( 
.A1(n_18505),
.A2(n_18483),
.B1(n_18577),
.B2(n_18509),
.Y(n_18635)
);

INVx1_ASAP7_75t_L g18636 ( 
.A(n_18568),
.Y(n_18636)
);

INVx2_ASAP7_75t_L g18637 ( 
.A(n_18527),
.Y(n_18637)
);

INVx1_ASAP7_75t_L g18638 ( 
.A(n_18520),
.Y(n_18638)
);

NAND2xp5_ASAP7_75t_L g18639 ( 
.A(n_18500),
.B(n_2912),
.Y(n_18639)
);

AND2x2_ASAP7_75t_L g18640 ( 
.A(n_18514),
.B(n_2913),
.Y(n_18640)
);

INVx1_ASAP7_75t_L g18641 ( 
.A(n_18578),
.Y(n_18641)
);

OAI32xp33_ASAP7_75t_L g18642 ( 
.A1(n_18494),
.A2(n_2916),
.A3(n_2914),
.B1(n_2915),
.B2(n_2917),
.Y(n_18642)
);

OAI22xp5_ASAP7_75t_L g18643 ( 
.A1(n_18544),
.A2(n_2917),
.B1(n_2915),
.B2(n_2916),
.Y(n_18643)
);

AOI21xp5_ASAP7_75t_L g18644 ( 
.A1(n_18517),
.A2(n_2918),
.B(n_2919),
.Y(n_18644)
);

INVxp67_ASAP7_75t_L g18645 ( 
.A(n_18583),
.Y(n_18645)
);

INVx2_ASAP7_75t_L g18646 ( 
.A(n_18563),
.Y(n_18646)
);

AOI21xp33_ASAP7_75t_L g18647 ( 
.A1(n_18512),
.A2(n_2919),
.B(n_2920),
.Y(n_18647)
);

INVx1_ASAP7_75t_L g18648 ( 
.A(n_18595),
.Y(n_18648)
);

AOI22xp5_ASAP7_75t_L g18649 ( 
.A1(n_18565),
.A2(n_2922),
.B1(n_2920),
.B2(n_2921),
.Y(n_18649)
);

NAND2xp5_ASAP7_75t_L g18650 ( 
.A(n_18499),
.B(n_2921),
.Y(n_18650)
);

INVx2_ASAP7_75t_L g18651 ( 
.A(n_18515),
.Y(n_18651)
);

AOI222xp33_ASAP7_75t_L g18652 ( 
.A1(n_18573),
.A2(n_2924),
.B1(n_2926),
.B2(n_2922),
.C1(n_2923),
.C2(n_2925),
.Y(n_18652)
);

AND2x2_ASAP7_75t_L g18653 ( 
.A(n_18472),
.B(n_2923),
.Y(n_18653)
);

AOI21xp5_ASAP7_75t_L g18654 ( 
.A1(n_18534),
.A2(n_2924),
.B(n_2925),
.Y(n_18654)
);

AOI222xp33_ASAP7_75t_L g18655 ( 
.A1(n_18508),
.A2(n_2928),
.B1(n_2930),
.B2(n_2926),
.C1(n_2927),
.C2(n_2929),
.Y(n_18655)
);

OAI22xp5_ASAP7_75t_L g18656 ( 
.A1(n_18473),
.A2(n_2929),
.B1(n_2927),
.B2(n_2928),
.Y(n_18656)
);

NOR2xp33_ASAP7_75t_L g18657 ( 
.A(n_18588),
.B(n_18589),
.Y(n_18657)
);

INVxp33_ASAP7_75t_L g18658 ( 
.A(n_18536),
.Y(n_18658)
);

NAND3xp33_ASAP7_75t_L g18659 ( 
.A(n_18497),
.B(n_2930),
.C(n_2931),
.Y(n_18659)
);

NAND2xp5_ASAP7_75t_L g18660 ( 
.A(n_18501),
.B(n_18579),
.Y(n_18660)
);

NAND2xp5_ASAP7_75t_L g18661 ( 
.A(n_18471),
.B(n_2932),
.Y(n_18661)
);

OAI21xp5_ASAP7_75t_SL g18662 ( 
.A1(n_18503),
.A2(n_18495),
.B(n_18574),
.Y(n_18662)
);

NAND2xp5_ASAP7_75t_SL g18663 ( 
.A(n_18567),
.B(n_2932),
.Y(n_18663)
);

AOI22xp5_ASAP7_75t_L g18664 ( 
.A1(n_18570),
.A2(n_2935),
.B1(n_2933),
.B2(n_2934),
.Y(n_18664)
);

INVx1_ASAP7_75t_L g18665 ( 
.A(n_18487),
.Y(n_18665)
);

AOI211xp5_ASAP7_75t_L g18666 ( 
.A1(n_18530),
.A2(n_2936),
.B(n_2933),
.C(n_2934),
.Y(n_18666)
);

NAND3xp33_ASAP7_75t_SL g18667 ( 
.A(n_18478),
.B(n_2936),
.C(n_2937),
.Y(n_18667)
);

INVx2_ASAP7_75t_L g18668 ( 
.A(n_18543),
.Y(n_18668)
);

INVx1_ASAP7_75t_L g18669 ( 
.A(n_18486),
.Y(n_18669)
);

AND2x2_ASAP7_75t_L g18670 ( 
.A(n_18519),
.B(n_2937),
.Y(n_18670)
);

NAND2xp5_ASAP7_75t_L g18671 ( 
.A(n_18581),
.B(n_2938),
.Y(n_18671)
);

AND2x4_ASAP7_75t_L g18672 ( 
.A(n_18485),
.B(n_18491),
.Y(n_18672)
);

A2O1A1Ixp33_ASAP7_75t_L g18673 ( 
.A1(n_18556),
.A2(n_2941),
.B(n_2938),
.C(n_2940),
.Y(n_18673)
);

AND2x2_ASAP7_75t_L g18674 ( 
.A(n_18490),
.B(n_2940),
.Y(n_18674)
);

AND2x2_ASAP7_75t_L g18675 ( 
.A(n_18523),
.B(n_2941),
.Y(n_18675)
);

OAI322xp33_ASAP7_75t_L g18676 ( 
.A1(n_18571),
.A2(n_2947),
.A3(n_2946),
.B1(n_2944),
.B2(n_2942),
.C1(n_2943),
.C2(n_2945),
.Y(n_18676)
);

NOR2xp67_ASAP7_75t_L g18677 ( 
.A(n_18466),
.B(n_2942),
.Y(n_18677)
);

OAI221xp5_ASAP7_75t_L g18678 ( 
.A1(n_18586),
.A2(n_18575),
.B1(n_18566),
.B2(n_18545),
.C(n_18585),
.Y(n_18678)
);

INVx1_ASAP7_75t_L g18679 ( 
.A(n_18560),
.Y(n_18679)
);

NOR2xp67_ASAP7_75t_L g18680 ( 
.A(n_18592),
.B(n_2943),
.Y(n_18680)
);

AND2x2_ASAP7_75t_L g18681 ( 
.A(n_18474),
.B(n_2945),
.Y(n_18681)
);

NOR2xp33_ASAP7_75t_L g18682 ( 
.A(n_18506),
.B(n_2946),
.Y(n_18682)
);

INVxp67_ASAP7_75t_SL g18683 ( 
.A(n_18532),
.Y(n_18683)
);

OAI22xp5_ASAP7_75t_L g18684 ( 
.A1(n_18576),
.A2(n_2950),
.B1(n_2947),
.B2(n_2948),
.Y(n_18684)
);

AOI21xp5_ASAP7_75t_L g18685 ( 
.A1(n_18484),
.A2(n_2948),
.B(n_2950),
.Y(n_18685)
);

AOI22xp33_ASAP7_75t_SL g18686 ( 
.A1(n_18582),
.A2(n_2953),
.B1(n_2951),
.B2(n_2952),
.Y(n_18686)
);

OR2x2_ASAP7_75t_L g18687 ( 
.A(n_18535),
.B(n_2951),
.Y(n_18687)
);

AND2x2_ASAP7_75t_L g18688 ( 
.A(n_18521),
.B(n_2954),
.Y(n_18688)
);

AOI22xp5_ASAP7_75t_L g18689 ( 
.A1(n_18580),
.A2(n_2956),
.B1(n_2954),
.B2(n_2955),
.Y(n_18689)
);

AOI221xp5_ASAP7_75t_L g18690 ( 
.A1(n_18524),
.A2(n_2957),
.B1(n_2955),
.B2(n_2956),
.C(n_2958),
.Y(n_18690)
);

AOI22xp5_ASAP7_75t_L g18691 ( 
.A1(n_18558),
.A2(n_2960),
.B1(n_2958),
.B2(n_2959),
.Y(n_18691)
);

NAND2xp5_ASAP7_75t_L g18692 ( 
.A(n_18480),
.B(n_2959),
.Y(n_18692)
);

INVx1_ASAP7_75t_L g18693 ( 
.A(n_18529),
.Y(n_18693)
);

INVx1_ASAP7_75t_L g18694 ( 
.A(n_18528),
.Y(n_18694)
);

AOI21xp33_ASAP7_75t_L g18695 ( 
.A1(n_18522),
.A2(n_2960),
.B(n_2961),
.Y(n_18695)
);

AOI21xp33_ASAP7_75t_L g18696 ( 
.A1(n_18538),
.A2(n_2961),
.B(n_2962),
.Y(n_18696)
);

OAI221xp5_ASAP7_75t_L g18697 ( 
.A1(n_18569),
.A2(n_2964),
.B1(n_2962),
.B2(n_2963),
.C(n_2965),
.Y(n_18697)
);

NAND2xp5_ASAP7_75t_L g18698 ( 
.A(n_18549),
.B(n_2963),
.Y(n_18698)
);

NOR3xp33_ASAP7_75t_SL g18699 ( 
.A(n_18557),
.B(n_2964),
.C(n_2965),
.Y(n_18699)
);

NOR2xp33_ASAP7_75t_SL g18700 ( 
.A(n_18537),
.B(n_2966),
.Y(n_18700)
);

AOI22xp5_ASAP7_75t_L g18701 ( 
.A1(n_18551),
.A2(n_2969),
.B1(n_2967),
.B2(n_2968),
.Y(n_18701)
);

NOR2xp33_ASAP7_75t_L g18702 ( 
.A(n_18540),
.B(n_18541),
.Y(n_18702)
);

INVx1_ASAP7_75t_L g18703 ( 
.A(n_18542),
.Y(n_18703)
);

AND2x2_ASAP7_75t_L g18704 ( 
.A(n_18552),
.B(n_2967),
.Y(n_18704)
);

AOI22xp5_ASAP7_75t_L g18705 ( 
.A1(n_18467),
.A2(n_2971),
.B1(n_2969),
.B2(n_2970),
.Y(n_18705)
);

INVx2_ASAP7_75t_L g18706 ( 
.A(n_18587),
.Y(n_18706)
);

INVx1_ASAP7_75t_L g18707 ( 
.A(n_18584),
.Y(n_18707)
);

INVxp67_ASAP7_75t_SL g18708 ( 
.A(n_18554),
.Y(n_18708)
);

INVx1_ASAP7_75t_L g18709 ( 
.A(n_18584),
.Y(n_18709)
);

INVx1_ASAP7_75t_SL g18710 ( 
.A(n_18482),
.Y(n_18710)
);

OAI22xp5_ASAP7_75t_L g18711 ( 
.A1(n_18467),
.A2(n_2973),
.B1(n_2970),
.B2(n_2972),
.Y(n_18711)
);

OR2x2_ASAP7_75t_L g18712 ( 
.A(n_18475),
.B(n_2972),
.Y(n_18712)
);

NAND3x2_ASAP7_75t_L g18713 ( 
.A(n_18573),
.B(n_2973),
.C(n_2974),
.Y(n_18713)
);

INVx2_ASAP7_75t_L g18714 ( 
.A(n_18587),
.Y(n_18714)
);

INVx1_ASAP7_75t_L g18715 ( 
.A(n_18584),
.Y(n_18715)
);

INVx3_ASAP7_75t_L g18716 ( 
.A(n_18475),
.Y(n_18716)
);

AOI22xp5_ASAP7_75t_L g18717 ( 
.A1(n_18716),
.A2(n_2976),
.B1(n_2974),
.B2(n_2975),
.Y(n_18717)
);

AOI221xp5_ASAP7_75t_L g18718 ( 
.A1(n_18635),
.A2(n_2977),
.B1(n_2975),
.B2(n_2976),
.C(n_2978),
.Y(n_18718)
);

INVx1_ASAP7_75t_L g18719 ( 
.A(n_18600),
.Y(n_18719)
);

OAI22xp33_ASAP7_75t_L g18720 ( 
.A1(n_18617),
.A2(n_2981),
.B1(n_2979),
.B2(n_2980),
.Y(n_18720)
);

OAI221xp5_ASAP7_75t_L g18721 ( 
.A1(n_18662),
.A2(n_2982),
.B1(n_2980),
.B2(n_2981),
.C(n_2983),
.Y(n_18721)
);

OAI21xp5_ASAP7_75t_L g18722 ( 
.A1(n_18596),
.A2(n_2982),
.B(n_2983),
.Y(n_18722)
);

OAI22xp33_ASAP7_75t_SL g18723 ( 
.A1(n_18597),
.A2(n_2986),
.B1(n_2984),
.B2(n_2985),
.Y(n_18723)
);

OAI21xp33_ASAP7_75t_SL g18724 ( 
.A1(n_18683),
.A2(n_18709),
.B(n_18707),
.Y(n_18724)
);

INVx1_ASAP7_75t_L g18725 ( 
.A(n_18712),
.Y(n_18725)
);

AOI21xp33_ASAP7_75t_SL g18726 ( 
.A1(n_18715),
.A2(n_2984),
.B(n_2985),
.Y(n_18726)
);

NOR2xp33_ASAP7_75t_SL g18727 ( 
.A(n_18602),
.B(n_2986),
.Y(n_18727)
);

INVx1_ASAP7_75t_L g18728 ( 
.A(n_18628),
.Y(n_18728)
);

XNOR2xp5_ASAP7_75t_L g18729 ( 
.A(n_18601),
.B(n_18713),
.Y(n_18729)
);

INVx1_ASAP7_75t_L g18730 ( 
.A(n_18653),
.Y(n_18730)
);

NAND3xp33_ASAP7_75t_L g18731 ( 
.A(n_18666),
.B(n_2987),
.C(n_2988),
.Y(n_18731)
);

AOI22xp33_ASAP7_75t_L g18732 ( 
.A1(n_18716),
.A2(n_2990),
.B1(n_2987),
.B2(n_2989),
.Y(n_18732)
);

AOI22xp5_ASAP7_75t_L g18733 ( 
.A1(n_18604),
.A2(n_2991),
.B1(n_2989),
.B2(n_2990),
.Y(n_18733)
);

INVx1_ASAP7_75t_L g18734 ( 
.A(n_18640),
.Y(n_18734)
);

OAI221xp5_ASAP7_75t_SL g18735 ( 
.A1(n_18614),
.A2(n_2993),
.B1(n_2991),
.B2(n_2992),
.C(n_2994),
.Y(n_18735)
);

OAI21xp33_ASAP7_75t_L g18736 ( 
.A1(n_18657),
.A2(n_2992),
.B(n_2993),
.Y(n_18736)
);

OAI22x1_ASAP7_75t_L g18737 ( 
.A1(n_18708),
.A2(n_2996),
.B1(n_2994),
.B2(n_2995),
.Y(n_18737)
);

INVx1_ASAP7_75t_L g18738 ( 
.A(n_18674),
.Y(n_18738)
);

NAND3xp33_ASAP7_75t_L g18739 ( 
.A(n_18699),
.B(n_2995),
.C(n_2996),
.Y(n_18739)
);

NAND2xp5_ASAP7_75t_L g18740 ( 
.A(n_18670),
.B(n_2997),
.Y(n_18740)
);

INVx1_ASAP7_75t_L g18741 ( 
.A(n_18675),
.Y(n_18741)
);

OAI22xp5_ASAP7_75t_L g18742 ( 
.A1(n_18625),
.A2(n_2999),
.B1(n_2997),
.B2(n_2998),
.Y(n_18742)
);

INVx1_ASAP7_75t_L g18743 ( 
.A(n_18681),
.Y(n_18743)
);

INVx2_ASAP7_75t_L g18744 ( 
.A(n_18688),
.Y(n_18744)
);

AOI21xp5_ASAP7_75t_L g18745 ( 
.A1(n_18618),
.A2(n_2998),
.B(n_2999),
.Y(n_18745)
);

INVx1_ASAP7_75t_L g18746 ( 
.A(n_18704),
.Y(n_18746)
);

OAI22xp33_ASAP7_75t_L g18747 ( 
.A1(n_18658),
.A2(n_3002),
.B1(n_3000),
.B2(n_3001),
.Y(n_18747)
);

AND2x2_ASAP7_75t_L g18748 ( 
.A(n_18706),
.B(n_3000),
.Y(n_18748)
);

INVx1_ASAP7_75t_L g18749 ( 
.A(n_18650),
.Y(n_18749)
);

AOI221xp5_ASAP7_75t_L g18750 ( 
.A1(n_18693),
.A2(n_3004),
.B1(n_3001),
.B2(n_3003),
.C(n_3005),
.Y(n_18750)
);

NAND2xp5_ASAP7_75t_L g18751 ( 
.A(n_18631),
.B(n_3004),
.Y(n_18751)
);

NOR2xp33_ASAP7_75t_L g18752 ( 
.A(n_18613),
.B(n_18710),
.Y(n_18752)
);

AOI21xp33_ASAP7_75t_L g18753 ( 
.A1(n_18606),
.A2(n_3006),
.B(n_3007),
.Y(n_18753)
);

OAI22xp5_ASAP7_75t_L g18754 ( 
.A1(n_18611),
.A2(n_3009),
.B1(n_3006),
.B2(n_3008),
.Y(n_18754)
);

INVxp67_ASAP7_75t_SL g18755 ( 
.A(n_18609),
.Y(n_18755)
);

NOR2xp33_ASAP7_75t_SL g18756 ( 
.A(n_18676),
.B(n_3008),
.Y(n_18756)
);

INVx1_ASAP7_75t_L g18757 ( 
.A(n_18630),
.Y(n_18757)
);

BUFx6f_ASAP7_75t_L g18758 ( 
.A(n_18672),
.Y(n_18758)
);

OR2x2_ASAP7_75t_L g18759 ( 
.A(n_18603),
.B(n_3009),
.Y(n_18759)
);

INVx1_ASAP7_75t_L g18760 ( 
.A(n_18639),
.Y(n_18760)
);

AOI211xp5_ASAP7_75t_L g18761 ( 
.A1(n_18667),
.A2(n_3012),
.B(n_3010),
.C(n_3011),
.Y(n_18761)
);

INVx1_ASAP7_75t_L g18762 ( 
.A(n_18687),
.Y(n_18762)
);

AOI221xp5_ASAP7_75t_L g18763 ( 
.A1(n_18694),
.A2(n_3014),
.B1(n_3012),
.B2(n_3013),
.C(n_3015),
.Y(n_18763)
);

AOI22xp5_ASAP7_75t_L g18764 ( 
.A1(n_18714),
.A2(n_18672),
.B1(n_18622),
.B2(n_18608),
.Y(n_18764)
);

A2O1A1Ixp33_ASAP7_75t_L g18765 ( 
.A1(n_18629),
.A2(n_3015),
.B(n_3013),
.C(n_3014),
.Y(n_18765)
);

AND2x2_ASAP7_75t_L g18766 ( 
.A(n_18598),
.B(n_3016),
.Y(n_18766)
);

INVx1_ASAP7_75t_L g18767 ( 
.A(n_18698),
.Y(n_18767)
);

NOR2xp33_ASAP7_75t_L g18768 ( 
.A(n_18610),
.B(n_3016),
.Y(n_18768)
);

NAND2xp5_ASAP7_75t_L g18769 ( 
.A(n_18686),
.B(n_3017),
.Y(n_18769)
);

NAND2xp5_ASAP7_75t_L g18770 ( 
.A(n_18644),
.B(n_3017),
.Y(n_18770)
);

INVx2_ASAP7_75t_L g18771 ( 
.A(n_18637),
.Y(n_18771)
);

A2O1A1Ixp33_ASAP7_75t_L g18772 ( 
.A1(n_18682),
.A2(n_3020),
.B(n_3018),
.C(n_3019),
.Y(n_18772)
);

OAI221xp5_ASAP7_75t_L g18773 ( 
.A1(n_18673),
.A2(n_18661),
.B1(n_18659),
.B2(n_18632),
.C(n_18671),
.Y(n_18773)
);

OAI21xp33_ASAP7_75t_L g18774 ( 
.A1(n_18634),
.A2(n_3019),
.B(n_3020),
.Y(n_18774)
);

OAI22xp5_ASAP7_75t_L g18775 ( 
.A1(n_18692),
.A2(n_3023),
.B1(n_3021),
.B2(n_3022),
.Y(n_18775)
);

INVx1_ASAP7_75t_L g18776 ( 
.A(n_18663),
.Y(n_18776)
);

INVx1_ASAP7_75t_SL g18777 ( 
.A(n_18660),
.Y(n_18777)
);

BUFx3_ASAP7_75t_L g18778 ( 
.A(n_18646),
.Y(n_18778)
);

AOI211xp5_ASAP7_75t_L g18779 ( 
.A1(n_18643),
.A2(n_3024),
.B(n_3022),
.C(n_3023),
.Y(n_18779)
);

AOI221xp5_ASAP7_75t_L g18780 ( 
.A1(n_18678),
.A2(n_3026),
.B1(n_3024),
.B2(n_3025),
.C(n_3027),
.Y(n_18780)
);

NOR2x1_ASAP7_75t_L g18781 ( 
.A(n_18648),
.B(n_3025),
.Y(n_18781)
);

NAND2xp5_ASAP7_75t_L g18782 ( 
.A(n_18685),
.B(n_3026),
.Y(n_18782)
);

AOI31xp33_ASAP7_75t_L g18783 ( 
.A1(n_18638),
.A2(n_3029),
.A3(n_3027),
.B(n_3028),
.Y(n_18783)
);

OR2x2_ASAP7_75t_L g18784 ( 
.A(n_18607),
.B(n_18612),
.Y(n_18784)
);

NOR2xp33_ASAP7_75t_L g18785 ( 
.A(n_18615),
.B(n_3028),
.Y(n_18785)
);

OAI221xp5_ASAP7_75t_L g18786 ( 
.A1(n_18621),
.A2(n_3031),
.B1(n_3029),
.B2(n_3030),
.C(n_3032),
.Y(n_18786)
);

INVx1_ASAP7_75t_L g18787 ( 
.A(n_18623),
.Y(n_18787)
);

INVx1_ASAP7_75t_L g18788 ( 
.A(n_18624),
.Y(n_18788)
);

NAND2xp5_ASAP7_75t_L g18789 ( 
.A(n_18700),
.B(n_18652),
.Y(n_18789)
);

INVx1_ASAP7_75t_L g18790 ( 
.A(n_18627),
.Y(n_18790)
);

NAND2xp5_ASAP7_75t_L g18791 ( 
.A(n_18649),
.B(n_3031),
.Y(n_18791)
);

NAND2xp5_ASAP7_75t_L g18792 ( 
.A(n_18677),
.B(n_3032),
.Y(n_18792)
);

INVx1_ASAP7_75t_L g18793 ( 
.A(n_18633),
.Y(n_18793)
);

AOI22xp5_ASAP7_75t_L g18794 ( 
.A1(n_18599),
.A2(n_3035),
.B1(n_3033),
.B2(n_3034),
.Y(n_18794)
);

AOI322xp5_ASAP7_75t_L g18795 ( 
.A1(n_18702),
.A2(n_3038),
.A3(n_3037),
.B1(n_3035),
.B2(n_3033),
.C1(n_3034),
.C2(n_3036),
.Y(n_18795)
);

AOI21x1_ASAP7_75t_L g18796 ( 
.A1(n_18654),
.A2(n_3036),
.B(n_3037),
.Y(n_18796)
);

OR2x2_ASAP7_75t_L g18797 ( 
.A(n_18668),
.B(n_3038),
.Y(n_18797)
);

INVxp67_ASAP7_75t_SL g18798 ( 
.A(n_18616),
.Y(n_18798)
);

OAI22xp33_ASAP7_75t_L g18799 ( 
.A1(n_18680),
.A2(n_3041),
.B1(n_3039),
.B2(n_3040),
.Y(n_18799)
);

OAI211xp5_ASAP7_75t_L g18800 ( 
.A1(n_18620),
.A2(n_3042),
.B(n_3039),
.C(n_3041),
.Y(n_18800)
);

OAI222xp33_ASAP7_75t_L g18801 ( 
.A1(n_18703),
.A2(n_3044),
.B1(n_3046),
.B2(n_3042),
.C1(n_3043),
.C2(n_3045),
.Y(n_18801)
);

INVx1_ASAP7_75t_L g18802 ( 
.A(n_18636),
.Y(n_18802)
);

INVxp67_ASAP7_75t_L g18803 ( 
.A(n_18697),
.Y(n_18803)
);

INVxp67_ASAP7_75t_L g18804 ( 
.A(n_18711),
.Y(n_18804)
);

INVx1_ASAP7_75t_L g18805 ( 
.A(n_18651),
.Y(n_18805)
);

INVx1_ASAP7_75t_L g18806 ( 
.A(n_18641),
.Y(n_18806)
);

INVx2_ASAP7_75t_L g18807 ( 
.A(n_18665),
.Y(n_18807)
);

NAND2xp5_ASAP7_75t_L g18808 ( 
.A(n_18655),
.B(n_3043),
.Y(n_18808)
);

OAI32xp33_ASAP7_75t_L g18809 ( 
.A1(n_18679),
.A2(n_3049),
.A3(n_3047),
.B1(n_3048),
.B2(n_3050),
.Y(n_18809)
);

OAI221xp5_ASAP7_75t_L g18810 ( 
.A1(n_18645),
.A2(n_3049),
.B1(n_3047),
.B2(n_3048),
.C(n_3051),
.Y(n_18810)
);

OAI21xp5_ASAP7_75t_L g18811 ( 
.A1(n_18669),
.A2(n_3051),
.B(n_3052),
.Y(n_18811)
);

NAND2xp5_ASAP7_75t_L g18812 ( 
.A(n_18690),
.B(n_3053),
.Y(n_18812)
);

NAND3xp33_ASAP7_75t_SL g18813 ( 
.A(n_18664),
.B(n_18689),
.C(n_18605),
.Y(n_18813)
);

INVx1_ASAP7_75t_L g18814 ( 
.A(n_18642),
.Y(n_18814)
);

INVx1_ASAP7_75t_L g18815 ( 
.A(n_18684),
.Y(n_18815)
);

AOI21xp5_ASAP7_75t_L g18816 ( 
.A1(n_18619),
.A2(n_3053),
.B(n_3054),
.Y(n_18816)
);

INVx1_ASAP7_75t_L g18817 ( 
.A(n_18626),
.Y(n_18817)
);

OAI22xp5_ASAP7_75t_L g18818 ( 
.A1(n_18705),
.A2(n_3056),
.B1(n_3054),
.B2(n_3055),
.Y(n_18818)
);

OAI221xp5_ASAP7_75t_L g18819 ( 
.A1(n_18647),
.A2(n_3057),
.B1(n_3055),
.B2(n_3056),
.C(n_3058),
.Y(n_18819)
);

AND2x2_ASAP7_75t_L g18820 ( 
.A(n_18696),
.B(n_3057),
.Y(n_18820)
);

INVxp67_ASAP7_75t_L g18821 ( 
.A(n_18656),
.Y(n_18821)
);

NAND2xp5_ASAP7_75t_L g18822 ( 
.A(n_18691),
.B(n_3058),
.Y(n_18822)
);

INVx1_ASAP7_75t_L g18823 ( 
.A(n_18701),
.Y(n_18823)
);

AOI21xp5_ASAP7_75t_L g18824 ( 
.A1(n_18695),
.A2(n_3059),
.B(n_3060),
.Y(n_18824)
);

NOR2xp33_ASAP7_75t_R g18825 ( 
.A(n_18716),
.B(n_3059),
.Y(n_18825)
);

OAI22xp5_ASAP7_75t_L g18826 ( 
.A1(n_18617),
.A2(n_3063),
.B1(n_3060),
.B2(n_3062),
.Y(n_18826)
);

AOI22xp5_ASAP7_75t_L g18827 ( 
.A1(n_18716),
.A2(n_3064),
.B1(n_3062),
.B2(n_3063),
.Y(n_18827)
);

OR2x2_ASAP7_75t_L g18828 ( 
.A(n_18712),
.B(n_3064),
.Y(n_18828)
);

A2O1A1Ixp33_ASAP7_75t_L g18829 ( 
.A1(n_18596),
.A2(n_3067),
.B(n_3065),
.C(n_3066),
.Y(n_18829)
);

NOR2xp33_ASAP7_75t_R g18830 ( 
.A(n_18716),
.B(n_3065),
.Y(n_18830)
);

OAI21xp33_ASAP7_75t_SL g18831 ( 
.A1(n_18617),
.A2(n_3066),
.B(n_3067),
.Y(n_18831)
);

AOI222xp33_ASAP7_75t_L g18832 ( 
.A1(n_18601),
.A2(n_3070),
.B1(n_3072),
.B2(n_3068),
.C1(n_3069),
.C2(n_3071),
.Y(n_18832)
);

NAND3xp33_ASAP7_75t_L g18833 ( 
.A(n_18617),
.B(n_3068),
.C(n_3069),
.Y(n_18833)
);

XOR2xp5_ASAP7_75t_L g18834 ( 
.A(n_18729),
.B(n_3072),
.Y(n_18834)
);

AOI221xp5_ASAP7_75t_L g18835 ( 
.A1(n_18724),
.A2(n_3075),
.B1(n_3073),
.B2(n_3074),
.C(n_3076),
.Y(n_18835)
);

AND2x2_ASAP7_75t_L g18836 ( 
.A(n_18771),
.B(n_3073),
.Y(n_18836)
);

INVx1_ASAP7_75t_L g18837 ( 
.A(n_18758),
.Y(n_18837)
);

OAI22xp5_ASAP7_75t_L g18838 ( 
.A1(n_18764),
.A2(n_3077),
.B1(n_3074),
.B2(n_3075),
.Y(n_18838)
);

INVx1_ASAP7_75t_L g18839 ( 
.A(n_18758),
.Y(n_18839)
);

INVx1_ASAP7_75t_SL g18840 ( 
.A(n_18825),
.Y(n_18840)
);

NAND2xp5_ASAP7_75t_L g18841 ( 
.A(n_18758),
.B(n_3077),
.Y(n_18841)
);

INVx1_ASAP7_75t_L g18842 ( 
.A(n_18781),
.Y(n_18842)
);

INVxp67_ASAP7_75t_L g18843 ( 
.A(n_18727),
.Y(n_18843)
);

NAND2xp5_ASAP7_75t_L g18844 ( 
.A(n_18766),
.B(n_3078),
.Y(n_18844)
);

INVxp67_ASAP7_75t_SL g18845 ( 
.A(n_18737),
.Y(n_18845)
);

OR2x2_ASAP7_75t_L g18846 ( 
.A(n_18828),
.B(n_3078),
.Y(n_18846)
);

NOR2xp33_ASAP7_75t_L g18847 ( 
.A(n_18735),
.B(n_3079),
.Y(n_18847)
);

INVx1_ASAP7_75t_L g18848 ( 
.A(n_18748),
.Y(n_18848)
);

AND2x2_ASAP7_75t_L g18849 ( 
.A(n_18778),
.B(n_3079),
.Y(n_18849)
);

NOR2xp33_ASAP7_75t_L g18850 ( 
.A(n_18831),
.B(n_3080),
.Y(n_18850)
);

INVx1_ASAP7_75t_L g18851 ( 
.A(n_18797),
.Y(n_18851)
);

NOR2xp33_ASAP7_75t_L g18852 ( 
.A(n_18800),
.B(n_3080),
.Y(n_18852)
);

INVx3_ASAP7_75t_L g18853 ( 
.A(n_18796),
.Y(n_18853)
);

AND2x2_ASAP7_75t_L g18854 ( 
.A(n_18719),
.B(n_18728),
.Y(n_18854)
);

HB1xp67_ASAP7_75t_SL g18855 ( 
.A(n_18784),
.Y(n_18855)
);

OR2x2_ASAP7_75t_L g18856 ( 
.A(n_18759),
.B(n_3081),
.Y(n_18856)
);

OR2x2_ASAP7_75t_L g18857 ( 
.A(n_18740),
.B(n_3081),
.Y(n_18857)
);

OAI221xp5_ASAP7_75t_SL g18858 ( 
.A1(n_18718),
.A2(n_18777),
.B1(n_18821),
.B2(n_18808),
.C(n_18804),
.Y(n_18858)
);

AOI221xp5_ASAP7_75t_L g18859 ( 
.A1(n_18752),
.A2(n_18814),
.B1(n_18793),
.B2(n_18739),
.C(n_18805),
.Y(n_18859)
);

NAND2xp5_ASAP7_75t_L g18860 ( 
.A(n_18726),
.B(n_3082),
.Y(n_18860)
);

INVx1_ASAP7_75t_SL g18861 ( 
.A(n_18830),
.Y(n_18861)
);

AND2x2_ASAP7_75t_L g18862 ( 
.A(n_18734),
.B(n_3082),
.Y(n_18862)
);

NOR2xp33_ASAP7_75t_L g18863 ( 
.A(n_18786),
.B(n_3083),
.Y(n_18863)
);

INVx2_ASAP7_75t_L g18864 ( 
.A(n_18744),
.Y(n_18864)
);

BUFx2_ASAP7_75t_L g18865 ( 
.A(n_18811),
.Y(n_18865)
);

INVx1_ASAP7_75t_SL g18866 ( 
.A(n_18792),
.Y(n_18866)
);

NAND2xp5_ASAP7_75t_SL g18867 ( 
.A(n_18723),
.B(n_3084),
.Y(n_18867)
);

INVx1_ASAP7_75t_L g18868 ( 
.A(n_18768),
.Y(n_18868)
);

AOI221x1_ASAP7_75t_SL g18869 ( 
.A1(n_18789),
.A2(n_3086),
.B1(n_3084),
.B2(n_3085),
.C(n_3087),
.Y(n_18869)
);

INVx1_ASAP7_75t_SL g18870 ( 
.A(n_18770),
.Y(n_18870)
);

INVx1_ASAP7_75t_L g18871 ( 
.A(n_18769),
.Y(n_18871)
);

NAND2xp5_ASAP7_75t_L g18872 ( 
.A(n_18783),
.B(n_3085),
.Y(n_18872)
);

NAND2xp5_ASAP7_75t_L g18873 ( 
.A(n_18720),
.B(n_3087),
.Y(n_18873)
);

INVx1_ASAP7_75t_L g18874 ( 
.A(n_18833),
.Y(n_18874)
);

INVx2_ASAP7_75t_L g18875 ( 
.A(n_18820),
.Y(n_18875)
);

NAND2xp5_ASAP7_75t_L g18876 ( 
.A(n_18829),
.B(n_3088),
.Y(n_18876)
);

OR2x2_ASAP7_75t_L g18877 ( 
.A(n_18751),
.B(n_3088),
.Y(n_18877)
);

INVx1_ASAP7_75t_L g18878 ( 
.A(n_18782),
.Y(n_18878)
);

INVx1_ASAP7_75t_L g18879 ( 
.A(n_18812),
.Y(n_18879)
);

OR2x2_ASAP7_75t_L g18880 ( 
.A(n_18791),
.B(n_3089),
.Y(n_18880)
);

NAND2xp5_ASAP7_75t_L g18881 ( 
.A(n_18774),
.B(n_3089),
.Y(n_18881)
);

NOR2x1_ASAP7_75t_L g18882 ( 
.A(n_18801),
.B(n_3090),
.Y(n_18882)
);

AND2x2_ASAP7_75t_L g18883 ( 
.A(n_18730),
.B(n_3090),
.Y(n_18883)
);

NAND2xp5_ASAP7_75t_L g18884 ( 
.A(n_18761),
.B(n_3091),
.Y(n_18884)
);

AND2x2_ASAP7_75t_L g18885 ( 
.A(n_18738),
.B(n_3091),
.Y(n_18885)
);

OR2x2_ASAP7_75t_L g18886 ( 
.A(n_18818),
.B(n_3092),
.Y(n_18886)
);

INVx2_ASAP7_75t_L g18887 ( 
.A(n_18746),
.Y(n_18887)
);

NAND2xp5_ASAP7_75t_L g18888 ( 
.A(n_18736),
.B(n_3092),
.Y(n_18888)
);

AOI222xp33_ASAP7_75t_L g18889 ( 
.A1(n_18813),
.A2(n_18806),
.B1(n_18787),
.B2(n_18788),
.C1(n_18802),
.C2(n_18790),
.Y(n_18889)
);

INVx4_ASAP7_75t_L g18890 ( 
.A(n_18807),
.Y(n_18890)
);

NAND2xp5_ASAP7_75t_L g18891 ( 
.A(n_18799),
.B(n_3093),
.Y(n_18891)
);

NAND2xp5_ASAP7_75t_SL g18892 ( 
.A(n_18779),
.B(n_3093),
.Y(n_18892)
);

NAND2xp5_ASAP7_75t_L g18893 ( 
.A(n_18745),
.B(n_3094),
.Y(n_18893)
);

AND2x2_ASAP7_75t_L g18894 ( 
.A(n_18725),
.B(n_3094),
.Y(n_18894)
);

INVx1_ASAP7_75t_SL g18895 ( 
.A(n_18822),
.Y(n_18895)
);

INVxp67_ASAP7_75t_L g18896 ( 
.A(n_18756),
.Y(n_18896)
);

AND2x2_ASAP7_75t_L g18897 ( 
.A(n_18741),
.B(n_18743),
.Y(n_18897)
);

AND2x2_ASAP7_75t_L g18898 ( 
.A(n_18722),
.B(n_3095),
.Y(n_18898)
);

HB1xp67_ASAP7_75t_L g18899 ( 
.A(n_18742),
.Y(n_18899)
);

INVx2_ASAP7_75t_SL g18900 ( 
.A(n_18762),
.Y(n_18900)
);

INVx1_ASAP7_75t_L g18901 ( 
.A(n_18785),
.Y(n_18901)
);

INVx1_ASAP7_75t_L g18902 ( 
.A(n_18775),
.Y(n_18902)
);

AOI22xp5_ASAP7_75t_L g18903 ( 
.A1(n_18755),
.A2(n_3097),
.B1(n_3095),
.B2(n_3096),
.Y(n_18903)
);

INVx1_ASAP7_75t_L g18904 ( 
.A(n_18731),
.Y(n_18904)
);

INVx1_ASAP7_75t_L g18905 ( 
.A(n_18765),
.Y(n_18905)
);

INVx2_ASAP7_75t_L g18906 ( 
.A(n_18757),
.Y(n_18906)
);

INVx1_ASAP7_75t_L g18907 ( 
.A(n_18721),
.Y(n_18907)
);

NAND2xp5_ASAP7_75t_L g18908 ( 
.A(n_18772),
.B(n_3096),
.Y(n_18908)
);

INVx1_ASAP7_75t_L g18909 ( 
.A(n_18826),
.Y(n_18909)
);

INVx1_ASAP7_75t_L g18910 ( 
.A(n_18798),
.Y(n_18910)
);

OR2x2_ASAP7_75t_L g18911 ( 
.A(n_18776),
.B(n_3097),
.Y(n_18911)
);

NAND2xp5_ASAP7_75t_L g18912 ( 
.A(n_18747),
.B(n_3098),
.Y(n_18912)
);

HB1xp67_ASAP7_75t_L g18913 ( 
.A(n_18754),
.Y(n_18913)
);

AND2x2_ASAP7_75t_L g18914 ( 
.A(n_18815),
.B(n_3098),
.Y(n_18914)
);

AOI22xp5_ASAP7_75t_L g18915 ( 
.A1(n_18817),
.A2(n_3101),
.B1(n_3099),
.B2(n_3100),
.Y(n_18915)
);

NAND2xp5_ASAP7_75t_L g18916 ( 
.A(n_18750),
.B(n_3099),
.Y(n_18916)
);

INVx2_ASAP7_75t_L g18917 ( 
.A(n_18760),
.Y(n_18917)
);

INVx1_ASAP7_75t_L g18918 ( 
.A(n_18819),
.Y(n_18918)
);

AND2x2_ASAP7_75t_L g18919 ( 
.A(n_18823),
.B(n_3100),
.Y(n_18919)
);

INVx1_ASAP7_75t_L g18920 ( 
.A(n_18749),
.Y(n_18920)
);

INVx1_ASAP7_75t_L g18921 ( 
.A(n_18733),
.Y(n_18921)
);

INVx1_ASAP7_75t_L g18922 ( 
.A(n_18767),
.Y(n_18922)
);

INVx1_ASAP7_75t_L g18923 ( 
.A(n_18794),
.Y(n_18923)
);

NAND2x1_ASAP7_75t_L g18924 ( 
.A(n_18816),
.B(n_18824),
.Y(n_18924)
);

NOR2x1_ASAP7_75t_L g18925 ( 
.A(n_18810),
.B(n_3101),
.Y(n_18925)
);

INVx1_ASAP7_75t_L g18926 ( 
.A(n_18717),
.Y(n_18926)
);

INVx2_ASAP7_75t_L g18927 ( 
.A(n_18827),
.Y(n_18927)
);

INVx2_ASAP7_75t_L g18928 ( 
.A(n_18803),
.Y(n_18928)
);

AND2x2_ASAP7_75t_L g18929 ( 
.A(n_18753),
.B(n_3102),
.Y(n_18929)
);

NAND2xp5_ASAP7_75t_L g18930 ( 
.A(n_18780),
.B(n_3102),
.Y(n_18930)
);

INVx1_ASAP7_75t_L g18931 ( 
.A(n_18773),
.Y(n_18931)
);

HB1xp67_ASAP7_75t_L g18932 ( 
.A(n_18809),
.Y(n_18932)
);

INVx1_ASAP7_75t_L g18933 ( 
.A(n_18832),
.Y(n_18933)
);

INVx1_ASAP7_75t_L g18934 ( 
.A(n_18732),
.Y(n_18934)
);

HB1xp67_ASAP7_75t_L g18935 ( 
.A(n_18763),
.Y(n_18935)
);

NAND2xp5_ASAP7_75t_L g18936 ( 
.A(n_18795),
.B(n_3103),
.Y(n_18936)
);

NOR2xp33_ASAP7_75t_L g18937 ( 
.A(n_18758),
.B(n_3103),
.Y(n_18937)
);

HB1xp67_ASAP7_75t_L g18938 ( 
.A(n_18758),
.Y(n_18938)
);

NAND2xp5_ASAP7_75t_L g18939 ( 
.A(n_18758),
.B(n_3104),
.Y(n_18939)
);

INVx1_ASAP7_75t_L g18940 ( 
.A(n_18758),
.Y(n_18940)
);

AND2x2_ASAP7_75t_L g18941 ( 
.A(n_18771),
.B(n_3105),
.Y(n_18941)
);

AND2x2_ASAP7_75t_L g18942 ( 
.A(n_18771),
.B(n_3105),
.Y(n_18942)
);

INVx1_ASAP7_75t_L g18943 ( 
.A(n_18758),
.Y(n_18943)
);

NAND2xp5_ASAP7_75t_L g18944 ( 
.A(n_18758),
.B(n_3106),
.Y(n_18944)
);

HB1xp67_ASAP7_75t_L g18945 ( 
.A(n_18758),
.Y(n_18945)
);

INVxp67_ASAP7_75t_L g18946 ( 
.A(n_18758),
.Y(n_18946)
);

INVx1_ASAP7_75t_L g18947 ( 
.A(n_18758),
.Y(n_18947)
);

INVx1_ASAP7_75t_L g18948 ( 
.A(n_18758),
.Y(n_18948)
);

INVx1_ASAP7_75t_L g18949 ( 
.A(n_18758),
.Y(n_18949)
);

NOR2xp33_ASAP7_75t_L g18950 ( 
.A(n_18758),
.B(n_3107),
.Y(n_18950)
);

NAND2xp5_ASAP7_75t_L g18951 ( 
.A(n_18758),
.B(n_3107),
.Y(n_18951)
);

INVx2_ASAP7_75t_SL g18952 ( 
.A(n_18758),
.Y(n_18952)
);

AND2x2_ASAP7_75t_L g18953 ( 
.A(n_18771),
.B(n_3108),
.Y(n_18953)
);

AND2x2_ASAP7_75t_L g18954 ( 
.A(n_18771),
.B(n_3108),
.Y(n_18954)
);

NAND2xp5_ASAP7_75t_L g18955 ( 
.A(n_18758),
.B(n_3110),
.Y(n_18955)
);

AND2x2_ASAP7_75t_L g18956 ( 
.A(n_18771),
.B(n_3110),
.Y(n_18956)
);

INVx1_ASAP7_75t_L g18957 ( 
.A(n_18758),
.Y(n_18957)
);

AOI222xp33_ASAP7_75t_L g18958 ( 
.A1(n_18724),
.A2(n_3114),
.B1(n_3116),
.B2(n_3111),
.C1(n_3112),
.C2(n_3115),
.Y(n_18958)
);

OR2x2_ASAP7_75t_L g18959 ( 
.A(n_18758),
.B(n_3111),
.Y(n_18959)
);

NAND2xp5_ASAP7_75t_L g18960 ( 
.A(n_18758),
.B(n_3112),
.Y(n_18960)
);

NOR2xp33_ASAP7_75t_SL g18961 ( 
.A(n_18801),
.B(n_3115),
.Y(n_18961)
);

INVx2_ASAP7_75t_L g18962 ( 
.A(n_18758),
.Y(n_18962)
);

AND2x2_ASAP7_75t_L g18963 ( 
.A(n_18771),
.B(n_3116),
.Y(n_18963)
);

INVx1_ASAP7_75t_L g18964 ( 
.A(n_18758),
.Y(n_18964)
);

INVx1_ASAP7_75t_L g18965 ( 
.A(n_18758),
.Y(n_18965)
);

NAND2xp5_ASAP7_75t_L g18966 ( 
.A(n_18758),
.B(n_3117),
.Y(n_18966)
);

NAND2xp5_ASAP7_75t_L g18967 ( 
.A(n_18758),
.B(n_3117),
.Y(n_18967)
);

OAI22xp5_ASAP7_75t_L g18968 ( 
.A1(n_18764),
.A2(n_3120),
.B1(n_3118),
.B2(n_3119),
.Y(n_18968)
);

INVx2_ASAP7_75t_L g18969 ( 
.A(n_18758),
.Y(n_18969)
);

OAI21xp33_ASAP7_75t_L g18970 ( 
.A1(n_18764),
.A2(n_3118),
.B(n_3119),
.Y(n_18970)
);

AND2x2_ASAP7_75t_L g18971 ( 
.A(n_18771),
.B(n_3120),
.Y(n_18971)
);

O2A1O1Ixp33_ASAP7_75t_L g18972 ( 
.A1(n_18938),
.A2(n_18945),
.B(n_18946),
.C(n_18952),
.Y(n_18972)
);

NAND2xp5_ASAP7_75t_SL g18973 ( 
.A(n_18962),
.B(n_3121),
.Y(n_18973)
);

NAND2x1_ASAP7_75t_SL g18974 ( 
.A(n_18853),
.B(n_3121),
.Y(n_18974)
);

AND2x2_ASAP7_75t_L g18975 ( 
.A(n_18969),
.B(n_3122),
.Y(n_18975)
);

INVx2_ASAP7_75t_L g18976 ( 
.A(n_18959),
.Y(n_18976)
);

OR2x2_ASAP7_75t_L g18977 ( 
.A(n_18841),
.B(n_3122),
.Y(n_18977)
);

OAI21xp33_ASAP7_75t_L g18978 ( 
.A1(n_18910),
.A2(n_3123),
.B(n_3124),
.Y(n_18978)
);

NOR2xp33_ASAP7_75t_L g18979 ( 
.A(n_18970),
.B(n_3123),
.Y(n_18979)
);

INVx1_ASAP7_75t_L g18980 ( 
.A(n_18919),
.Y(n_18980)
);

OAI21xp5_ASAP7_75t_L g18981 ( 
.A1(n_18837),
.A2(n_3124),
.B(n_3125),
.Y(n_18981)
);

O2A1O1Ixp33_ASAP7_75t_L g18982 ( 
.A1(n_18939),
.A2(n_3127),
.B(n_3125),
.C(n_3126),
.Y(n_18982)
);

O2A1O1Ixp33_ASAP7_75t_L g18983 ( 
.A1(n_18944),
.A2(n_18955),
.B(n_18960),
.C(n_18951),
.Y(n_18983)
);

NAND2xp5_ASAP7_75t_L g18984 ( 
.A(n_18849),
.B(n_3126),
.Y(n_18984)
);

BUFx3_ASAP7_75t_L g18985 ( 
.A(n_18839),
.Y(n_18985)
);

NOR2xp67_ASAP7_75t_L g18986 ( 
.A(n_18842),
.B(n_18890),
.Y(n_18986)
);

AND2x2_ASAP7_75t_L g18987 ( 
.A(n_18845),
.B(n_3127),
.Y(n_18987)
);

INVx1_ASAP7_75t_L g18988 ( 
.A(n_18966),
.Y(n_18988)
);

INVxp67_ASAP7_75t_SL g18989 ( 
.A(n_18937),
.Y(n_18989)
);

NAND2xp5_ASAP7_75t_L g18990 ( 
.A(n_18914),
.B(n_3128),
.Y(n_18990)
);

INVx1_ASAP7_75t_L g18991 ( 
.A(n_18967),
.Y(n_18991)
);

AOI22xp5_ASAP7_75t_L g18992 ( 
.A1(n_18834),
.A2(n_18900),
.B1(n_18943),
.B2(n_18940),
.Y(n_18992)
);

INVx1_ASAP7_75t_SL g18993 ( 
.A(n_18855),
.Y(n_18993)
);

NAND2xp5_ASAP7_75t_L g18994 ( 
.A(n_18950),
.B(n_3128),
.Y(n_18994)
);

OAI222xp33_ASAP7_75t_L g18995 ( 
.A1(n_18947),
.A2(n_3131),
.B1(n_3133),
.B2(n_3129),
.C1(n_3130),
.C2(n_3132),
.Y(n_18995)
);

INVx2_ASAP7_75t_L g18996 ( 
.A(n_18862),
.Y(n_18996)
);

OR2x2_ASAP7_75t_L g18997 ( 
.A(n_18872),
.B(n_3129),
.Y(n_18997)
);

AOI21xp5_ASAP7_75t_L g18998 ( 
.A1(n_18948),
.A2(n_18957),
.B(n_18949),
.Y(n_18998)
);

AOI22xp33_ASAP7_75t_SL g18999 ( 
.A1(n_18964),
.A2(n_3133),
.B1(n_3130),
.B2(n_3131),
.Y(n_18999)
);

INVx1_ASAP7_75t_L g19000 ( 
.A(n_18846),
.Y(n_19000)
);

OR2x2_ASAP7_75t_L g19001 ( 
.A(n_18844),
.B(n_3134),
.Y(n_19001)
);

O2A1O1Ixp33_ASAP7_75t_L g19002 ( 
.A1(n_18965),
.A2(n_18867),
.B(n_18936),
.C(n_18860),
.Y(n_19002)
);

OAI21xp33_ASAP7_75t_L g19003 ( 
.A1(n_18889),
.A2(n_3134),
.B(n_3135),
.Y(n_19003)
);

AOI222xp33_ASAP7_75t_L g19004 ( 
.A1(n_18859),
.A2(n_3137),
.B1(n_3139),
.B2(n_3135),
.C1(n_3136),
.C2(n_3138),
.Y(n_19004)
);

INVx1_ASAP7_75t_L g19005 ( 
.A(n_18857),
.Y(n_19005)
);

INVx1_ASAP7_75t_L g19006 ( 
.A(n_18877),
.Y(n_19006)
);

OAI21xp33_ASAP7_75t_L g19007 ( 
.A1(n_18854),
.A2(n_3136),
.B(n_3140),
.Y(n_19007)
);

NOR4xp25_ASAP7_75t_L g19008 ( 
.A(n_18858),
.B(n_3142),
.C(n_3140),
.D(n_3141),
.Y(n_19008)
);

INVx2_ASAP7_75t_L g19009 ( 
.A(n_18911),
.Y(n_19009)
);

INVx1_ASAP7_75t_L g19010 ( 
.A(n_18856),
.Y(n_19010)
);

NAND2xp5_ASAP7_75t_L g19011 ( 
.A(n_18958),
.B(n_3141),
.Y(n_19011)
);

INVx1_ASAP7_75t_L g19012 ( 
.A(n_18882),
.Y(n_19012)
);

INVx2_ASAP7_75t_SL g19013 ( 
.A(n_18836),
.Y(n_19013)
);

NAND2xp5_ASAP7_75t_L g19014 ( 
.A(n_18869),
.B(n_3142),
.Y(n_19014)
);

INVx1_ASAP7_75t_L g19015 ( 
.A(n_18941),
.Y(n_19015)
);

INVx1_ASAP7_75t_L g19016 ( 
.A(n_18942),
.Y(n_19016)
);

NAND2xp5_ASAP7_75t_SL g19017 ( 
.A(n_18890),
.B(n_3143),
.Y(n_19017)
);

AOI211xp5_ASAP7_75t_L g19018 ( 
.A1(n_18835),
.A2(n_3147),
.B(n_3145),
.C(n_3146),
.Y(n_19018)
);

INVx2_ASAP7_75t_SL g19019 ( 
.A(n_18953),
.Y(n_19019)
);

XOR2xp5_ASAP7_75t_L g19020 ( 
.A(n_18932),
.B(n_3145),
.Y(n_19020)
);

INVxp67_ASAP7_75t_L g19021 ( 
.A(n_18954),
.Y(n_19021)
);

OAI21xp33_ASAP7_75t_SL g19022 ( 
.A1(n_18850),
.A2(n_3146),
.B(n_3147),
.Y(n_19022)
);

AND2x2_ASAP7_75t_L g19023 ( 
.A(n_18897),
.B(n_3148),
.Y(n_19023)
);

NAND2xp5_ASAP7_75t_L g19024 ( 
.A(n_18956),
.B(n_3148),
.Y(n_19024)
);

AOI221x1_ASAP7_75t_L g19025 ( 
.A1(n_18931),
.A2(n_3151),
.B1(n_3149),
.B2(n_3150),
.C(n_3152),
.Y(n_19025)
);

OR2x2_ASAP7_75t_L g19026 ( 
.A(n_18880),
.B(n_3149),
.Y(n_19026)
);

NOR3xp33_ASAP7_75t_L g19027 ( 
.A(n_18896),
.B(n_3150),
.C(n_3151),
.Y(n_19027)
);

AOI322xp5_ASAP7_75t_L g19028 ( 
.A1(n_18847),
.A2(n_3157),
.A3(n_3156),
.B1(n_3154),
.B2(n_3152),
.C1(n_3153),
.C2(n_3155),
.Y(n_19028)
);

INVx1_ASAP7_75t_L g19029 ( 
.A(n_18963),
.Y(n_19029)
);

OR2x2_ASAP7_75t_L g19030 ( 
.A(n_18891),
.B(n_3153),
.Y(n_19030)
);

AOI211xp5_ASAP7_75t_L g19031 ( 
.A1(n_18852),
.A2(n_18863),
.B(n_18968),
.C(n_18838),
.Y(n_19031)
);

INVx1_ASAP7_75t_L g19032 ( 
.A(n_18971),
.Y(n_19032)
);

NAND2xp5_ASAP7_75t_L g19033 ( 
.A(n_18883),
.B(n_3154),
.Y(n_19033)
);

INVx1_ASAP7_75t_L g19034 ( 
.A(n_18885),
.Y(n_19034)
);

NAND2xp5_ASAP7_75t_L g19035 ( 
.A(n_18894),
.B(n_3155),
.Y(n_19035)
);

INVx1_ASAP7_75t_L g19036 ( 
.A(n_18881),
.Y(n_19036)
);

XNOR2xp5_ASAP7_75t_L g19037 ( 
.A(n_18928),
.B(n_3156),
.Y(n_19037)
);

NAND2xp5_ASAP7_75t_L g19038 ( 
.A(n_18898),
.B(n_3158),
.Y(n_19038)
);

AOI222xp33_ASAP7_75t_L g19039 ( 
.A1(n_18843),
.A2(n_3160),
.B1(n_3162),
.B2(n_3158),
.C1(n_3159),
.C2(n_3161),
.Y(n_19039)
);

INVx1_ASAP7_75t_L g19040 ( 
.A(n_18888),
.Y(n_19040)
);

AOI21xp5_ASAP7_75t_L g19041 ( 
.A1(n_18893),
.A2(n_3160),
.B(n_3162),
.Y(n_19041)
);

AOI22xp5_ASAP7_75t_L g19042 ( 
.A1(n_18961),
.A2(n_3165),
.B1(n_3163),
.B2(n_3164),
.Y(n_19042)
);

OR2x2_ASAP7_75t_L g19043 ( 
.A(n_18884),
.B(n_3164),
.Y(n_19043)
);

AOI22x1_ASAP7_75t_L g19044 ( 
.A1(n_18887),
.A2(n_3167),
.B1(n_3165),
.B2(n_3166),
.Y(n_19044)
);

NAND2xp5_ASAP7_75t_L g19045 ( 
.A(n_18840),
.B(n_3166),
.Y(n_19045)
);

INVx1_ASAP7_75t_SL g19046 ( 
.A(n_18861),
.Y(n_19046)
);

AOI22xp33_ASAP7_75t_L g19047 ( 
.A1(n_18864),
.A2(n_3169),
.B1(n_3167),
.B2(n_3168),
.Y(n_19047)
);

INVx1_ASAP7_75t_SL g19048 ( 
.A(n_18929),
.Y(n_19048)
);

OAI21xp33_ASAP7_75t_L g19049 ( 
.A1(n_18934),
.A2(n_3168),
.B(n_3169),
.Y(n_19049)
);

NAND2xp5_ASAP7_75t_L g19050 ( 
.A(n_18848),
.B(n_3170),
.Y(n_19050)
);

NAND2xp5_ASAP7_75t_SL g19051 ( 
.A(n_18906),
.B(n_3171),
.Y(n_19051)
);

NAND2xp5_ASAP7_75t_L g19052 ( 
.A(n_18851),
.B(n_3171),
.Y(n_19052)
);

INVx2_ASAP7_75t_SL g19053 ( 
.A(n_18886),
.Y(n_19053)
);

AOI21xp5_ASAP7_75t_L g19054 ( 
.A1(n_18930),
.A2(n_3172),
.B(n_3173),
.Y(n_19054)
);

O2A1O1Ixp33_ASAP7_75t_L g19055 ( 
.A1(n_18899),
.A2(n_3174),
.B(n_3172),
.C(n_3173),
.Y(n_19055)
);

AOI21xp33_ASAP7_75t_SL g19056 ( 
.A1(n_18873),
.A2(n_3174),
.B(n_3175),
.Y(n_19056)
);

NOR2xp67_ASAP7_75t_L g19057 ( 
.A(n_18903),
.B(n_3175),
.Y(n_19057)
);

INVx1_ASAP7_75t_L g19058 ( 
.A(n_18912),
.Y(n_19058)
);

INVxp67_ASAP7_75t_L g19059 ( 
.A(n_18913),
.Y(n_19059)
);

NAND2xp5_ASAP7_75t_L g19060 ( 
.A(n_18915),
.B(n_3176),
.Y(n_19060)
);

INVx1_ASAP7_75t_L g19061 ( 
.A(n_18876),
.Y(n_19061)
);

NAND2xp5_ASAP7_75t_L g19062 ( 
.A(n_18933),
.B(n_18866),
.Y(n_19062)
);

AOI211xp5_ASAP7_75t_L g19063 ( 
.A1(n_18892),
.A2(n_18920),
.B(n_18905),
.C(n_18874),
.Y(n_19063)
);

INVx1_ASAP7_75t_L g19064 ( 
.A(n_18908),
.Y(n_19064)
);

INVx1_ASAP7_75t_L g19065 ( 
.A(n_18925),
.Y(n_19065)
);

AND2x2_ASAP7_75t_L g19066 ( 
.A(n_18865),
.B(n_18927),
.Y(n_19066)
);

INVx1_ASAP7_75t_L g19067 ( 
.A(n_18916),
.Y(n_19067)
);

INVx1_ASAP7_75t_L g19068 ( 
.A(n_18924),
.Y(n_19068)
);

INVx1_ASAP7_75t_SL g19069 ( 
.A(n_18870),
.Y(n_19069)
);

NOR2xp33_ASAP7_75t_L g19070 ( 
.A(n_18926),
.B(n_3176),
.Y(n_19070)
);

INVx1_ASAP7_75t_L g19071 ( 
.A(n_18935),
.Y(n_19071)
);

AOI221xp5_ASAP7_75t_L g19072 ( 
.A1(n_18904),
.A2(n_3179),
.B1(n_3177),
.B2(n_3178),
.C(n_3180),
.Y(n_19072)
);

O2A1O1Ixp33_ASAP7_75t_L g19073 ( 
.A1(n_18917),
.A2(n_3179),
.B(n_3177),
.C(n_3178),
.Y(n_19073)
);

AOI222xp33_ASAP7_75t_L g19074 ( 
.A1(n_18907),
.A2(n_3183),
.B1(n_3185),
.B2(n_3181),
.C1(n_3182),
.C2(n_3184),
.Y(n_19074)
);

INVx1_ASAP7_75t_L g19075 ( 
.A(n_18909),
.Y(n_19075)
);

NAND2xp5_ASAP7_75t_L g19076 ( 
.A(n_18878),
.B(n_3181),
.Y(n_19076)
);

INVx1_ASAP7_75t_L g19077 ( 
.A(n_18921),
.Y(n_19077)
);

INVx1_ASAP7_75t_L g19078 ( 
.A(n_18922),
.Y(n_19078)
);

INVx1_ASAP7_75t_L g19079 ( 
.A(n_18923),
.Y(n_19079)
);

AOI222xp33_ASAP7_75t_L g19080 ( 
.A1(n_18918),
.A2(n_3184),
.B1(n_3186),
.B2(n_3182),
.C1(n_3183),
.C2(n_3185),
.Y(n_19080)
);

O2A1O1Ixp33_ASAP7_75t_L g19081 ( 
.A1(n_18902),
.A2(n_18871),
.B(n_18868),
.C(n_18875),
.Y(n_19081)
);

OAI22xp5_ASAP7_75t_L g19082 ( 
.A1(n_18895),
.A2(n_3188),
.B1(n_3186),
.B2(n_3187),
.Y(n_19082)
);

INVx1_ASAP7_75t_L g19083 ( 
.A(n_18901),
.Y(n_19083)
);

INVx1_ASAP7_75t_L g19084 ( 
.A(n_18879),
.Y(n_19084)
);

NAND3xp33_ASAP7_75t_L g19085 ( 
.A(n_18958),
.B(n_3188),
.C(n_3189),
.Y(n_19085)
);

INVx1_ASAP7_75t_L g19086 ( 
.A(n_18959),
.Y(n_19086)
);

NOR2xp33_ASAP7_75t_SL g19087 ( 
.A(n_18938),
.B(n_3189),
.Y(n_19087)
);

INVx1_ASAP7_75t_L g19088 ( 
.A(n_18959),
.Y(n_19088)
);

NOR2xp33_ASAP7_75t_L g19089 ( 
.A(n_18970),
.B(n_3190),
.Y(n_19089)
);

NAND2x1_ASAP7_75t_L g19090 ( 
.A(n_18853),
.B(n_3190),
.Y(n_19090)
);

AOI22xp5_ASAP7_75t_L g19091 ( 
.A1(n_18952),
.A2(n_3193),
.B1(n_3191),
.B2(n_3192),
.Y(n_19091)
);

OAI211xp5_ASAP7_75t_L g19092 ( 
.A1(n_18958),
.A2(n_3193),
.B(n_3191),
.C(n_3192),
.Y(n_19092)
);

AOI22xp33_ASAP7_75t_L g19093 ( 
.A1(n_18952),
.A2(n_3196),
.B1(n_3194),
.B2(n_3195),
.Y(n_19093)
);

NAND2xp5_ASAP7_75t_SL g19094 ( 
.A(n_18952),
.B(n_3194),
.Y(n_19094)
);

INVxp67_ASAP7_75t_L g19095 ( 
.A(n_18937),
.Y(n_19095)
);

INVx1_ASAP7_75t_L g19096 ( 
.A(n_18959),
.Y(n_19096)
);

XNOR2x1_ASAP7_75t_L g19097 ( 
.A(n_18834),
.B(n_3195),
.Y(n_19097)
);

NAND2xp5_ASAP7_75t_L g19098 ( 
.A(n_18849),
.B(n_3196),
.Y(n_19098)
);

NAND2xp5_ASAP7_75t_SL g19099 ( 
.A(n_18952),
.B(n_3197),
.Y(n_19099)
);

AND2x2_ASAP7_75t_L g19100 ( 
.A(n_18962),
.B(n_3197),
.Y(n_19100)
);

NAND2xp5_ASAP7_75t_L g19101 ( 
.A(n_18849),
.B(n_3198),
.Y(n_19101)
);

INVx2_ASAP7_75t_L g19102 ( 
.A(n_18959),
.Y(n_19102)
);

INVx1_ASAP7_75t_L g19103 ( 
.A(n_18959),
.Y(n_19103)
);

AND2x2_ASAP7_75t_L g19104 ( 
.A(n_18962),
.B(n_3198),
.Y(n_19104)
);

OAI211xp5_ASAP7_75t_L g19105 ( 
.A1(n_18958),
.A2(n_3201),
.B(n_3199),
.C(n_3200),
.Y(n_19105)
);

AOI211x1_ASAP7_75t_L g19106 ( 
.A1(n_18867),
.A2(n_3201),
.B(n_3199),
.C(n_3200),
.Y(n_19106)
);

INVx1_ASAP7_75t_L g19107 ( 
.A(n_18959),
.Y(n_19107)
);

INVx2_ASAP7_75t_SL g19108 ( 
.A(n_18959),
.Y(n_19108)
);

INVx1_ASAP7_75t_SL g19109 ( 
.A(n_18855),
.Y(n_19109)
);

OR2x2_ASAP7_75t_L g19110 ( 
.A(n_18841),
.B(n_3203),
.Y(n_19110)
);

INVxp67_ASAP7_75t_L g19111 ( 
.A(n_18937),
.Y(n_19111)
);

AOI21xp5_ASAP7_75t_L g19112 ( 
.A1(n_18938),
.A2(n_3203),
.B(n_3204),
.Y(n_19112)
);

AOI21xp5_ASAP7_75t_L g19113 ( 
.A1(n_18938),
.A2(n_3204),
.B(n_3205),
.Y(n_19113)
);

OAI21xp33_ASAP7_75t_SL g19114 ( 
.A1(n_18889),
.A2(n_3205),
.B(n_3206),
.Y(n_19114)
);

AOI322xp5_ASAP7_75t_L g19115 ( 
.A1(n_18845),
.A2(n_3211),
.A3(n_3210),
.B1(n_3208),
.B2(n_3206),
.C1(n_3207),
.C2(n_3209),
.Y(n_19115)
);

INVx1_ASAP7_75t_L g19116 ( 
.A(n_18959),
.Y(n_19116)
);

OAI21xp5_ASAP7_75t_L g19117 ( 
.A1(n_18998),
.A2(n_19059),
.B(n_18972),
.Y(n_19117)
);

INVx1_ASAP7_75t_L g19118 ( 
.A(n_18974),
.Y(n_19118)
);

AOI33xp33_ASAP7_75t_L g19119 ( 
.A1(n_18993),
.A2(n_3209),
.A3(n_3211),
.B1(n_3207),
.B2(n_3208),
.B3(n_3210),
.Y(n_19119)
);

AOI221xp5_ASAP7_75t_L g19120 ( 
.A1(n_19008),
.A2(n_3214),
.B1(n_3212),
.B2(n_3213),
.C(n_3215),
.Y(n_19120)
);

NAND2xp5_ASAP7_75t_L g19121 ( 
.A(n_18987),
.B(n_3212),
.Y(n_19121)
);

INVx2_ASAP7_75t_SL g19122 ( 
.A(n_19090),
.Y(n_19122)
);

INVx1_ASAP7_75t_L g19123 ( 
.A(n_19020),
.Y(n_19123)
);

OAI211xp5_ASAP7_75t_L g19124 ( 
.A1(n_19114),
.A2(n_3216),
.B(n_3213),
.C(n_3214),
.Y(n_19124)
);

NAND2xp5_ASAP7_75t_SL g19125 ( 
.A(n_19004),
.B(n_3216),
.Y(n_19125)
);

OAI21xp33_ASAP7_75t_SL g19126 ( 
.A1(n_19042),
.A2(n_3217),
.B(n_3218),
.Y(n_19126)
);

OAI21xp5_ASAP7_75t_SL g19127 ( 
.A1(n_19109),
.A2(n_3217),
.B(n_3218),
.Y(n_19127)
);

OAI21xp5_ASAP7_75t_L g19128 ( 
.A1(n_19085),
.A2(n_3219),
.B(n_3220),
.Y(n_19128)
);

OAI211xp5_ASAP7_75t_L g19129 ( 
.A1(n_19003),
.A2(n_3221),
.B(n_3219),
.C(n_3220),
.Y(n_19129)
);

OAI222xp33_ASAP7_75t_L g19130 ( 
.A1(n_18992),
.A2(n_3223),
.B1(n_3225),
.B2(n_3221),
.C1(n_3222),
.C2(n_3224),
.Y(n_19130)
);

O2A1O1Ixp33_ASAP7_75t_SL g19131 ( 
.A1(n_19014),
.A2(n_3225),
.B(n_3222),
.C(n_3223),
.Y(n_19131)
);

A2O1A1Ixp33_ASAP7_75t_L g19132 ( 
.A1(n_19073),
.A2(n_3228),
.B(n_3226),
.C(n_3227),
.Y(n_19132)
);

OAI211xp5_ASAP7_75t_L g19133 ( 
.A1(n_19022),
.A2(n_3230),
.B(n_3227),
.C(n_3229),
.Y(n_19133)
);

AOI211xp5_ASAP7_75t_SL g19134 ( 
.A1(n_18986),
.A2(n_19045),
.B(n_19078),
.C(n_19071),
.Y(n_19134)
);

OAI211xp5_ASAP7_75t_L g19135 ( 
.A1(n_19056),
.A2(n_3232),
.B(n_3230),
.C(n_3231),
.Y(n_19135)
);

OR2x2_ASAP7_75t_L g19136 ( 
.A(n_19033),
.B(n_3231),
.Y(n_19136)
);

AO22x2_ASAP7_75t_L g19137 ( 
.A1(n_19097),
.A2(n_3234),
.B1(n_3232),
.B2(n_3233),
.Y(n_19137)
);

AOI221xp5_ASAP7_75t_L g19138 ( 
.A1(n_19106),
.A2(n_3236),
.B1(n_3233),
.B2(n_3235),
.C(n_3237),
.Y(n_19138)
);

AOI22xp5_ASAP7_75t_L g19139 ( 
.A1(n_19079),
.A2(n_3238),
.B1(n_3235),
.B2(n_3237),
.Y(n_19139)
);

AOI221xp5_ASAP7_75t_L g19140 ( 
.A1(n_19092),
.A2(n_3240),
.B1(n_3238),
.B2(n_3239),
.C(n_3241),
.Y(n_19140)
);

AOI21xp5_ASAP7_75t_L g19141 ( 
.A1(n_19062),
.A2(n_3239),
.B(n_3240),
.Y(n_19141)
);

O2A1O1Ixp33_ASAP7_75t_L g19142 ( 
.A1(n_19051),
.A2(n_18990),
.B(n_19035),
.C(n_19012),
.Y(n_19142)
);

OAI21xp5_ASAP7_75t_SL g19143 ( 
.A1(n_19105),
.A2(n_3241),
.B(n_3242),
.Y(n_19143)
);

NOR2xp33_ASAP7_75t_SL g19144 ( 
.A(n_18995),
.B(n_3242),
.Y(n_19144)
);

AOI21xp5_ASAP7_75t_L g19145 ( 
.A1(n_19011),
.A2(n_3243),
.B(n_3244),
.Y(n_19145)
);

AOI22xp33_ASAP7_75t_L g19146 ( 
.A1(n_18985),
.A2(n_3246),
.B1(n_3244),
.B2(n_3245),
.Y(n_19146)
);

O2A1O1Ixp33_ASAP7_75t_L g19147 ( 
.A1(n_18984),
.A2(n_3247),
.B(n_3245),
.C(n_3246),
.Y(n_19147)
);

NAND2xp33_ASAP7_75t_SL g19148 ( 
.A(n_19026),
.B(n_3247),
.Y(n_19148)
);

AOI21xp5_ASAP7_75t_SL g19149 ( 
.A1(n_19025),
.A2(n_3248),
.B(n_3249),
.Y(n_19149)
);

OAI22xp5_ASAP7_75t_L g19150 ( 
.A1(n_19077),
.A2(n_3251),
.B1(n_3248),
.B2(n_3250),
.Y(n_19150)
);

AOI21xp5_ASAP7_75t_L g19151 ( 
.A1(n_19081),
.A2(n_3250),
.B(n_3251),
.Y(n_19151)
);

NOR4xp25_ASAP7_75t_L g19152 ( 
.A(n_19002),
.B(n_3255),
.C(n_3253),
.D(n_3254),
.Y(n_19152)
);

AOI211xp5_ASAP7_75t_SL g19153 ( 
.A1(n_19075),
.A2(n_3256),
.B(n_3254),
.C(n_3255),
.Y(n_19153)
);

INVx1_ASAP7_75t_SL g19154 ( 
.A(n_19023),
.Y(n_19154)
);

INVxp67_ASAP7_75t_SL g19155 ( 
.A(n_19037),
.Y(n_19155)
);

AOI21xp33_ASAP7_75t_L g19156 ( 
.A1(n_18997),
.A2(n_3256),
.B(n_3257),
.Y(n_19156)
);

OR2x2_ASAP7_75t_L g19157 ( 
.A(n_19098),
.B(n_3257),
.Y(n_19157)
);

AOI22xp5_ASAP7_75t_L g19158 ( 
.A1(n_19066),
.A2(n_3260),
.B1(n_3258),
.B2(n_3259),
.Y(n_19158)
);

AO22x2_ASAP7_75t_L g19159 ( 
.A1(n_19034),
.A2(n_3261),
.B1(n_3258),
.B2(n_3260),
.Y(n_19159)
);

NAND3xp33_ASAP7_75t_SL g19160 ( 
.A(n_19063),
.B(n_3262),
.C(n_3263),
.Y(n_19160)
);

AOI211x1_ASAP7_75t_SL g19161 ( 
.A1(n_19057),
.A2(n_3264),
.B(n_3262),
.C(n_3263),
.Y(n_19161)
);

OA21x2_ASAP7_75t_SL g19162 ( 
.A1(n_19046),
.A2(n_3264),
.B(n_3265),
.Y(n_19162)
);

OAI22xp33_ASAP7_75t_L g19163 ( 
.A1(n_19087),
.A2(n_3267),
.B1(n_3265),
.B2(n_3266),
.Y(n_19163)
);

INVx1_ASAP7_75t_L g19164 ( 
.A(n_18977),
.Y(n_19164)
);

AOI21xp5_ASAP7_75t_SL g19165 ( 
.A1(n_19017),
.A2(n_19055),
.B(n_18982),
.Y(n_19165)
);

OAI21xp33_ASAP7_75t_L g19166 ( 
.A1(n_19069),
.A2(n_3266),
.B(n_3267),
.Y(n_19166)
);

AOI222xp33_ASAP7_75t_L g19167 ( 
.A1(n_19068),
.A2(n_3270),
.B1(n_3272),
.B2(n_3268),
.C1(n_3269),
.C2(n_3271),
.Y(n_19167)
);

OAI22xp5_ASAP7_75t_L g19168 ( 
.A1(n_19101),
.A2(n_3270),
.B1(n_3268),
.B2(n_3269),
.Y(n_19168)
);

NAND3xp33_ASAP7_75t_L g19169 ( 
.A(n_19027),
.B(n_3272),
.C(n_3273),
.Y(n_19169)
);

OAI22xp5_ASAP7_75t_L g19170 ( 
.A1(n_19024),
.A2(n_3275),
.B1(n_3273),
.B2(n_3274),
.Y(n_19170)
);

INVx2_ASAP7_75t_L g19171 ( 
.A(n_18975),
.Y(n_19171)
);

OAI22xp33_ASAP7_75t_SL g19172 ( 
.A1(n_19030),
.A2(n_3277),
.B1(n_3274),
.B2(n_3276),
.Y(n_19172)
);

OAI21xp33_ASAP7_75t_L g19173 ( 
.A1(n_19083),
.A2(n_19089),
.B(n_18979),
.Y(n_19173)
);

O2A1O1Ixp5_ASAP7_75t_L g19174 ( 
.A1(n_19060),
.A2(n_19065),
.B(n_18996),
.C(n_19054),
.Y(n_19174)
);

OAI22xp33_ASAP7_75t_L g19175 ( 
.A1(n_19043),
.A2(n_3278),
.B1(n_3276),
.B2(n_3277),
.Y(n_19175)
);

OAI211xp5_ASAP7_75t_SL g19176 ( 
.A1(n_19031),
.A2(n_3280),
.B(n_3278),
.C(n_3279),
.Y(n_19176)
);

AOI211xp5_ASAP7_75t_L g19177 ( 
.A1(n_19041),
.A2(n_3281),
.B(n_3279),
.C(n_3280),
.Y(n_19177)
);

AOI21xp5_ASAP7_75t_L g19178 ( 
.A1(n_19038),
.A2(n_3281),
.B(n_3282),
.Y(n_19178)
);

NOR4xp25_ASAP7_75t_L g19179 ( 
.A(n_18983),
.B(n_3284),
.C(n_3282),
.D(n_3283),
.Y(n_19179)
);

NOR2xp33_ASAP7_75t_L g19180 ( 
.A(n_19049),
.B(n_3283),
.Y(n_19180)
);

AOI221xp5_ASAP7_75t_SL g19181 ( 
.A1(n_19021),
.A2(n_3286),
.B1(n_3284),
.B2(n_3285),
.C(n_3287),
.Y(n_19181)
);

OAI322xp33_ASAP7_75t_L g19182 ( 
.A1(n_19095),
.A2(n_3291),
.A3(n_3290),
.B1(n_3288),
.B2(n_3285),
.C1(n_3286),
.C2(n_3289),
.Y(n_19182)
);

NAND2xp5_ASAP7_75t_L g19183 ( 
.A(n_19028),
.B(n_3288),
.Y(n_19183)
);

OAI211xp5_ASAP7_75t_L g19184 ( 
.A1(n_19080),
.A2(n_3292),
.B(n_3289),
.C(n_3291),
.Y(n_19184)
);

OAI22xp5_ASAP7_75t_L g19185 ( 
.A1(n_18994),
.A2(n_3294),
.B1(n_3292),
.B2(n_3293),
.Y(n_19185)
);

OAI22xp33_ASAP7_75t_L g19186 ( 
.A1(n_19084),
.A2(n_19013),
.B1(n_19019),
.B2(n_18980),
.Y(n_19186)
);

NAND2x1p5_ASAP7_75t_L g19187 ( 
.A(n_19094),
.B(n_3293),
.Y(n_19187)
);

NOR2xp33_ASAP7_75t_L g19188 ( 
.A(n_19110),
.B(n_3294),
.Y(n_19188)
);

NOR2xp33_ASAP7_75t_L g19189 ( 
.A(n_19099),
.B(n_3295),
.Y(n_19189)
);

INVxp33_ASAP7_75t_L g19190 ( 
.A(n_19070),
.Y(n_19190)
);

OAI221xp5_ASAP7_75t_L g19191 ( 
.A1(n_19018),
.A2(n_3297),
.B1(n_3295),
.B2(n_3296),
.C(n_3298),
.Y(n_19191)
);

INVx1_ASAP7_75t_L g19192 ( 
.A(n_19001),
.Y(n_19192)
);

INVx1_ASAP7_75t_SL g19193 ( 
.A(n_19100),
.Y(n_19193)
);

AOI22xp5_ASAP7_75t_L g19194 ( 
.A1(n_19000),
.A2(n_3299),
.B1(n_3296),
.B2(n_3297),
.Y(n_19194)
);

INVx2_ASAP7_75t_SL g19195 ( 
.A(n_19104),
.Y(n_19195)
);

AOI21xp5_ASAP7_75t_L g19196 ( 
.A1(n_18989),
.A2(n_3299),
.B(n_3300),
.Y(n_19196)
);

OAI22x1_ASAP7_75t_SL g19197 ( 
.A1(n_19015),
.A2(n_3302),
.B1(n_3300),
.B2(n_3301),
.Y(n_19197)
);

INVx2_ASAP7_75t_SL g19198 ( 
.A(n_18973),
.Y(n_19198)
);

OAI22xp5_ASAP7_75t_L g19199 ( 
.A1(n_19111),
.A2(n_3303),
.B1(n_3301),
.B2(n_3302),
.Y(n_19199)
);

AOI222xp33_ASAP7_75t_SL g19200 ( 
.A1(n_19048),
.A2(n_3305),
.B1(n_3307),
.B2(n_3303),
.C1(n_3304),
.C2(n_3306),
.Y(n_19200)
);

AOI32xp33_ASAP7_75t_L g19201 ( 
.A1(n_19010),
.A2(n_3307),
.A3(n_3304),
.B1(n_3306),
.B2(n_3308),
.Y(n_19201)
);

AOI21xp33_ASAP7_75t_L g19202 ( 
.A1(n_19108),
.A2(n_3308),
.B(n_3309),
.Y(n_19202)
);

OAI21xp33_ASAP7_75t_L g19203 ( 
.A1(n_19016),
.A2(n_3309),
.B(n_3310),
.Y(n_19203)
);

OAI21xp5_ASAP7_75t_L g19204 ( 
.A1(n_19029),
.A2(n_3310),
.B(n_3311),
.Y(n_19204)
);

AOI322xp5_ASAP7_75t_L g19205 ( 
.A1(n_19053),
.A2(n_3316),
.A3(n_3315),
.B1(n_3313),
.B2(n_3311),
.C1(n_3312),
.C2(n_3314),
.Y(n_19205)
);

AOI211xp5_ASAP7_75t_L g19206 ( 
.A1(n_19112),
.A2(n_3314),
.B(n_3312),
.C(n_3313),
.Y(n_19206)
);

OAI21xp33_ASAP7_75t_L g19207 ( 
.A1(n_19032),
.A2(n_3315),
.B(n_3316),
.Y(n_19207)
);

OAI221xp5_ASAP7_75t_L g19208 ( 
.A1(n_19044),
.A2(n_3319),
.B1(n_3317),
.B2(n_3318),
.C(n_3320),
.Y(n_19208)
);

AOI211xp5_ASAP7_75t_L g19209 ( 
.A1(n_19113),
.A2(n_19007),
.B(n_19088),
.C(n_19086),
.Y(n_19209)
);

INVx1_ASAP7_75t_L g19210 ( 
.A(n_19052),
.Y(n_19210)
);

OAI211xp5_ASAP7_75t_SL g19211 ( 
.A1(n_19096),
.A2(n_3319),
.B(n_3317),
.C(n_3318),
.Y(n_19211)
);

OAI21xp5_ASAP7_75t_L g19212 ( 
.A1(n_19103),
.A2(n_3320),
.B(n_3321),
.Y(n_19212)
);

OAI221xp5_ASAP7_75t_L g19213 ( 
.A1(n_18978),
.A2(n_3323),
.B1(n_3321),
.B2(n_3322),
.C(n_3325),
.Y(n_19213)
);

NAND2xp5_ASAP7_75t_L g19214 ( 
.A(n_19050),
.B(n_3323),
.Y(n_19214)
);

OAI22xp33_ASAP7_75t_L g19215 ( 
.A1(n_19009),
.A2(n_3327),
.B1(n_3325),
.B2(n_3326),
.Y(n_19215)
);

AOI21xp33_ASAP7_75t_SL g19216 ( 
.A1(n_19074),
.A2(n_3326),
.B(n_3327),
.Y(n_19216)
);

AOI211xp5_ASAP7_75t_L g19217 ( 
.A1(n_19107),
.A2(n_19116),
.B(n_19058),
.C(n_19082),
.Y(n_19217)
);

AOI22xp5_ASAP7_75t_L g19218 ( 
.A1(n_18976),
.A2(n_3330),
.B1(n_3328),
.B2(n_3329),
.Y(n_19218)
);

OAI22xp5_ASAP7_75t_L g19219 ( 
.A1(n_19102),
.A2(n_3330),
.B1(n_3328),
.B2(n_3329),
.Y(n_19219)
);

O2A1O1Ixp33_ASAP7_75t_L g19220 ( 
.A1(n_18988),
.A2(n_3333),
.B(n_3331),
.C(n_3332),
.Y(n_19220)
);

AOI211xp5_ASAP7_75t_L g19221 ( 
.A1(n_18991),
.A2(n_19005),
.B(n_19006),
.C(n_18981),
.Y(n_19221)
);

OAI221xp5_ASAP7_75t_SL g19222 ( 
.A1(n_19061),
.A2(n_3333),
.B1(n_3331),
.B2(n_3332),
.C(n_3334),
.Y(n_19222)
);

OAI21xp5_ASAP7_75t_SL g19223 ( 
.A1(n_19064),
.A2(n_3334),
.B(n_3335),
.Y(n_19223)
);

INVx2_ASAP7_75t_SL g19224 ( 
.A(n_19076),
.Y(n_19224)
);

AOI221xp5_ASAP7_75t_L g19225 ( 
.A1(n_19067),
.A2(n_3337),
.B1(n_3335),
.B2(n_3336),
.C(n_3338),
.Y(n_19225)
);

INVxp67_ASAP7_75t_L g19226 ( 
.A(n_19039),
.Y(n_19226)
);

INVx1_ASAP7_75t_L g19227 ( 
.A(n_19036),
.Y(n_19227)
);

NAND3xp33_ASAP7_75t_L g19228 ( 
.A(n_19072),
.B(n_3336),
.C(n_3337),
.Y(n_19228)
);

AND2x2_ASAP7_75t_L g19229 ( 
.A(n_19040),
.B(n_3338),
.Y(n_19229)
);

AOI22xp5_ASAP7_75t_L g19230 ( 
.A1(n_18999),
.A2(n_19091),
.B1(n_19093),
.B2(n_19047),
.Y(n_19230)
);

OAI21xp5_ASAP7_75t_L g19231 ( 
.A1(n_19115),
.A2(n_3339),
.B(n_3340),
.Y(n_19231)
);

OAI22xp5_ASAP7_75t_L g19232 ( 
.A1(n_19020),
.A2(n_3342),
.B1(n_3340),
.B2(n_3341),
.Y(n_19232)
);

NAND3xp33_ASAP7_75t_L g19233 ( 
.A(n_19004),
.B(n_3341),
.C(n_3342),
.Y(n_19233)
);

OAI311xp33_ASAP7_75t_L g19234 ( 
.A1(n_18992),
.A2(n_3345),
.A3(n_3343),
.B1(n_3344),
.C1(n_3346),
.Y(n_19234)
);

INVx2_ASAP7_75t_L g19235 ( 
.A(n_19023),
.Y(n_19235)
);

O2A1O1Ixp33_ASAP7_75t_L g19236 ( 
.A1(n_19090),
.A2(n_3345),
.B(n_3343),
.C(n_3344),
.Y(n_19236)
);

AOI22xp5_ASAP7_75t_L g19237 ( 
.A1(n_18993),
.A2(n_3348),
.B1(n_3346),
.B2(n_3347),
.Y(n_19237)
);

OAI21xp33_ASAP7_75t_SL g19238 ( 
.A1(n_18974),
.A2(n_3347),
.B(n_3349),
.Y(n_19238)
);

AOI21xp5_ASAP7_75t_L g19239 ( 
.A1(n_18972),
.A2(n_3349),
.B(n_3350),
.Y(n_19239)
);

OAI22xp5_ASAP7_75t_L g19240 ( 
.A1(n_19020),
.A2(n_3352),
.B1(n_3350),
.B2(n_3351),
.Y(n_19240)
);

OAI22xp33_ASAP7_75t_L g19241 ( 
.A1(n_19042),
.A2(n_3353),
.B1(n_3351),
.B2(n_3352),
.Y(n_19241)
);

INVx1_ASAP7_75t_L g19242 ( 
.A(n_18974),
.Y(n_19242)
);

AOI322xp5_ASAP7_75t_L g19243 ( 
.A1(n_18993),
.A2(n_3358),
.A3(n_3357),
.B1(n_3355),
.B2(n_3353),
.C1(n_3354),
.C2(n_3356),
.Y(n_19243)
);

OAI221xp5_ASAP7_75t_L g19244 ( 
.A1(n_19003),
.A2(n_3357),
.B1(n_3354),
.B2(n_3356),
.C(n_3358),
.Y(n_19244)
);

OR2x2_ASAP7_75t_L g19245 ( 
.A(n_19152),
.B(n_3359),
.Y(n_19245)
);

NAND2xp33_ASAP7_75t_SL g19246 ( 
.A(n_19122),
.B(n_3359),
.Y(n_19246)
);

INVx1_ASAP7_75t_L g19247 ( 
.A(n_19121),
.Y(n_19247)
);

NAND2xp5_ASAP7_75t_L g19248 ( 
.A(n_19179),
.B(n_3360),
.Y(n_19248)
);

AND2x2_ASAP7_75t_L g19249 ( 
.A(n_19137),
.B(n_3360),
.Y(n_19249)
);

NOR2x1_ASAP7_75t_L g19250 ( 
.A(n_19149),
.B(n_3361),
.Y(n_19250)
);

INVx1_ASAP7_75t_L g19251 ( 
.A(n_19137),
.Y(n_19251)
);

INVx1_ASAP7_75t_SL g19252 ( 
.A(n_19197),
.Y(n_19252)
);

INVx2_ASAP7_75t_L g19253 ( 
.A(n_19159),
.Y(n_19253)
);

OR2x2_ASAP7_75t_L g19254 ( 
.A(n_19160),
.B(n_3361),
.Y(n_19254)
);

INVx1_ASAP7_75t_L g19255 ( 
.A(n_19131),
.Y(n_19255)
);

NAND2xp5_ASAP7_75t_SL g19256 ( 
.A(n_19117),
.B(n_3362),
.Y(n_19256)
);

INVx1_ASAP7_75t_L g19257 ( 
.A(n_19136),
.Y(n_19257)
);

NAND2xp5_ASAP7_75t_L g19258 ( 
.A(n_19188),
.B(n_3362),
.Y(n_19258)
);

NAND3x1_ASAP7_75t_L g19259 ( 
.A(n_19118),
.B(n_3363),
.C(n_3364),
.Y(n_19259)
);

INVx2_ASAP7_75t_L g19260 ( 
.A(n_19159),
.Y(n_19260)
);

INVxp67_ASAP7_75t_L g19261 ( 
.A(n_19157),
.Y(n_19261)
);

INVx1_ASAP7_75t_L g19262 ( 
.A(n_19187),
.Y(n_19262)
);

OAI22xp5_ASAP7_75t_L g19263 ( 
.A1(n_19226),
.A2(n_3365),
.B1(n_3363),
.B2(n_3364),
.Y(n_19263)
);

NAND3xp33_ASAP7_75t_L g19264 ( 
.A(n_19134),
.B(n_3366),
.C(n_3367),
.Y(n_19264)
);

NOR2xp33_ASAP7_75t_L g19265 ( 
.A(n_19238),
.B(n_3367),
.Y(n_19265)
);

NOR2xp33_ASAP7_75t_L g19266 ( 
.A(n_19133),
.B(n_3368),
.Y(n_19266)
);

NAND3xp33_ASAP7_75t_L g19267 ( 
.A(n_19239),
.B(n_3368),
.C(n_3369),
.Y(n_19267)
);

NAND2xp5_ASAP7_75t_L g19268 ( 
.A(n_19223),
.B(n_3369),
.Y(n_19268)
);

NOR2xp33_ASAP7_75t_L g19269 ( 
.A(n_19143),
.B(n_3370),
.Y(n_19269)
);

NAND3xp33_ASAP7_75t_L g19270 ( 
.A(n_19151),
.B(n_3370),
.C(n_3371),
.Y(n_19270)
);

NAND2xp5_ASAP7_75t_L g19271 ( 
.A(n_19166),
.B(n_3371),
.Y(n_19271)
);

NOR2xp33_ASAP7_75t_L g19272 ( 
.A(n_19126),
.B(n_3372),
.Y(n_19272)
);

INVx1_ASAP7_75t_SL g19273 ( 
.A(n_19229),
.Y(n_19273)
);

INVx1_ASAP7_75t_L g19274 ( 
.A(n_19214),
.Y(n_19274)
);

AOI221x1_ASAP7_75t_L g19275 ( 
.A1(n_19173),
.A2(n_3374),
.B1(n_3372),
.B2(n_3373),
.C(n_3375),
.Y(n_19275)
);

INVx1_ASAP7_75t_L g19276 ( 
.A(n_19124),
.Y(n_19276)
);

NAND2xp5_ASAP7_75t_L g19277 ( 
.A(n_19172),
.B(n_3374),
.Y(n_19277)
);

AND2x2_ASAP7_75t_L g19278 ( 
.A(n_19235),
.B(n_3375),
.Y(n_19278)
);

NAND2xp5_ASAP7_75t_L g19279 ( 
.A(n_19196),
.B(n_3376),
.Y(n_19279)
);

INVx1_ASAP7_75t_L g19280 ( 
.A(n_19183),
.Y(n_19280)
);

NAND2xp5_ASAP7_75t_L g19281 ( 
.A(n_19203),
.B(n_3376),
.Y(n_19281)
);

INVx1_ASAP7_75t_SL g19282 ( 
.A(n_19148),
.Y(n_19282)
);

INVx1_ASAP7_75t_L g19283 ( 
.A(n_19135),
.Y(n_19283)
);

INVx2_ASAP7_75t_L g19284 ( 
.A(n_19171),
.Y(n_19284)
);

INVxp67_ASAP7_75t_SL g19285 ( 
.A(n_19236),
.Y(n_19285)
);

AND2x2_ASAP7_75t_L g19286 ( 
.A(n_19154),
.B(n_3377),
.Y(n_19286)
);

NAND2xp33_ASAP7_75t_L g19287 ( 
.A(n_19201),
.B(n_3377),
.Y(n_19287)
);

NOR2x1_ASAP7_75t_L g19288 ( 
.A(n_19242),
.B(n_3378),
.Y(n_19288)
);

NAND4xp25_ASAP7_75t_L g19289 ( 
.A(n_19162),
.B(n_3380),
.C(n_3378),
.D(n_3379),
.Y(n_19289)
);

NAND2xp5_ASAP7_75t_L g19290 ( 
.A(n_19207),
.B(n_19120),
.Y(n_19290)
);

AND2x2_ASAP7_75t_L g19291 ( 
.A(n_19231),
.B(n_3379),
.Y(n_19291)
);

HB1xp67_ASAP7_75t_L g19292 ( 
.A(n_19153),
.Y(n_19292)
);

NAND2x1_ASAP7_75t_L g19293 ( 
.A(n_19165),
.B(n_3380),
.Y(n_19293)
);

NAND2xp5_ASAP7_75t_L g19294 ( 
.A(n_19140),
.B(n_3381),
.Y(n_19294)
);

INVx2_ASAP7_75t_L g19295 ( 
.A(n_19195),
.Y(n_19295)
);

AND2x2_ASAP7_75t_L g19296 ( 
.A(n_19128),
.B(n_3381),
.Y(n_19296)
);

NOR2x1_ASAP7_75t_L g19297 ( 
.A(n_19127),
.B(n_3382),
.Y(n_19297)
);

NAND2xp5_ASAP7_75t_L g19298 ( 
.A(n_19181),
.B(n_3382),
.Y(n_19298)
);

OR2x2_ASAP7_75t_L g19299 ( 
.A(n_19169),
.B(n_3383),
.Y(n_19299)
);

NAND2xp5_ASAP7_75t_L g19300 ( 
.A(n_19163),
.B(n_3383),
.Y(n_19300)
);

AND2x2_ASAP7_75t_L g19301 ( 
.A(n_19189),
.B(n_3384),
.Y(n_19301)
);

NAND2xp5_ASAP7_75t_L g19302 ( 
.A(n_19141),
.B(n_3384),
.Y(n_19302)
);

NOR2xp33_ASAP7_75t_SL g19303 ( 
.A(n_19130),
.B(n_3385),
.Y(n_19303)
);

INVx1_ASAP7_75t_L g19304 ( 
.A(n_19129),
.Y(n_19304)
);

INVxp67_ASAP7_75t_L g19305 ( 
.A(n_19144),
.Y(n_19305)
);

INVx1_ASAP7_75t_L g19306 ( 
.A(n_19161),
.Y(n_19306)
);

NAND2xp5_ASAP7_75t_SL g19307 ( 
.A(n_19186),
.B(n_3385),
.Y(n_19307)
);

NAND2xp5_ASAP7_75t_L g19308 ( 
.A(n_19178),
.B(n_3386),
.Y(n_19308)
);

AOI22xp5_ASAP7_75t_L g19309 ( 
.A1(n_19180),
.A2(n_3388),
.B1(n_3386),
.B2(n_3387),
.Y(n_19309)
);

NOR3xp33_ASAP7_75t_L g19310 ( 
.A(n_19174),
.B(n_3387),
.C(n_3388),
.Y(n_19310)
);

NAND2xp5_ASAP7_75t_L g19311 ( 
.A(n_19206),
.B(n_3389),
.Y(n_19311)
);

NAND2xp5_ASAP7_75t_L g19312 ( 
.A(n_19177),
.B(n_3389),
.Y(n_19312)
);

AOI221xp5_ASAP7_75t_SL g19313 ( 
.A1(n_19216),
.A2(n_3392),
.B1(n_3390),
.B2(n_3391),
.C(n_3393),
.Y(n_19313)
);

NOR2xp33_ASAP7_75t_L g19314 ( 
.A(n_19191),
.B(n_3390),
.Y(n_19314)
);

NOR2xp33_ASAP7_75t_L g19315 ( 
.A(n_19244),
.B(n_3391),
.Y(n_19315)
);

NAND2xp5_ASAP7_75t_L g19316 ( 
.A(n_19138),
.B(n_3392),
.Y(n_19316)
);

INVx1_ASAP7_75t_L g19317 ( 
.A(n_19184),
.Y(n_19317)
);

NOR2xp33_ASAP7_75t_L g19318 ( 
.A(n_19233),
.B(n_19213),
.Y(n_19318)
);

NAND2xp5_ASAP7_75t_SL g19319 ( 
.A(n_19241),
.B(n_3393),
.Y(n_19319)
);

NOR2xp33_ASAP7_75t_L g19320 ( 
.A(n_19193),
.B(n_3394),
.Y(n_19320)
);

NAND2xp5_ASAP7_75t_L g19321 ( 
.A(n_19175),
.B(n_3394),
.Y(n_19321)
);

OAI21xp33_ASAP7_75t_L g19322 ( 
.A1(n_19190),
.A2(n_3395),
.B(n_3397),
.Y(n_19322)
);

NAND2xp5_ASAP7_75t_L g19323 ( 
.A(n_19119),
.B(n_19132),
.Y(n_19323)
);

AOI221xp5_ASAP7_75t_L g19324 ( 
.A1(n_19145),
.A2(n_3398),
.B1(n_3395),
.B2(n_3397),
.C(n_3399),
.Y(n_19324)
);

NAND2xp5_ASAP7_75t_L g19325 ( 
.A(n_19232),
.B(n_3399),
.Y(n_19325)
);

AND2x2_ASAP7_75t_L g19326 ( 
.A(n_19198),
.B(n_3400),
.Y(n_19326)
);

AND2x2_ASAP7_75t_L g19327 ( 
.A(n_19155),
.B(n_3400),
.Y(n_19327)
);

AND2x2_ASAP7_75t_L g19328 ( 
.A(n_19123),
.B(n_3401),
.Y(n_19328)
);

OAI221xp5_ASAP7_75t_SL g19329 ( 
.A1(n_19230),
.A2(n_3403),
.B1(n_3401),
.B2(n_3402),
.C(n_3404),
.Y(n_19329)
);

NAND2xp5_ASAP7_75t_L g19330 ( 
.A(n_19240),
.B(n_3402),
.Y(n_19330)
);

NAND2xp5_ASAP7_75t_L g19331 ( 
.A(n_19156),
.B(n_3403),
.Y(n_19331)
);

NAND2xp5_ASAP7_75t_L g19332 ( 
.A(n_19147),
.B(n_3404),
.Y(n_19332)
);

NOR3xp33_ASAP7_75t_L g19333 ( 
.A(n_19142),
.B(n_3405),
.C(n_3406),
.Y(n_19333)
);

NAND2xp5_ASAP7_75t_L g19334 ( 
.A(n_19204),
.B(n_3405),
.Y(n_19334)
);

NAND2xp5_ASAP7_75t_L g19335 ( 
.A(n_19202),
.B(n_3407),
.Y(n_19335)
);

NAND2xp5_ASAP7_75t_L g19336 ( 
.A(n_19212),
.B(n_3407),
.Y(n_19336)
);

OR2x2_ASAP7_75t_L g19337 ( 
.A(n_19228),
.B(n_3408),
.Y(n_19337)
);

AOI22xp5_ASAP7_75t_L g19338 ( 
.A1(n_19176),
.A2(n_3410),
.B1(n_3408),
.B2(n_3409),
.Y(n_19338)
);

INVx2_ASAP7_75t_L g19339 ( 
.A(n_19192),
.Y(n_19339)
);

INVx1_ASAP7_75t_L g19340 ( 
.A(n_19208),
.Y(n_19340)
);

NAND2xp5_ASAP7_75t_L g19341 ( 
.A(n_19237),
.B(n_3410),
.Y(n_19341)
);

INVx1_ASAP7_75t_SL g19342 ( 
.A(n_19170),
.Y(n_19342)
);

NOR2x1_ASAP7_75t_L g19343 ( 
.A(n_19211),
.B(n_3411),
.Y(n_19343)
);

INVx1_ASAP7_75t_L g19344 ( 
.A(n_19125),
.Y(n_19344)
);

INVxp67_ASAP7_75t_L g19345 ( 
.A(n_19200),
.Y(n_19345)
);

NOR3x1_ASAP7_75t_L g19346 ( 
.A(n_19224),
.B(n_3411),
.C(n_3412),
.Y(n_19346)
);

INVx1_ASAP7_75t_L g19347 ( 
.A(n_19164),
.Y(n_19347)
);

AND2x2_ASAP7_75t_L g19348 ( 
.A(n_19227),
.B(n_3412),
.Y(n_19348)
);

NAND2xp33_ASAP7_75t_L g19349 ( 
.A(n_19185),
.B(n_3413),
.Y(n_19349)
);

INVx1_ASAP7_75t_L g19350 ( 
.A(n_19220),
.Y(n_19350)
);

NAND2xp5_ASAP7_75t_SL g19351 ( 
.A(n_19217),
.B(n_3414),
.Y(n_19351)
);

INVx1_ASAP7_75t_L g19352 ( 
.A(n_19168),
.Y(n_19352)
);

INVx1_ASAP7_75t_L g19353 ( 
.A(n_19210),
.Y(n_19353)
);

INVx1_ASAP7_75t_L g19354 ( 
.A(n_19158),
.Y(n_19354)
);

NAND2x1_ASAP7_75t_SL g19355 ( 
.A(n_19218),
.B(n_3415),
.Y(n_19355)
);

INVx2_ASAP7_75t_L g19356 ( 
.A(n_19139),
.Y(n_19356)
);

OR2x2_ASAP7_75t_L g19357 ( 
.A(n_19222),
.B(n_3415),
.Y(n_19357)
);

NAND2xp5_ASAP7_75t_L g19358 ( 
.A(n_19215),
.B(n_3416),
.Y(n_19358)
);

NAND2x1_ASAP7_75t_SL g19359 ( 
.A(n_19194),
.B(n_3416),
.Y(n_19359)
);

OR2x2_ASAP7_75t_L g19360 ( 
.A(n_19219),
.B(n_19146),
.Y(n_19360)
);

INVx2_ASAP7_75t_SL g19361 ( 
.A(n_19150),
.Y(n_19361)
);

NOR2x1_ASAP7_75t_L g19362 ( 
.A(n_19182),
.B(n_3417),
.Y(n_19362)
);

NAND2xp5_ASAP7_75t_L g19363 ( 
.A(n_19167),
.B(n_3417),
.Y(n_19363)
);

NAND2xp5_ASAP7_75t_L g19364 ( 
.A(n_19209),
.B(n_3418),
.Y(n_19364)
);

OAI22xp5_ASAP7_75t_L g19365 ( 
.A1(n_19221),
.A2(n_3422),
.B1(n_3419),
.B2(n_3420),
.Y(n_19365)
);

NAND2xp5_ASAP7_75t_L g19366 ( 
.A(n_19225),
.B(n_3419),
.Y(n_19366)
);

NAND2xp5_ASAP7_75t_L g19367 ( 
.A(n_19199),
.B(n_3420),
.Y(n_19367)
);

NAND2xp5_ASAP7_75t_L g19368 ( 
.A(n_19243),
.B(n_3422),
.Y(n_19368)
);

INVxp67_ASAP7_75t_L g19369 ( 
.A(n_19234),
.Y(n_19369)
);

NOR2xp33_ASAP7_75t_L g19370 ( 
.A(n_19205),
.B(n_3423),
.Y(n_19370)
);

NAND2xp5_ASAP7_75t_L g19371 ( 
.A(n_19152),
.B(n_3423),
.Y(n_19371)
);

NAND2xp5_ASAP7_75t_L g19372 ( 
.A(n_19152),
.B(n_3424),
.Y(n_19372)
);

INVx1_ASAP7_75t_L g19373 ( 
.A(n_19121),
.Y(n_19373)
);

NOR2xp33_ASAP7_75t_L g19374 ( 
.A(n_19121),
.B(n_3424),
.Y(n_19374)
);

INVx2_ASAP7_75t_L g19375 ( 
.A(n_19159),
.Y(n_19375)
);

OAI21xp5_ASAP7_75t_L g19376 ( 
.A1(n_19117),
.A2(n_3425),
.B(n_3426),
.Y(n_19376)
);

NAND3xp33_ASAP7_75t_L g19377 ( 
.A(n_19134),
.B(n_3425),
.C(n_3426),
.Y(n_19377)
);

INVx1_ASAP7_75t_L g19378 ( 
.A(n_19121),
.Y(n_19378)
);

NAND2xp5_ASAP7_75t_L g19379 ( 
.A(n_19152),
.B(n_3427),
.Y(n_19379)
);

NOR2x1_ASAP7_75t_L g19380 ( 
.A(n_19149),
.B(n_3428),
.Y(n_19380)
);

NOR2xp33_ASAP7_75t_L g19381 ( 
.A(n_19121),
.B(n_3428),
.Y(n_19381)
);

NOR3xp33_ASAP7_75t_L g19382 ( 
.A(n_19364),
.B(n_3429),
.C(n_3430),
.Y(n_19382)
);

AOI22xp33_ASAP7_75t_L g19383 ( 
.A1(n_19310),
.A2(n_3432),
.B1(n_3430),
.B2(n_3431),
.Y(n_19383)
);

NAND4xp25_ASAP7_75t_SL g19384 ( 
.A(n_19313),
.B(n_3435),
.C(n_3433),
.D(n_3434),
.Y(n_19384)
);

NOR3xp33_ASAP7_75t_L g19385 ( 
.A(n_19347),
.B(n_3433),
.C(n_3434),
.Y(n_19385)
);

NAND3xp33_ASAP7_75t_L g19386 ( 
.A(n_19264),
.B(n_3436),
.C(n_3437),
.Y(n_19386)
);

NOR3xp33_ASAP7_75t_L g19387 ( 
.A(n_19284),
.B(n_19339),
.C(n_19295),
.Y(n_19387)
);

NAND2xp5_ASAP7_75t_L g19388 ( 
.A(n_19320),
.B(n_3436),
.Y(n_19388)
);

NOR3x1_ASAP7_75t_L g19389 ( 
.A(n_19377),
.B(n_3437),
.C(n_3438),
.Y(n_19389)
);

OAI21xp33_ASAP7_75t_L g19390 ( 
.A1(n_19303),
.A2(n_3439),
.B(n_3440),
.Y(n_19390)
);

NAND4xp75_ASAP7_75t_L g19391 ( 
.A(n_19307),
.B(n_3441),
.C(n_3439),
.D(n_3440),
.Y(n_19391)
);

NAND3xp33_ASAP7_75t_L g19392 ( 
.A(n_19333),
.B(n_3441),
.C(n_3442),
.Y(n_19392)
);

OAI211xp5_ASAP7_75t_L g19393 ( 
.A1(n_19376),
.A2(n_3444),
.B(n_3442),
.C(n_3443),
.Y(n_19393)
);

INVx1_ASAP7_75t_L g19394 ( 
.A(n_19249),
.Y(n_19394)
);

OR2x2_ASAP7_75t_L g19395 ( 
.A(n_19289),
.B(n_19371),
.Y(n_19395)
);

AND2x2_ASAP7_75t_L g19396 ( 
.A(n_19301),
.B(n_3443),
.Y(n_19396)
);

NOR3x1_ASAP7_75t_L g19397 ( 
.A(n_19293),
.B(n_3444),
.C(n_3445),
.Y(n_19397)
);

AOI211xp5_ASAP7_75t_L g19398 ( 
.A1(n_19266),
.A2(n_3447),
.B(n_3445),
.C(n_3446),
.Y(n_19398)
);

OAI211xp5_ASAP7_75t_SL g19399 ( 
.A1(n_19345),
.A2(n_3448),
.B(n_3446),
.C(n_3447),
.Y(n_19399)
);

NAND3xp33_ASAP7_75t_L g19400 ( 
.A(n_19265),
.B(n_3448),
.C(n_3449),
.Y(n_19400)
);

NOR3xp33_ASAP7_75t_L g19401 ( 
.A(n_19305),
.B(n_3449),
.C(n_3450),
.Y(n_19401)
);

AOI211x1_ASAP7_75t_SL g19402 ( 
.A1(n_19316),
.A2(n_3452),
.B(n_3450),
.C(n_3451),
.Y(n_19402)
);

OAI211xp5_ASAP7_75t_L g19403 ( 
.A1(n_19256),
.A2(n_3453),
.B(n_3451),
.C(n_3452),
.Y(n_19403)
);

NOR2x1_ASAP7_75t_L g19404 ( 
.A(n_19288),
.B(n_3454),
.Y(n_19404)
);

NAND3xp33_ASAP7_75t_L g19405 ( 
.A(n_19246),
.B(n_19351),
.C(n_19324),
.Y(n_19405)
);

NOR2x1_ASAP7_75t_L g19406 ( 
.A(n_19253),
.B(n_3454),
.Y(n_19406)
);

OR2x2_ASAP7_75t_L g19407 ( 
.A(n_19372),
.B(n_3455),
.Y(n_19407)
);

AOI221xp5_ASAP7_75t_L g19408 ( 
.A1(n_19370),
.A2(n_3457),
.B1(n_3455),
.B2(n_3456),
.C(n_3458),
.Y(n_19408)
);

NOR2x1_ASAP7_75t_L g19409 ( 
.A(n_19260),
.B(n_3457),
.Y(n_19409)
);

NOR2x1_ASAP7_75t_L g19410 ( 
.A(n_19375),
.B(n_3458),
.Y(n_19410)
);

AOI32xp33_ASAP7_75t_L g19411 ( 
.A1(n_19250),
.A2(n_3461),
.A3(n_3459),
.B1(n_3460),
.B2(n_3462),
.Y(n_19411)
);

NOR2x1_ASAP7_75t_L g19412 ( 
.A(n_19255),
.B(n_3459),
.Y(n_19412)
);

NOR2x1_ASAP7_75t_L g19413 ( 
.A(n_19251),
.B(n_3460),
.Y(n_19413)
);

NOR2x1_ASAP7_75t_L g19414 ( 
.A(n_19380),
.B(n_3461),
.Y(n_19414)
);

NAND2xp5_ASAP7_75t_L g19415 ( 
.A(n_19374),
.B(n_3462),
.Y(n_19415)
);

INVx1_ASAP7_75t_L g19416 ( 
.A(n_19248),
.Y(n_19416)
);

NAND2xp5_ASAP7_75t_SL g19417 ( 
.A(n_19338),
.B(n_3463),
.Y(n_19417)
);

INVx1_ASAP7_75t_L g19418 ( 
.A(n_19379),
.Y(n_19418)
);

NAND5xp2_ASAP7_75t_L g19419 ( 
.A(n_19269),
.B(n_3465),
.C(n_3463),
.D(n_3464),
.E(n_3466),
.Y(n_19419)
);

NAND2xp5_ASAP7_75t_SL g19420 ( 
.A(n_19263),
.B(n_3464),
.Y(n_19420)
);

OAI211xp5_ASAP7_75t_L g19421 ( 
.A1(n_19368),
.A2(n_3468),
.B(n_3466),
.C(n_3467),
.Y(n_19421)
);

AOI22xp5_ASAP7_75t_L g19422 ( 
.A1(n_19369),
.A2(n_3469),
.B1(n_3467),
.B2(n_3468),
.Y(n_19422)
);

AOI221xp5_ASAP7_75t_L g19423 ( 
.A1(n_19270),
.A2(n_3471),
.B1(n_3469),
.B2(n_3470),
.C(n_3472),
.Y(n_19423)
);

NAND2xp5_ASAP7_75t_L g19424 ( 
.A(n_19381),
.B(n_19286),
.Y(n_19424)
);

NOR3xp33_ASAP7_75t_L g19425 ( 
.A(n_19317),
.B(n_3470),
.C(n_3471),
.Y(n_19425)
);

NAND3xp33_ASAP7_75t_SL g19426 ( 
.A(n_19252),
.B(n_3472),
.C(n_3473),
.Y(n_19426)
);

OAI221xp5_ASAP7_75t_L g19427 ( 
.A1(n_19267),
.A2(n_3475),
.B1(n_3473),
.B2(n_3474),
.C(n_3476),
.Y(n_19427)
);

NAND4xp25_ASAP7_75t_L g19428 ( 
.A(n_19315),
.B(n_19318),
.C(n_19314),
.D(n_19298),
.Y(n_19428)
);

AOI21xp5_ASAP7_75t_L g19429 ( 
.A1(n_19287),
.A2(n_3474),
.B(n_3476),
.Y(n_19429)
);

NAND2xp5_ASAP7_75t_L g19430 ( 
.A(n_19309),
.B(n_3477),
.Y(n_19430)
);

OAI211xp5_ASAP7_75t_SL g19431 ( 
.A1(n_19276),
.A2(n_3479),
.B(n_3477),
.C(n_3478),
.Y(n_19431)
);

OAI21xp33_ASAP7_75t_SL g19432 ( 
.A1(n_19359),
.A2(n_3478),
.B(n_3479),
.Y(n_19432)
);

NAND2xp5_ASAP7_75t_L g19433 ( 
.A(n_19322),
.B(n_3480),
.Y(n_19433)
);

A2O1A1Ixp33_ASAP7_75t_L g19434 ( 
.A1(n_19272),
.A2(n_3482),
.B(n_3480),
.C(n_3481),
.Y(n_19434)
);

BUFx2_ASAP7_75t_L g19435 ( 
.A(n_19259),
.Y(n_19435)
);

NAND4xp25_ASAP7_75t_L g19436 ( 
.A(n_19362),
.B(n_3483),
.C(n_3481),
.D(n_3482),
.Y(n_19436)
);

NAND3xp33_ASAP7_75t_L g19437 ( 
.A(n_19292),
.B(n_3483),
.C(n_3484),
.Y(n_19437)
);

NAND4xp25_ASAP7_75t_L g19438 ( 
.A(n_19271),
.B(n_19281),
.C(n_19277),
.D(n_19335),
.Y(n_19438)
);

NOR3xp33_ASAP7_75t_L g19439 ( 
.A(n_19353),
.B(n_3484),
.C(n_3485),
.Y(n_19439)
);

NOR3x1_ASAP7_75t_L g19440 ( 
.A(n_19325),
.B(n_3485),
.C(n_3486),
.Y(n_19440)
);

NAND3xp33_ASAP7_75t_SL g19441 ( 
.A(n_19282),
.B(n_3486),
.C(n_3487),
.Y(n_19441)
);

NAND4xp25_ASAP7_75t_L g19442 ( 
.A(n_19343),
.B(n_3490),
.C(n_3488),
.D(n_3489),
.Y(n_19442)
);

INVx1_ASAP7_75t_L g19443 ( 
.A(n_19245),
.Y(n_19443)
);

NAND3xp33_ASAP7_75t_SL g19444 ( 
.A(n_19273),
.B(n_3488),
.C(n_3489),
.Y(n_19444)
);

NAND4xp25_ASAP7_75t_L g19445 ( 
.A(n_19294),
.B(n_3492),
.C(n_3490),
.D(n_3491),
.Y(n_19445)
);

OAI21xp33_ASAP7_75t_L g19446 ( 
.A1(n_19306),
.A2(n_19291),
.B(n_19247),
.Y(n_19446)
);

INVx1_ASAP7_75t_L g19447 ( 
.A(n_19346),
.Y(n_19447)
);

NOR2xp67_ASAP7_75t_L g19448 ( 
.A(n_19365),
.B(n_3492),
.Y(n_19448)
);

NAND3xp33_ASAP7_75t_L g19449 ( 
.A(n_19349),
.B(n_3493),
.C(n_3494),
.Y(n_19449)
);

OA211x2_ASAP7_75t_L g19450 ( 
.A1(n_19258),
.A2(n_3495),
.B(n_3493),
.C(n_3494),
.Y(n_19450)
);

NAND2xp5_ASAP7_75t_L g19451 ( 
.A(n_19296),
.B(n_3495),
.Y(n_19451)
);

NOR3x1_ASAP7_75t_L g19452 ( 
.A(n_19330),
.B(n_3496),
.C(n_3497),
.Y(n_19452)
);

INVxp67_ASAP7_75t_L g19453 ( 
.A(n_19327),
.Y(n_19453)
);

AOI22xp5_ASAP7_75t_L g19454 ( 
.A1(n_19304),
.A2(n_3498),
.B1(n_3496),
.B2(n_3497),
.Y(n_19454)
);

AND4x1_ASAP7_75t_L g19455 ( 
.A(n_19262),
.B(n_3500),
.C(n_3498),
.D(n_3499),
.Y(n_19455)
);

NOR3xp33_ASAP7_75t_SL g19456 ( 
.A(n_19283),
.B(n_3499),
.C(n_3500),
.Y(n_19456)
);

OAI221xp5_ASAP7_75t_SL g19457 ( 
.A1(n_19254),
.A2(n_3503),
.B1(n_3501),
.B2(n_3502),
.C(n_3504),
.Y(n_19457)
);

NAND3xp33_ASAP7_75t_SL g19458 ( 
.A(n_19342),
.B(n_3501),
.C(n_3502),
.Y(n_19458)
);

NAND4xp25_ASAP7_75t_L g19459 ( 
.A(n_19331),
.B(n_3506),
.C(n_3504),
.D(n_3505),
.Y(n_19459)
);

NAND4xp25_ASAP7_75t_L g19460 ( 
.A(n_19268),
.B(n_19363),
.C(n_19297),
.D(n_19312),
.Y(n_19460)
);

NAND2xp5_ASAP7_75t_L g19461 ( 
.A(n_19355),
.B(n_3505),
.Y(n_19461)
);

NOR3xp33_ASAP7_75t_L g19462 ( 
.A(n_19344),
.B(n_3506),
.C(n_3507),
.Y(n_19462)
);

INVx1_ASAP7_75t_L g19463 ( 
.A(n_19279),
.Y(n_19463)
);

NAND2xp5_ASAP7_75t_L g19464 ( 
.A(n_19285),
.B(n_3508),
.Y(n_19464)
);

AOI21xp5_ASAP7_75t_L g19465 ( 
.A1(n_19332),
.A2(n_3509),
.B(n_3510),
.Y(n_19465)
);

NOR3xp33_ASAP7_75t_L g19466 ( 
.A(n_19280),
.B(n_3509),
.C(n_3510),
.Y(n_19466)
);

NAND2xp5_ASAP7_75t_L g19467 ( 
.A(n_19257),
.B(n_3511),
.Y(n_19467)
);

NAND3x1_ASAP7_75t_L g19468 ( 
.A(n_19300),
.B(n_3511),
.C(n_3512),
.Y(n_19468)
);

INVx1_ASAP7_75t_L g19469 ( 
.A(n_19334),
.Y(n_19469)
);

NAND2xp5_ASAP7_75t_L g19470 ( 
.A(n_19261),
.B(n_3512),
.Y(n_19470)
);

NAND3xp33_ASAP7_75t_L g19471 ( 
.A(n_19350),
.B(n_3513),
.C(n_3514),
.Y(n_19471)
);

NAND2xp5_ASAP7_75t_L g19472 ( 
.A(n_19361),
.B(n_3513),
.Y(n_19472)
);

AOI221xp5_ASAP7_75t_L g19473 ( 
.A1(n_19319),
.A2(n_19358),
.B1(n_19367),
.B2(n_19340),
.C(n_19341),
.Y(n_19473)
);

OAI221xp5_ASAP7_75t_L g19474 ( 
.A1(n_19321),
.A2(n_3517),
.B1(n_3515),
.B2(n_3516),
.C(n_3518),
.Y(n_19474)
);

NOR3xp33_ASAP7_75t_L g19475 ( 
.A(n_19352),
.B(n_3515),
.C(n_3516),
.Y(n_19475)
);

NAND2xp5_ASAP7_75t_L g19476 ( 
.A(n_19336),
.B(n_3518),
.Y(n_19476)
);

NAND2xp5_ASAP7_75t_L g19477 ( 
.A(n_19373),
.B(n_19378),
.Y(n_19477)
);

NOR3x1_ASAP7_75t_L g19478 ( 
.A(n_19311),
.B(n_3519),
.C(n_3520),
.Y(n_19478)
);

NOR3x1_ASAP7_75t_L g19479 ( 
.A(n_19308),
.B(n_3521),
.C(n_3522),
.Y(n_19479)
);

AOI211xp5_ASAP7_75t_SL g19480 ( 
.A1(n_19354),
.A2(n_3524),
.B(n_3521),
.C(n_3523),
.Y(n_19480)
);

NOR2xp33_ASAP7_75t_L g19481 ( 
.A(n_19299),
.B(n_3523),
.Y(n_19481)
);

NOR2xp33_ASAP7_75t_L g19482 ( 
.A(n_19357),
.B(n_3524),
.Y(n_19482)
);

NOR3xp33_ASAP7_75t_L g19483 ( 
.A(n_19274),
.B(n_3525),
.C(n_3526),
.Y(n_19483)
);

NOR3xp33_ASAP7_75t_L g19484 ( 
.A(n_19356),
.B(n_3525),
.C(n_3526),
.Y(n_19484)
);

AOI22xp5_ASAP7_75t_L g19485 ( 
.A1(n_19323),
.A2(n_3529),
.B1(n_3527),
.B2(n_3528),
.Y(n_19485)
);

AOI211xp5_ASAP7_75t_SL g19486 ( 
.A1(n_19290),
.A2(n_3529),
.B(n_3527),
.C(n_3528),
.Y(n_19486)
);

NOR5xp2_ASAP7_75t_L g19487 ( 
.A(n_19329),
.B(n_3532),
.C(n_3530),
.D(n_3531),
.E(n_3533),
.Y(n_19487)
);

NAND4xp25_ASAP7_75t_L g19488 ( 
.A(n_19366),
.B(n_3533),
.C(n_3531),
.D(n_3532),
.Y(n_19488)
);

AOI221x1_ASAP7_75t_L g19489 ( 
.A1(n_19302),
.A2(n_3536),
.B1(n_3534),
.B2(n_3535),
.C(n_3537),
.Y(n_19489)
);

NAND2xp5_ASAP7_75t_L g19490 ( 
.A(n_19278),
.B(n_3534),
.Y(n_19490)
);

NAND2xp5_ASAP7_75t_L g19491 ( 
.A(n_19328),
.B(n_3535),
.Y(n_19491)
);

NAND4xp25_ASAP7_75t_SL g19492 ( 
.A(n_19337),
.B(n_3539),
.C(n_3536),
.D(n_3538),
.Y(n_19492)
);

NOR5xp2_ASAP7_75t_L g19493 ( 
.A(n_19360),
.B(n_3541),
.C(n_3538),
.D(n_3540),
.E(n_3542),
.Y(n_19493)
);

NOR3x1_ASAP7_75t_L g19494 ( 
.A(n_19275),
.B(n_3540),
.C(n_3541),
.Y(n_19494)
);

NOR5xp2_ASAP7_75t_L g19495 ( 
.A(n_19326),
.B(n_3544),
.C(n_3542),
.D(n_3543),
.E(n_3545),
.Y(n_19495)
);

NOR4xp25_ASAP7_75t_L g19496 ( 
.A(n_19348),
.B(n_3545),
.C(n_3543),
.D(n_3544),
.Y(n_19496)
);

NOR3xp33_ASAP7_75t_L g19497 ( 
.A(n_19364),
.B(n_3546),
.C(n_3547),
.Y(n_19497)
);

NAND2xp5_ASAP7_75t_L g19498 ( 
.A(n_19320),
.B(n_3547),
.Y(n_19498)
);

NOR2xp67_ASAP7_75t_L g19499 ( 
.A(n_19289),
.B(n_3548),
.Y(n_19499)
);

OAI211xp5_ASAP7_75t_L g19500 ( 
.A1(n_19376),
.A2(n_3550),
.B(n_3548),
.C(n_3549),
.Y(n_19500)
);

OAI211xp5_ASAP7_75t_SL g19501 ( 
.A1(n_19364),
.A2(n_3551),
.B(n_3549),
.C(n_3550),
.Y(n_19501)
);

OR2x2_ASAP7_75t_L g19502 ( 
.A(n_19289),
.B(n_3551),
.Y(n_19502)
);

NAND2xp5_ASAP7_75t_SL g19503 ( 
.A(n_19338),
.B(n_3552),
.Y(n_19503)
);

NOR2x1_ASAP7_75t_L g19504 ( 
.A(n_19288),
.B(n_3552),
.Y(n_19504)
);

NOR2xp33_ASAP7_75t_L g19505 ( 
.A(n_19256),
.B(n_3553),
.Y(n_19505)
);

NAND2xp5_ASAP7_75t_SL g19506 ( 
.A(n_19338),
.B(n_3554),
.Y(n_19506)
);

AOI211xp5_ASAP7_75t_L g19507 ( 
.A1(n_19310),
.A2(n_3557),
.B(n_3555),
.C(n_3556),
.Y(n_19507)
);

NOR2xp33_ASAP7_75t_SL g19508 ( 
.A(n_19252),
.B(n_3555),
.Y(n_19508)
);

NAND4xp25_ASAP7_75t_SL g19509 ( 
.A(n_19313),
.B(n_3558),
.C(n_3556),
.D(n_3557),
.Y(n_19509)
);

NOR2xp33_ASAP7_75t_L g19510 ( 
.A(n_19256),
.B(n_3558),
.Y(n_19510)
);

INVx1_ASAP7_75t_L g19511 ( 
.A(n_19249),
.Y(n_19511)
);

OAI21xp5_ASAP7_75t_L g19512 ( 
.A1(n_19369),
.A2(n_3559),
.B(n_3560),
.Y(n_19512)
);

NAND2xp5_ASAP7_75t_L g19513 ( 
.A(n_19320),
.B(n_3559),
.Y(n_19513)
);

OAI321xp33_ASAP7_75t_L g19514 ( 
.A1(n_19289),
.A2(n_3562),
.A3(n_3564),
.B1(n_3560),
.B2(n_3561),
.C(n_3563),
.Y(n_19514)
);

NAND2xp5_ASAP7_75t_L g19515 ( 
.A(n_19320),
.B(n_3563),
.Y(n_19515)
);

NOR4xp25_ASAP7_75t_L g19516 ( 
.A(n_19307),
.B(n_3566),
.C(n_3564),
.D(n_3565),
.Y(n_19516)
);

OAI221xp5_ASAP7_75t_L g19517 ( 
.A1(n_19310),
.A2(n_3568),
.B1(n_3566),
.B2(n_3567),
.C(n_3569),
.Y(n_19517)
);

AOI221x1_ASAP7_75t_L g19518 ( 
.A1(n_19364),
.A2(n_3569),
.B1(n_3567),
.B2(n_3568),
.C(n_3570),
.Y(n_19518)
);

AOI211xp5_ASAP7_75t_L g19519 ( 
.A1(n_19310),
.A2(n_3572),
.B(n_3570),
.C(n_3571),
.Y(n_19519)
);

NOR3xp33_ASAP7_75t_L g19520 ( 
.A(n_19364),
.B(n_3571),
.C(n_3572),
.Y(n_19520)
);

NAND4xp25_ASAP7_75t_L g19521 ( 
.A(n_19310),
.B(n_3575),
.C(n_3573),
.D(n_3574),
.Y(n_19521)
);

NAND4xp25_ASAP7_75t_L g19522 ( 
.A(n_19310),
.B(n_3576),
.C(n_3573),
.D(n_3574),
.Y(n_19522)
);

OAI21xp33_ASAP7_75t_L g19523 ( 
.A1(n_19284),
.A2(n_3576),
.B(n_3577),
.Y(n_19523)
);

NOR2x1_ASAP7_75t_L g19524 ( 
.A(n_19288),
.B(n_3577),
.Y(n_19524)
);

AOI221x1_ASAP7_75t_L g19525 ( 
.A1(n_19364),
.A2(n_3580),
.B1(n_3578),
.B2(n_3579),
.C(n_3582),
.Y(n_19525)
);

NAND2xp5_ASAP7_75t_L g19526 ( 
.A(n_19320),
.B(n_3578),
.Y(n_19526)
);

NAND2xp5_ASAP7_75t_L g19527 ( 
.A(n_19320),
.B(n_3582),
.Y(n_19527)
);

OAI21xp5_ASAP7_75t_L g19528 ( 
.A1(n_19369),
.A2(n_3583),
.B(n_3584),
.Y(n_19528)
);

INVx1_ASAP7_75t_L g19529 ( 
.A(n_19249),
.Y(n_19529)
);

NAND4xp25_ASAP7_75t_L g19530 ( 
.A(n_19310),
.B(n_3585),
.C(n_3583),
.D(n_3584),
.Y(n_19530)
);

NOR2xp33_ASAP7_75t_L g19531 ( 
.A(n_19256),
.B(n_3586),
.Y(n_19531)
);

AOI21xp5_ASAP7_75t_L g19532 ( 
.A1(n_19287),
.A2(n_3586),
.B(n_3587),
.Y(n_19532)
);

NOR2x1_ASAP7_75t_L g19533 ( 
.A(n_19288),
.B(n_3587),
.Y(n_19533)
);

NOR2xp33_ASAP7_75t_L g19534 ( 
.A(n_19256),
.B(n_3588),
.Y(n_19534)
);

NOR3xp33_ASAP7_75t_SL g19535 ( 
.A(n_19307),
.B(n_3589),
.C(n_3590),
.Y(n_19535)
);

OA211x2_ASAP7_75t_L g19536 ( 
.A1(n_19293),
.A2(n_3591),
.B(n_3589),
.C(n_3590),
.Y(n_19536)
);

NAND3xp33_ASAP7_75t_SL g19537 ( 
.A(n_19252),
.B(n_3591),
.C(n_3592),
.Y(n_19537)
);

NAND2xp5_ASAP7_75t_L g19538 ( 
.A(n_19320),
.B(n_3592),
.Y(n_19538)
);

NAND2xp5_ASAP7_75t_SL g19539 ( 
.A(n_19338),
.B(n_3593),
.Y(n_19539)
);

NOR3xp33_ASAP7_75t_L g19540 ( 
.A(n_19364),
.B(n_3593),
.C(n_3594),
.Y(n_19540)
);

NAND4xp25_ASAP7_75t_L g19541 ( 
.A(n_19310),
.B(n_3596),
.C(n_3594),
.D(n_3595),
.Y(n_19541)
);

OAI21xp33_ASAP7_75t_L g19542 ( 
.A1(n_19284),
.A2(n_3597),
.B(n_3598),
.Y(n_19542)
);

NOR2x1_ASAP7_75t_L g19543 ( 
.A(n_19288),
.B(n_3598),
.Y(n_19543)
);

NAND3xp33_ASAP7_75t_L g19544 ( 
.A(n_19264),
.B(n_3599),
.C(n_3600),
.Y(n_19544)
);

NAND2xp5_ASAP7_75t_L g19545 ( 
.A(n_19320),
.B(n_3599),
.Y(n_19545)
);

NAND4xp75_ASAP7_75t_L g19546 ( 
.A(n_19307),
.B(n_3602),
.C(n_3600),
.D(n_3601),
.Y(n_19546)
);

NAND3xp33_ASAP7_75t_SL g19547 ( 
.A(n_19252),
.B(n_3603),
.C(n_3604),
.Y(n_19547)
);

AOI211xp5_ASAP7_75t_L g19548 ( 
.A1(n_19310),
.A2(n_3606),
.B(n_3603),
.C(n_3605),
.Y(n_19548)
);

NOR2x1_ASAP7_75t_L g19549 ( 
.A(n_19288),
.B(n_3605),
.Y(n_19549)
);

NAND3xp33_ASAP7_75t_L g19550 ( 
.A(n_19264),
.B(n_3606),
.C(n_3607),
.Y(n_19550)
);

NAND2xp5_ASAP7_75t_SL g19551 ( 
.A(n_19338),
.B(n_3607),
.Y(n_19551)
);

NOR3xp33_ASAP7_75t_SL g19552 ( 
.A(n_19307),
.B(n_3608),
.C(n_3609),
.Y(n_19552)
);

OAI211xp5_ASAP7_75t_L g19553 ( 
.A1(n_19376),
.A2(n_3611),
.B(n_3609),
.C(n_3610),
.Y(n_19553)
);

AO221x1_ASAP7_75t_L g19554 ( 
.A1(n_19369),
.A2(n_3613),
.B1(n_3610),
.B2(n_3612),
.C(n_3614),
.Y(n_19554)
);

NAND3xp33_ASAP7_75t_L g19555 ( 
.A(n_19264),
.B(n_3613),
.C(n_3614),
.Y(n_19555)
);

NOR3xp33_ASAP7_75t_L g19556 ( 
.A(n_19364),
.B(n_3615),
.C(n_3616),
.Y(n_19556)
);

NAND3xp33_ASAP7_75t_SL g19557 ( 
.A(n_19252),
.B(n_3615),
.C(n_3616),
.Y(n_19557)
);

NOR2xp67_ASAP7_75t_L g19558 ( 
.A(n_19289),
.B(n_3617),
.Y(n_19558)
);

NAND3xp33_ASAP7_75t_L g19559 ( 
.A(n_19264),
.B(n_3618),
.C(n_3619),
.Y(n_19559)
);

NOR3x1_ASAP7_75t_SL g19560 ( 
.A(n_19292),
.B(n_3618),
.C(n_3620),
.Y(n_19560)
);

OAI211xp5_ASAP7_75t_SL g19561 ( 
.A1(n_19364),
.A2(n_3622),
.B(n_3620),
.C(n_3621),
.Y(n_19561)
);

NAND4xp25_ASAP7_75t_L g19562 ( 
.A(n_19310),
.B(n_3623),
.C(n_3621),
.D(n_3622),
.Y(n_19562)
);

OAI211xp5_ASAP7_75t_SL g19563 ( 
.A1(n_19364),
.A2(n_3625),
.B(n_3623),
.C(n_3624),
.Y(n_19563)
);

NAND2xp5_ASAP7_75t_L g19564 ( 
.A(n_19320),
.B(n_3624),
.Y(n_19564)
);

NAND2xp5_ASAP7_75t_SL g19565 ( 
.A(n_19338),
.B(n_3625),
.Y(n_19565)
);

NAND4xp25_ASAP7_75t_L g19566 ( 
.A(n_19310),
.B(n_3628),
.C(n_3626),
.D(n_3627),
.Y(n_19566)
);

OAI211xp5_ASAP7_75t_L g19567 ( 
.A1(n_19376),
.A2(n_3630),
.B(n_3628),
.C(n_3629),
.Y(n_19567)
);

AOI211xp5_ASAP7_75t_L g19568 ( 
.A1(n_19310),
.A2(n_3632),
.B(n_3630),
.C(n_3631),
.Y(n_19568)
);

NAND2xp5_ASAP7_75t_L g19569 ( 
.A(n_19320),
.B(n_3631),
.Y(n_19569)
);

NAND2xp5_ASAP7_75t_SL g19570 ( 
.A(n_19338),
.B(n_3632),
.Y(n_19570)
);

NOR3x1_ASAP7_75t_SL g19571 ( 
.A(n_19292),
.B(n_3633),
.C(n_3634),
.Y(n_19571)
);

NOR3xp33_ASAP7_75t_L g19572 ( 
.A(n_19364),
.B(n_3633),
.C(n_3634),
.Y(n_19572)
);

NOR3xp33_ASAP7_75t_L g19573 ( 
.A(n_19364),
.B(n_3635),
.C(n_3636),
.Y(n_19573)
);

NOR4xp25_ASAP7_75t_L g19574 ( 
.A(n_19307),
.B(n_3637),
.C(n_3635),
.D(n_3636),
.Y(n_19574)
);

NOR3x1_ASAP7_75t_L g19575 ( 
.A(n_19264),
.B(n_3638),
.C(n_3639),
.Y(n_19575)
);

NOR3xp33_ASAP7_75t_L g19576 ( 
.A(n_19364),
.B(n_3638),
.C(n_3639),
.Y(n_19576)
);

NOR2xp67_ASAP7_75t_L g19577 ( 
.A(n_19289),
.B(n_3640),
.Y(n_19577)
);

INVx1_ASAP7_75t_L g19578 ( 
.A(n_19249),
.Y(n_19578)
);

NOR2xp33_ASAP7_75t_SL g19579 ( 
.A(n_19252),
.B(n_3641),
.Y(n_19579)
);

NAND3xp33_ASAP7_75t_L g19580 ( 
.A(n_19264),
.B(n_3642),
.C(n_3643),
.Y(n_19580)
);

NAND5xp2_ASAP7_75t_L g19581 ( 
.A(n_19303),
.B(n_3644),
.C(n_3642),
.D(n_3643),
.E(n_3645),
.Y(n_19581)
);

AOI21xp5_ASAP7_75t_L g19582 ( 
.A1(n_19287),
.A2(n_3644),
.B(n_3645),
.Y(n_19582)
);

NOR4xp25_ASAP7_75t_L g19583 ( 
.A(n_19307),
.B(n_3648),
.C(n_3646),
.D(n_3647),
.Y(n_19583)
);

NAND3xp33_ASAP7_75t_L g19584 ( 
.A(n_19264),
.B(n_3647),
.C(n_3648),
.Y(n_19584)
);

INVx1_ASAP7_75t_L g19585 ( 
.A(n_19249),
.Y(n_19585)
);

OAI211xp5_ASAP7_75t_L g19586 ( 
.A1(n_19376),
.A2(n_3651),
.B(n_3649),
.C(n_3650),
.Y(n_19586)
);

NOR3xp33_ASAP7_75t_L g19587 ( 
.A(n_19364),
.B(n_3649),
.C(n_3650),
.Y(n_19587)
);

NAND4xp75_ASAP7_75t_L g19588 ( 
.A(n_19307),
.B(n_3653),
.C(n_3651),
.D(n_3652),
.Y(n_19588)
);

NOR2xp33_ASAP7_75t_L g19589 ( 
.A(n_19256),
.B(n_3652),
.Y(n_19589)
);

NAND3xp33_ASAP7_75t_L g19590 ( 
.A(n_19264),
.B(n_3653),
.C(n_3654),
.Y(n_19590)
);

NOR2xp33_ASAP7_75t_L g19591 ( 
.A(n_19442),
.B(n_3654),
.Y(n_19591)
);

OAI22xp33_ASAP7_75t_L g19592 ( 
.A1(n_19508),
.A2(n_3657),
.B1(n_3655),
.B2(n_3656),
.Y(n_19592)
);

NAND2xp5_ASAP7_75t_L g19593 ( 
.A(n_19396),
.B(n_3655),
.Y(n_19593)
);

OAI22xp5_ASAP7_75t_L g19594 ( 
.A1(n_19383),
.A2(n_3658),
.B1(n_3656),
.B2(n_3657),
.Y(n_19594)
);

NAND2xp5_ASAP7_75t_L g19595 ( 
.A(n_19411),
.B(n_3658),
.Y(n_19595)
);

A2O1A1Ixp33_ASAP7_75t_L g19596 ( 
.A1(n_19481),
.A2(n_3661),
.B(n_3659),
.C(n_3660),
.Y(n_19596)
);

INVxp67_ASAP7_75t_SL g19597 ( 
.A(n_19413),
.Y(n_19597)
);

INVx1_ASAP7_75t_L g19598 ( 
.A(n_19560),
.Y(n_19598)
);

INVx1_ASAP7_75t_L g19599 ( 
.A(n_19571),
.Y(n_19599)
);

INVx1_ASAP7_75t_L g19600 ( 
.A(n_19536),
.Y(n_19600)
);

NOR2xp33_ASAP7_75t_L g19601 ( 
.A(n_19436),
.B(n_3659),
.Y(n_19601)
);

AOI22xp5_ASAP7_75t_L g19602 ( 
.A1(n_19387),
.A2(n_3663),
.B1(n_3660),
.B2(n_3662),
.Y(n_19602)
);

INVx1_ASAP7_75t_L g19603 ( 
.A(n_19412),
.Y(n_19603)
);

AO22x1_ASAP7_75t_L g19604 ( 
.A1(n_19414),
.A2(n_3665),
.B1(n_3663),
.B2(n_3664),
.Y(n_19604)
);

INVx1_ASAP7_75t_L g19605 ( 
.A(n_19406),
.Y(n_19605)
);

AOI22xp5_ASAP7_75t_L g19606 ( 
.A1(n_19499),
.A2(n_3666),
.B1(n_3664),
.B2(n_3665),
.Y(n_19606)
);

INVx2_ASAP7_75t_L g19607 ( 
.A(n_19554),
.Y(n_19607)
);

AOI22xp5_ASAP7_75t_L g19608 ( 
.A1(n_19558),
.A2(n_3668),
.B1(n_3666),
.B2(n_3667),
.Y(n_19608)
);

INVx1_ASAP7_75t_L g19609 ( 
.A(n_19409),
.Y(n_19609)
);

NOR2x1_ASAP7_75t_L g19610 ( 
.A(n_19410),
.B(n_3667),
.Y(n_19610)
);

INVx1_ASAP7_75t_L g19611 ( 
.A(n_19404),
.Y(n_19611)
);

INVx1_ASAP7_75t_L g19612 ( 
.A(n_19504),
.Y(n_19612)
);

AOI22xp5_ASAP7_75t_L g19613 ( 
.A1(n_19577),
.A2(n_3670),
.B1(n_3668),
.B2(n_3669),
.Y(n_19613)
);

OAI22xp5_ASAP7_75t_L g19614 ( 
.A1(n_19464),
.A2(n_3671),
.B1(n_3669),
.B2(n_3670),
.Y(n_19614)
);

INVx1_ASAP7_75t_L g19615 ( 
.A(n_19524),
.Y(n_19615)
);

INVx1_ASAP7_75t_L g19616 ( 
.A(n_19533),
.Y(n_19616)
);

NOR2xp67_ASAP7_75t_L g19617 ( 
.A(n_19441),
.B(n_3671),
.Y(n_19617)
);

NOR2xp33_ASAP7_75t_L g19618 ( 
.A(n_19432),
.B(n_3673),
.Y(n_19618)
);

AO22x2_ASAP7_75t_L g19619 ( 
.A1(n_19394),
.A2(n_3677),
.B1(n_3674),
.B2(n_3676),
.Y(n_19619)
);

AOI22xp33_ASAP7_75t_L g19620 ( 
.A1(n_19384),
.A2(n_3677),
.B1(n_3674),
.B2(n_3676),
.Y(n_19620)
);

INVx2_ASAP7_75t_L g19621 ( 
.A(n_19397),
.Y(n_19621)
);

INVx1_ASAP7_75t_L g19622 ( 
.A(n_19543),
.Y(n_19622)
);

NAND2xp5_ASAP7_75t_L g19623 ( 
.A(n_19496),
.B(n_3678),
.Y(n_19623)
);

INVx1_ASAP7_75t_L g19624 ( 
.A(n_19549),
.Y(n_19624)
);

NOR2x1_ASAP7_75t_L g19625 ( 
.A(n_19435),
.B(n_3679),
.Y(n_19625)
);

INVx1_ASAP7_75t_L g19626 ( 
.A(n_19450),
.Y(n_19626)
);

OA22x2_ASAP7_75t_L g19627 ( 
.A1(n_19393),
.A2(n_3681),
.B1(n_3679),
.B2(n_3680),
.Y(n_19627)
);

NAND2xp5_ASAP7_75t_L g19628 ( 
.A(n_19456),
.B(n_3680),
.Y(n_19628)
);

INVx1_ASAP7_75t_L g19629 ( 
.A(n_19451),
.Y(n_19629)
);

INVx2_ASAP7_75t_L g19630 ( 
.A(n_19391),
.Y(n_19630)
);

NOR4xp25_ASAP7_75t_L g19631 ( 
.A(n_19390),
.B(n_3683),
.C(n_3681),
.D(n_3682),
.Y(n_19631)
);

AOI22xp5_ASAP7_75t_L g19632 ( 
.A1(n_19579),
.A2(n_3684),
.B1(n_3682),
.B2(n_3683),
.Y(n_19632)
);

INVx1_ASAP7_75t_L g19633 ( 
.A(n_19461),
.Y(n_19633)
);

O2A1O1Ixp33_ASAP7_75t_L g19634 ( 
.A1(n_19434),
.A2(n_3686),
.B(n_3684),
.C(n_3685),
.Y(n_19634)
);

INVx1_ASAP7_75t_L g19635 ( 
.A(n_19490),
.Y(n_19635)
);

INVxp67_ASAP7_75t_L g19636 ( 
.A(n_19491),
.Y(n_19636)
);

INVx1_ASAP7_75t_L g19637 ( 
.A(n_19502),
.Y(n_19637)
);

NAND2xp5_ASAP7_75t_SL g19638 ( 
.A(n_19514),
.B(n_3685),
.Y(n_19638)
);

INVxp67_ASAP7_75t_SL g19639 ( 
.A(n_19468),
.Y(n_19639)
);

AOI22xp5_ASAP7_75t_L g19640 ( 
.A1(n_19426),
.A2(n_19537),
.B1(n_19557),
.B2(n_19547),
.Y(n_19640)
);

INVx1_ASAP7_75t_L g19641 ( 
.A(n_19476),
.Y(n_19641)
);

INVx2_ASAP7_75t_L g19642 ( 
.A(n_19546),
.Y(n_19642)
);

OAI22xp5_ASAP7_75t_L g19643 ( 
.A1(n_19400),
.A2(n_3688),
.B1(n_3686),
.B2(n_3687),
.Y(n_19643)
);

INVx1_ASAP7_75t_L g19644 ( 
.A(n_19388),
.Y(n_19644)
);

INVx1_ASAP7_75t_L g19645 ( 
.A(n_19498),
.Y(n_19645)
);

AOI221xp5_ASAP7_75t_L g19646 ( 
.A1(n_19516),
.A2(n_19574),
.B1(n_19583),
.B2(n_19509),
.C(n_19581),
.Y(n_19646)
);

OAI211xp5_ASAP7_75t_SL g19647 ( 
.A1(n_19446),
.A2(n_3689),
.B(n_3687),
.C(n_3688),
.Y(n_19647)
);

AO22x2_ASAP7_75t_L g19648 ( 
.A1(n_19511),
.A2(n_3692),
.B1(n_3690),
.B2(n_3691),
.Y(n_19648)
);

AOI22xp5_ASAP7_75t_L g19649 ( 
.A1(n_19382),
.A2(n_3693),
.B1(n_3690),
.B2(n_3692),
.Y(n_19649)
);

NAND2xp5_ASAP7_75t_L g19650 ( 
.A(n_19425),
.B(n_3693),
.Y(n_19650)
);

INVx2_ASAP7_75t_L g19651 ( 
.A(n_19588),
.Y(n_19651)
);

INVx1_ASAP7_75t_L g19652 ( 
.A(n_19513),
.Y(n_19652)
);

INVx2_ASAP7_75t_L g19653 ( 
.A(n_19472),
.Y(n_19653)
);

AO22x2_ASAP7_75t_L g19654 ( 
.A1(n_19529),
.A2(n_3696),
.B1(n_3694),
.B2(n_3695),
.Y(n_19654)
);

AOI22xp33_ASAP7_75t_SL g19655 ( 
.A1(n_19421),
.A2(n_3698),
.B1(n_3695),
.B2(n_3697),
.Y(n_19655)
);

AOI31xp33_ASAP7_75t_L g19656 ( 
.A1(n_19447),
.A2(n_3700),
.A3(n_3698),
.B(n_3699),
.Y(n_19656)
);

NAND2xp5_ASAP7_75t_L g19657 ( 
.A(n_19398),
.B(n_3699),
.Y(n_19657)
);

INVx1_ASAP7_75t_L g19658 ( 
.A(n_19515),
.Y(n_19658)
);

OAI22xp5_ASAP7_75t_L g19659 ( 
.A1(n_19386),
.A2(n_3702),
.B1(n_3700),
.B2(n_3701),
.Y(n_19659)
);

AO22x2_ASAP7_75t_L g19660 ( 
.A1(n_19578),
.A2(n_3703),
.B1(n_3701),
.B2(n_3702),
.Y(n_19660)
);

INVx1_ASAP7_75t_L g19661 ( 
.A(n_19526),
.Y(n_19661)
);

INVx1_ASAP7_75t_L g19662 ( 
.A(n_19527),
.Y(n_19662)
);

INVx1_ASAP7_75t_L g19663 ( 
.A(n_19538),
.Y(n_19663)
);

NOR2xp33_ASAP7_75t_SL g19664 ( 
.A(n_19457),
.B(n_3703),
.Y(n_19664)
);

AOI22xp5_ASAP7_75t_L g19665 ( 
.A1(n_19497),
.A2(n_3706),
.B1(n_3704),
.B2(n_3705),
.Y(n_19665)
);

INVx1_ASAP7_75t_L g19666 ( 
.A(n_19545),
.Y(n_19666)
);

NAND2xp5_ASAP7_75t_L g19667 ( 
.A(n_19507),
.B(n_19519),
.Y(n_19667)
);

AO22x1_ASAP7_75t_L g19668 ( 
.A1(n_19494),
.A2(n_3707),
.B1(n_3704),
.B2(n_3706),
.Y(n_19668)
);

AOI22xp5_ASAP7_75t_L g19669 ( 
.A1(n_19520),
.A2(n_3709),
.B1(n_3707),
.B2(n_3708),
.Y(n_19669)
);

INVx2_ASAP7_75t_L g19670 ( 
.A(n_19470),
.Y(n_19670)
);

INVx1_ASAP7_75t_L g19671 ( 
.A(n_19564),
.Y(n_19671)
);

INVx1_ASAP7_75t_L g19672 ( 
.A(n_19569),
.Y(n_19672)
);

NOR2x1_ASAP7_75t_L g19673 ( 
.A(n_19458),
.B(n_3708),
.Y(n_19673)
);

AOI22xp5_ASAP7_75t_L g19674 ( 
.A1(n_19540),
.A2(n_19556),
.B1(n_19573),
.B2(n_19572),
.Y(n_19674)
);

INVx1_ASAP7_75t_L g19675 ( 
.A(n_19407),
.Y(n_19675)
);

NAND2xp5_ASAP7_75t_L g19676 ( 
.A(n_19548),
.B(n_3709),
.Y(n_19676)
);

INVx1_ASAP7_75t_L g19677 ( 
.A(n_19415),
.Y(n_19677)
);

INVx1_ASAP7_75t_L g19678 ( 
.A(n_19440),
.Y(n_19678)
);

AOI22xp5_ASAP7_75t_L g19679 ( 
.A1(n_19576),
.A2(n_3712),
.B1(n_3710),
.B2(n_3711),
.Y(n_19679)
);

OA22x2_ASAP7_75t_L g19680 ( 
.A1(n_19500),
.A2(n_3712),
.B1(n_3710),
.B2(n_3711),
.Y(n_19680)
);

NOR2x1_ASAP7_75t_L g19681 ( 
.A(n_19437),
.B(n_3713),
.Y(n_19681)
);

NAND2xp5_ASAP7_75t_SL g19682 ( 
.A(n_19408),
.B(n_3713),
.Y(n_19682)
);

AOI22xp33_ASAP7_75t_L g19683 ( 
.A1(n_19482),
.A2(n_3716),
.B1(n_3714),
.B2(n_3715),
.Y(n_19683)
);

AOI22xp5_ASAP7_75t_L g19684 ( 
.A1(n_19587),
.A2(n_3716),
.B1(n_3714),
.B2(n_3715),
.Y(n_19684)
);

INVx1_ASAP7_75t_L g19685 ( 
.A(n_19452),
.Y(n_19685)
);

INVx1_ASAP7_75t_L g19686 ( 
.A(n_19479),
.Y(n_19686)
);

INVx1_ASAP7_75t_L g19687 ( 
.A(n_19433),
.Y(n_19687)
);

NAND4xp25_ASAP7_75t_SL g19688 ( 
.A(n_19568),
.B(n_3719),
.C(n_3717),
.D(n_3718),
.Y(n_19688)
);

INVx1_ASAP7_75t_L g19689 ( 
.A(n_19544),
.Y(n_19689)
);

NOR4xp25_ASAP7_75t_L g19690 ( 
.A(n_19460),
.B(n_3719),
.C(n_3717),
.D(n_3718),
.Y(n_19690)
);

NAND2xp5_ASAP7_75t_L g19691 ( 
.A(n_19402),
.B(n_3720),
.Y(n_19691)
);

OAI21xp5_ASAP7_75t_SL g19692 ( 
.A1(n_19501),
.A2(n_3720),
.B(n_3721),
.Y(n_19692)
);

NOR4xp25_ASAP7_75t_L g19693 ( 
.A(n_19428),
.B(n_3723),
.C(n_3721),
.D(n_3722),
.Y(n_19693)
);

HB1xp67_ASAP7_75t_L g19694 ( 
.A(n_19455),
.Y(n_19694)
);

AO22x1_ASAP7_75t_L g19695 ( 
.A1(n_19478),
.A2(n_3725),
.B1(n_3722),
.B2(n_3724),
.Y(n_19695)
);

AOI22xp5_ASAP7_75t_L g19696 ( 
.A1(n_19505),
.A2(n_3727),
.B1(n_3725),
.B2(n_3726),
.Y(n_19696)
);

NOR4xp25_ASAP7_75t_L g19697 ( 
.A(n_19585),
.B(n_3728),
.C(n_3726),
.D(n_3727),
.Y(n_19697)
);

NOR4xp25_ASAP7_75t_L g19698 ( 
.A(n_19438),
.B(n_3731),
.C(n_3728),
.D(n_3729),
.Y(n_19698)
);

NAND2xp5_ASAP7_75t_SL g19699 ( 
.A(n_19423),
.B(n_3729),
.Y(n_19699)
);

NOR2x1_ASAP7_75t_L g19700 ( 
.A(n_19471),
.B(n_3732),
.Y(n_19700)
);

AO22x2_ASAP7_75t_L g19701 ( 
.A1(n_19443),
.A2(n_3734),
.B1(n_3732),
.B2(n_3733),
.Y(n_19701)
);

INVx1_ASAP7_75t_L g19702 ( 
.A(n_19550),
.Y(n_19702)
);

AO22x1_ASAP7_75t_L g19703 ( 
.A1(n_19389),
.A2(n_3736),
.B1(n_3733),
.B2(n_3735),
.Y(n_19703)
);

AOI22xp5_ASAP7_75t_L g19704 ( 
.A1(n_19510),
.A2(n_19534),
.B1(n_19589),
.B2(n_19531),
.Y(n_19704)
);

NAND2xp5_ASAP7_75t_L g19705 ( 
.A(n_19466),
.B(n_3736),
.Y(n_19705)
);

AND2x4_ASAP7_75t_L g19706 ( 
.A(n_19535),
.B(n_3737),
.Y(n_19706)
);

AOI22xp5_ASAP7_75t_L g19707 ( 
.A1(n_19444),
.A2(n_3739),
.B1(n_3737),
.B2(n_3738),
.Y(n_19707)
);

INVx2_ASAP7_75t_L g19708 ( 
.A(n_19467),
.Y(n_19708)
);

AOI22xp5_ASAP7_75t_L g19709 ( 
.A1(n_19521),
.A2(n_3740),
.B1(n_3738),
.B2(n_3739),
.Y(n_19709)
);

AO22x2_ASAP7_75t_L g19710 ( 
.A1(n_19416),
.A2(n_3742),
.B1(n_3740),
.B2(n_3741),
.Y(n_19710)
);

OA22x2_ASAP7_75t_L g19711 ( 
.A1(n_19553),
.A2(n_3743),
.B1(n_3741),
.B2(n_3742),
.Y(n_19711)
);

OAI22xp5_ASAP7_75t_SL g19712 ( 
.A1(n_19449),
.A2(n_3745),
.B1(n_3743),
.B2(n_3744),
.Y(n_19712)
);

INVx1_ASAP7_75t_SL g19713 ( 
.A(n_19395),
.Y(n_19713)
);

INVx2_ASAP7_75t_L g19714 ( 
.A(n_19575),
.Y(n_19714)
);

NOR2xp33_ASAP7_75t_L g19715 ( 
.A(n_19488),
.B(n_3744),
.Y(n_19715)
);

INVx1_ASAP7_75t_L g19716 ( 
.A(n_19555),
.Y(n_19716)
);

NOR2x1_ASAP7_75t_L g19717 ( 
.A(n_19492),
.B(n_3745),
.Y(n_19717)
);

AO22x2_ASAP7_75t_L g19718 ( 
.A1(n_19418),
.A2(n_3748),
.B1(n_3746),
.B2(n_3747),
.Y(n_19718)
);

AOI22xp5_ASAP7_75t_L g19719 ( 
.A1(n_19522),
.A2(n_3749),
.B1(n_3747),
.B2(n_3748),
.Y(n_19719)
);

INVx1_ASAP7_75t_L g19720 ( 
.A(n_19559),
.Y(n_19720)
);

NOR4xp25_ASAP7_75t_L g19721 ( 
.A(n_19453),
.B(n_3751),
.C(n_3749),
.D(n_3750),
.Y(n_19721)
);

NAND2xp5_ASAP7_75t_L g19722 ( 
.A(n_19475),
.B(n_3750),
.Y(n_19722)
);

AOI22xp5_ASAP7_75t_L g19723 ( 
.A1(n_19530),
.A2(n_3753),
.B1(n_3751),
.B2(n_3752),
.Y(n_19723)
);

AOI22xp5_ASAP7_75t_L g19724 ( 
.A1(n_19541),
.A2(n_3754),
.B1(n_3752),
.B2(n_3753),
.Y(n_19724)
);

AOI22xp5_ASAP7_75t_L g19725 ( 
.A1(n_19562),
.A2(n_19566),
.B1(n_19561),
.B2(n_19563),
.Y(n_19725)
);

AOI221xp5_ASAP7_75t_L g19726 ( 
.A1(n_19392),
.A2(n_3756),
.B1(n_3754),
.B2(n_3755),
.C(n_3757),
.Y(n_19726)
);

NAND2xp5_ASAP7_75t_L g19727 ( 
.A(n_19401),
.B(n_3755),
.Y(n_19727)
);

AO22x2_ASAP7_75t_L g19728 ( 
.A1(n_19463),
.A2(n_3758),
.B1(n_3756),
.B2(n_3757),
.Y(n_19728)
);

OAI22xp5_ASAP7_75t_SL g19729 ( 
.A1(n_19580),
.A2(n_3760),
.B1(n_3758),
.B2(n_3759),
.Y(n_19729)
);

NAND2xp5_ASAP7_75t_SL g19730 ( 
.A(n_19484),
.B(n_3759),
.Y(n_19730)
);

AOI22xp5_ASAP7_75t_L g19731 ( 
.A1(n_19399),
.A2(n_3762),
.B1(n_3760),
.B2(n_3761),
.Y(n_19731)
);

OAI22xp5_ASAP7_75t_L g19732 ( 
.A1(n_19584),
.A2(n_3763),
.B1(n_3761),
.B2(n_3762),
.Y(n_19732)
);

NAND2xp5_ASAP7_75t_SL g19733 ( 
.A(n_19590),
.B(n_3763),
.Y(n_19733)
);

INVx1_ASAP7_75t_L g19734 ( 
.A(n_19445),
.Y(n_19734)
);

INVx2_ASAP7_75t_L g19735 ( 
.A(n_19422),
.Y(n_19735)
);

AOI22xp5_ASAP7_75t_L g19736 ( 
.A1(n_19567),
.A2(n_3766),
.B1(n_3764),
.B2(n_3765),
.Y(n_19736)
);

NAND2xp5_ASAP7_75t_L g19737 ( 
.A(n_19439),
.B(n_3764),
.Y(n_19737)
);

OA22x2_ASAP7_75t_SL g19738 ( 
.A1(n_19469),
.A2(n_19495),
.B1(n_19493),
.B2(n_19487),
.Y(n_19738)
);

INVx1_ASAP7_75t_L g19739 ( 
.A(n_19552),
.Y(n_19739)
);

NOR2x1_ASAP7_75t_L g19740 ( 
.A(n_19459),
.B(n_19512),
.Y(n_19740)
);

INVx1_ASAP7_75t_L g19741 ( 
.A(n_19430),
.Y(n_19741)
);

NAND2xp5_ASAP7_75t_L g19742 ( 
.A(n_19385),
.B(n_3767),
.Y(n_19742)
);

INVx1_ASAP7_75t_L g19743 ( 
.A(n_19419),
.Y(n_19743)
);

INVx1_ASAP7_75t_L g19744 ( 
.A(n_19403),
.Y(n_19744)
);

OAI211xp5_ASAP7_75t_L g19745 ( 
.A1(n_19429),
.A2(n_3769),
.B(n_3767),
.C(n_3768),
.Y(n_19745)
);

INVx1_ASAP7_75t_L g19746 ( 
.A(n_19448),
.Y(n_19746)
);

AO22x2_ASAP7_75t_L g19747 ( 
.A1(n_19532),
.A2(n_3771),
.B1(n_3769),
.B2(n_3770),
.Y(n_19747)
);

NAND2xp5_ASAP7_75t_L g19748 ( 
.A(n_19462),
.B(n_19483),
.Y(n_19748)
);

NAND2xp5_ASAP7_75t_SL g19749 ( 
.A(n_19582),
.B(n_19465),
.Y(n_19749)
);

INVxp67_ASAP7_75t_L g19750 ( 
.A(n_19474),
.Y(n_19750)
);

AOI22xp5_ASAP7_75t_L g19751 ( 
.A1(n_19586),
.A2(n_19431),
.B1(n_19503),
.B2(n_19417),
.Y(n_19751)
);

OR2x6_ASAP7_75t_L g19752 ( 
.A(n_19477),
.B(n_3770),
.Y(n_19752)
);

NOR4xp25_ASAP7_75t_L g19753 ( 
.A(n_19405),
.B(n_3774),
.C(n_3772),
.D(n_3773),
.Y(n_19753)
);

OAI22xp5_ASAP7_75t_L g19754 ( 
.A1(n_19517),
.A2(n_3777),
.B1(n_3775),
.B2(n_3776),
.Y(n_19754)
);

OAI22xp5_ASAP7_75t_SL g19755 ( 
.A1(n_19427),
.A2(n_19424),
.B1(n_19528),
.B2(n_19454),
.Y(n_19755)
);

INVx1_ASAP7_75t_L g19756 ( 
.A(n_19420),
.Y(n_19756)
);

INVx1_ASAP7_75t_L g19757 ( 
.A(n_19506),
.Y(n_19757)
);

AOI221xp5_ASAP7_75t_L g19758 ( 
.A1(n_19539),
.A2(n_19565),
.B1(n_19570),
.B2(n_19551),
.C(n_19473),
.Y(n_19758)
);

OR2x2_ASAP7_75t_L g19759 ( 
.A(n_19523),
.B(n_3775),
.Y(n_19759)
);

AO22x1_ASAP7_75t_L g19760 ( 
.A1(n_19489),
.A2(n_19525),
.B1(n_19518),
.B2(n_19486),
.Y(n_19760)
);

OAI22xp5_ASAP7_75t_L g19761 ( 
.A1(n_19485),
.A2(n_3778),
.B1(n_3776),
.B2(n_3777),
.Y(n_19761)
);

AOI22xp5_ASAP7_75t_L g19762 ( 
.A1(n_19542),
.A2(n_3781),
.B1(n_3779),
.B2(n_3780),
.Y(n_19762)
);

INVx2_ASAP7_75t_L g19763 ( 
.A(n_19480),
.Y(n_19763)
);

AOI22xp5_ASAP7_75t_L g19764 ( 
.A1(n_19387),
.A2(n_3781),
.B1(n_3779),
.B2(n_3780),
.Y(n_19764)
);

AOI22xp5_ASAP7_75t_L g19765 ( 
.A1(n_19387),
.A2(n_3784),
.B1(n_3782),
.B2(n_3783),
.Y(n_19765)
);

AOI22xp5_ASAP7_75t_L g19766 ( 
.A1(n_19387),
.A2(n_3784),
.B1(n_3782),
.B2(n_3783),
.Y(n_19766)
);

OA22x2_ASAP7_75t_L g19767 ( 
.A1(n_19393),
.A2(n_3787),
.B1(n_3785),
.B2(n_3786),
.Y(n_19767)
);

INVx1_ASAP7_75t_L g19768 ( 
.A(n_19625),
.Y(n_19768)
);

AOI21xp5_ASAP7_75t_L g19769 ( 
.A1(n_19598),
.A2(n_3788),
.B(n_3789),
.Y(n_19769)
);

INVx1_ASAP7_75t_L g19770 ( 
.A(n_19627),
.Y(n_19770)
);

NAND2xp5_ASAP7_75t_L g19771 ( 
.A(n_19604),
.B(n_3788),
.Y(n_19771)
);

INVx1_ASAP7_75t_L g19772 ( 
.A(n_19680),
.Y(n_19772)
);

NOR3xp33_ASAP7_75t_L g19773 ( 
.A(n_19599),
.B(n_3789),
.C(n_3790),
.Y(n_19773)
);

INVx1_ASAP7_75t_L g19774 ( 
.A(n_19711),
.Y(n_19774)
);

NAND2xp5_ASAP7_75t_SL g19775 ( 
.A(n_19693),
.B(n_3790),
.Y(n_19775)
);

INVx1_ASAP7_75t_L g19776 ( 
.A(n_19767),
.Y(n_19776)
);

OAI21xp5_ASAP7_75t_L g19777 ( 
.A1(n_19601),
.A2(n_3791),
.B(n_3792),
.Y(n_19777)
);

NAND2xp5_ASAP7_75t_L g19778 ( 
.A(n_19695),
.B(n_3791),
.Y(n_19778)
);

NAND2xp5_ASAP7_75t_L g19779 ( 
.A(n_19668),
.B(n_3792),
.Y(n_19779)
);

OAI21xp33_ASAP7_75t_SL g19780 ( 
.A1(n_19610),
.A2(n_19623),
.B(n_19620),
.Y(n_19780)
);

AND2x2_ASAP7_75t_L g19781 ( 
.A(n_19626),
.B(n_3793),
.Y(n_19781)
);

AND2x2_ASAP7_75t_L g19782 ( 
.A(n_19706),
.B(n_19600),
.Y(n_19782)
);

INVx1_ASAP7_75t_L g19783 ( 
.A(n_19691),
.Y(n_19783)
);

INVx2_ASAP7_75t_L g19784 ( 
.A(n_19752),
.Y(n_19784)
);

INVx2_ASAP7_75t_SL g19785 ( 
.A(n_19717),
.Y(n_19785)
);

NAND3xp33_ASAP7_75t_L g19786 ( 
.A(n_19758),
.B(n_3793),
.C(n_3795),
.Y(n_19786)
);

INVx2_ASAP7_75t_L g19787 ( 
.A(n_19752),
.Y(n_19787)
);

INVx2_ASAP7_75t_SL g19788 ( 
.A(n_19673),
.Y(n_19788)
);

NAND3x1_ASAP7_75t_SL g19789 ( 
.A(n_19681),
.B(n_3795),
.C(n_3796),
.Y(n_19789)
);

NOR2x1p5_ASAP7_75t_L g19790 ( 
.A(n_19628),
.B(n_3796),
.Y(n_19790)
);

NOR3xp33_ASAP7_75t_SL g19791 ( 
.A(n_19618),
.B(n_3797),
.C(n_3798),
.Y(n_19791)
);

NAND3xp33_ASAP7_75t_L g19792 ( 
.A(n_19726),
.B(n_3797),
.C(n_3798),
.Y(n_19792)
);

NAND2xp5_ASAP7_75t_L g19793 ( 
.A(n_19703),
.B(n_3799),
.Y(n_19793)
);

INVx1_ASAP7_75t_L g19794 ( 
.A(n_19747),
.Y(n_19794)
);

HB1xp67_ASAP7_75t_L g19795 ( 
.A(n_19747),
.Y(n_19795)
);

NAND2xp5_ASAP7_75t_L g19796 ( 
.A(n_19606),
.B(n_3799),
.Y(n_19796)
);

AOI221xp5_ASAP7_75t_L g19797 ( 
.A1(n_19631),
.A2(n_3802),
.B1(n_3800),
.B2(n_3801),
.C(n_3803),
.Y(n_19797)
);

INVx1_ASAP7_75t_L g19798 ( 
.A(n_19729),
.Y(n_19798)
);

NOR2x1_ASAP7_75t_L g19799 ( 
.A(n_19605),
.B(n_3801),
.Y(n_19799)
);

INVx2_ASAP7_75t_L g19800 ( 
.A(n_19619),
.Y(n_19800)
);

AND2x2_ASAP7_75t_L g19801 ( 
.A(n_19591),
.B(n_3803),
.Y(n_19801)
);

NAND2xp5_ASAP7_75t_L g19802 ( 
.A(n_19608),
.B(n_3804),
.Y(n_19802)
);

OR2x2_ASAP7_75t_L g19803 ( 
.A(n_19698),
.B(n_3804),
.Y(n_19803)
);

NOR2x1_ASAP7_75t_L g19804 ( 
.A(n_19609),
.B(n_19603),
.Y(n_19804)
);

NAND2xp5_ASAP7_75t_L g19805 ( 
.A(n_19613),
.B(n_3805),
.Y(n_19805)
);

AND2x2_ASAP7_75t_L g19806 ( 
.A(n_19715),
.B(n_3805),
.Y(n_19806)
);

NAND2xp5_ASAP7_75t_L g19807 ( 
.A(n_19655),
.B(n_3806),
.Y(n_19807)
);

NAND2xp5_ASAP7_75t_L g19808 ( 
.A(n_19736),
.B(n_3806),
.Y(n_19808)
);

AND2x2_ASAP7_75t_L g19809 ( 
.A(n_19607),
.B(n_3807),
.Y(n_19809)
);

NAND2xp5_ASAP7_75t_L g19810 ( 
.A(n_19707),
.B(n_3807),
.Y(n_19810)
);

NOR3xp33_ASAP7_75t_L g19811 ( 
.A(n_19639),
.B(n_3808),
.C(n_3809),
.Y(n_19811)
);

NAND2xp5_ASAP7_75t_SL g19812 ( 
.A(n_19690),
.B(n_19709),
.Y(n_19812)
);

OAI221xp5_ASAP7_75t_L g19813 ( 
.A1(n_19731),
.A2(n_3810),
.B1(n_3808),
.B2(n_3809),
.C(n_3811),
.Y(n_19813)
);

NAND2xp5_ASAP7_75t_L g19814 ( 
.A(n_19760),
.B(n_3810),
.Y(n_19814)
);

AND2x4_ASAP7_75t_L g19815 ( 
.A(n_19617),
.B(n_19597),
.Y(n_19815)
);

INVx2_ASAP7_75t_L g19816 ( 
.A(n_19619),
.Y(n_19816)
);

NAND2xp5_ASAP7_75t_L g19817 ( 
.A(n_19719),
.B(n_3812),
.Y(n_19817)
);

AND2x2_ASAP7_75t_L g19818 ( 
.A(n_19763),
.B(n_3813),
.Y(n_19818)
);

NAND2xp5_ASAP7_75t_L g19819 ( 
.A(n_19723),
.B(n_3813),
.Y(n_19819)
);

OAI21xp5_ASAP7_75t_L g19820 ( 
.A1(n_19692),
.A2(n_3814),
.B(n_3815),
.Y(n_19820)
);

O2A1O1Ixp5_ASAP7_75t_L g19821 ( 
.A1(n_19638),
.A2(n_3817),
.B(n_3814),
.C(n_3816),
.Y(n_19821)
);

INVx1_ASAP7_75t_L g19822 ( 
.A(n_19712),
.Y(n_19822)
);

INVx3_ASAP7_75t_L g19823 ( 
.A(n_19621),
.Y(n_19823)
);

INVx1_ASAP7_75t_L g19824 ( 
.A(n_19759),
.Y(n_19824)
);

NOR2xp33_ASAP7_75t_L g19825 ( 
.A(n_19664),
.B(n_3816),
.Y(n_19825)
);

NAND2xp5_ASAP7_75t_L g19826 ( 
.A(n_19724),
.B(n_3817),
.Y(n_19826)
);

NOR2xp67_ASAP7_75t_SL g19827 ( 
.A(n_19611),
.B(n_19612),
.Y(n_19827)
);

INVx1_ASAP7_75t_L g19828 ( 
.A(n_19722),
.Y(n_19828)
);

NOR2x1p5_ASAP7_75t_L g19829 ( 
.A(n_19595),
.B(n_3818),
.Y(n_19829)
);

HB1xp67_ASAP7_75t_L g19830 ( 
.A(n_19697),
.Y(n_19830)
);

INVx1_ASAP7_75t_L g19831 ( 
.A(n_19737),
.Y(n_19831)
);

NAND3xp33_ASAP7_75t_L g19832 ( 
.A(n_19615),
.B(n_3818),
.C(n_3819),
.Y(n_19832)
);

AOI221xp5_ASAP7_75t_L g19833 ( 
.A1(n_19754),
.A2(n_3821),
.B1(n_3819),
.B2(n_3820),
.C(n_3822),
.Y(n_19833)
);

NAND2xp33_ASAP7_75t_L g19834 ( 
.A(n_19596),
.B(n_3820),
.Y(n_19834)
);

NAND2xp5_ASAP7_75t_L g19835 ( 
.A(n_19649),
.B(n_3821),
.Y(n_19835)
);

NAND2xp5_ASAP7_75t_L g19836 ( 
.A(n_19665),
.B(n_3822),
.Y(n_19836)
);

AND4x2_ASAP7_75t_L g19837 ( 
.A(n_19700),
.B(n_3825),
.C(n_3823),
.D(n_3824),
.Y(n_19837)
);

NAND2xp5_ASAP7_75t_L g19838 ( 
.A(n_19669),
.B(n_3823),
.Y(n_19838)
);

INVx1_ASAP7_75t_L g19839 ( 
.A(n_19742),
.Y(n_19839)
);

AND2x2_ASAP7_75t_L g19840 ( 
.A(n_19694),
.B(n_3825),
.Y(n_19840)
);

AOI21xp5_ASAP7_75t_L g19841 ( 
.A1(n_19749),
.A2(n_3826),
.B(n_3827),
.Y(n_19841)
);

NOR2xp33_ASAP7_75t_L g19842 ( 
.A(n_19688),
.B(n_3827),
.Y(n_19842)
);

NOR2x1_ASAP7_75t_L g19843 ( 
.A(n_19616),
.B(n_3828),
.Y(n_19843)
);

INVx1_ASAP7_75t_L g19844 ( 
.A(n_19650),
.Y(n_19844)
);

NAND2xp5_ASAP7_75t_SL g19845 ( 
.A(n_19753),
.B(n_3828),
.Y(n_19845)
);

NAND2xp5_ASAP7_75t_L g19846 ( 
.A(n_19679),
.B(n_3829),
.Y(n_19846)
);

INVx4_ASAP7_75t_L g19847 ( 
.A(n_19622),
.Y(n_19847)
);

INVx1_ASAP7_75t_SL g19848 ( 
.A(n_19593),
.Y(n_19848)
);

XOR2x2_ASAP7_75t_L g19849 ( 
.A(n_19640),
.B(n_3829),
.Y(n_19849)
);

NAND2xp5_ASAP7_75t_L g19850 ( 
.A(n_19684),
.B(n_19762),
.Y(n_19850)
);

NOR2xp33_ASAP7_75t_L g19851 ( 
.A(n_19705),
.B(n_3830),
.Y(n_19851)
);

INVx2_ASAP7_75t_L g19852 ( 
.A(n_19648),
.Y(n_19852)
);

OAI322xp33_ASAP7_75t_L g19853 ( 
.A1(n_19738),
.A2(n_3836),
.A3(n_3835),
.B1(n_3832),
.B2(n_3830),
.C1(n_3831),
.C2(n_3833),
.Y(n_19853)
);

AND3x1_ASAP7_75t_L g19854 ( 
.A(n_19630),
.B(n_3831),
.C(n_3832),
.Y(n_19854)
);

INVx1_ASAP7_75t_L g19855 ( 
.A(n_19727),
.Y(n_19855)
);

OR2x2_ASAP7_75t_L g19856 ( 
.A(n_19721),
.B(n_3833),
.Y(n_19856)
);

NAND2xp5_ASAP7_75t_L g19857 ( 
.A(n_19643),
.B(n_19592),
.Y(n_19857)
);

INVx1_ASAP7_75t_L g19858 ( 
.A(n_19676),
.Y(n_19858)
);

AOI211xp5_ASAP7_75t_L g19859 ( 
.A1(n_19659),
.A2(n_3838),
.B(n_3836),
.C(n_3837),
.Y(n_19859)
);

NAND2xp5_ASAP7_75t_L g19860 ( 
.A(n_19732),
.B(n_3837),
.Y(n_19860)
);

AND2x2_ASAP7_75t_L g19861 ( 
.A(n_19743),
.B(n_3838),
.Y(n_19861)
);

AND2x2_ASAP7_75t_L g19862 ( 
.A(n_19642),
.B(n_3839),
.Y(n_19862)
);

BUFx12f_ASAP7_75t_L g19863 ( 
.A(n_19713),
.Y(n_19863)
);

INVx1_ASAP7_75t_L g19864 ( 
.A(n_19657),
.Y(n_19864)
);

OAI21xp33_ASAP7_75t_SL g19865 ( 
.A1(n_19646),
.A2(n_3839),
.B(n_3840),
.Y(n_19865)
);

NOR2x1_ASAP7_75t_L g19866 ( 
.A(n_19624),
.B(n_3840),
.Y(n_19866)
);

NOR2xp33_ASAP7_75t_L g19867 ( 
.A(n_19730),
.B(n_3841),
.Y(n_19867)
);

INVx1_ASAP7_75t_L g19868 ( 
.A(n_19745),
.Y(n_19868)
);

INVx1_ASAP7_75t_L g19869 ( 
.A(n_19634),
.Y(n_19869)
);

NAND2xp5_ASAP7_75t_L g19870 ( 
.A(n_19632),
.B(n_3841),
.Y(n_19870)
);

NAND2xp5_ASAP7_75t_L g19871 ( 
.A(n_19696),
.B(n_3842),
.Y(n_19871)
);

NAND2xp5_ASAP7_75t_L g19872 ( 
.A(n_19594),
.B(n_3842),
.Y(n_19872)
);

XOR2x2_ASAP7_75t_L g19873 ( 
.A(n_19740),
.B(n_3843),
.Y(n_19873)
);

INVx1_ASAP7_75t_L g19874 ( 
.A(n_19733),
.Y(n_19874)
);

NAND2xp5_ASAP7_75t_L g19875 ( 
.A(n_19683),
.B(n_3843),
.Y(n_19875)
);

INVx1_ASAP7_75t_L g19876 ( 
.A(n_19648),
.Y(n_19876)
);

NAND2xp5_ASAP7_75t_L g19877 ( 
.A(n_19725),
.B(n_3844),
.Y(n_19877)
);

NAND2xp5_ASAP7_75t_L g19878 ( 
.A(n_19761),
.B(n_3844),
.Y(n_19878)
);

NAND2xp5_ASAP7_75t_L g19879 ( 
.A(n_19686),
.B(n_3845),
.Y(n_19879)
);

INVx1_ASAP7_75t_L g19880 ( 
.A(n_19654),
.Y(n_19880)
);

NAND2xp5_ASAP7_75t_L g19881 ( 
.A(n_19678),
.B(n_3845),
.Y(n_19881)
);

XNOR2xp5_ASAP7_75t_L g19882 ( 
.A(n_19751),
.B(n_3846),
.Y(n_19882)
);

INVxp67_ASAP7_75t_L g19883 ( 
.A(n_19651),
.Y(n_19883)
);

INVx5_ASAP7_75t_L g19884 ( 
.A(n_19714),
.Y(n_19884)
);

NOR2x1p5_ASAP7_75t_L g19885 ( 
.A(n_19748),
.B(n_19667),
.Y(n_19885)
);

INVx2_ASAP7_75t_SL g19886 ( 
.A(n_19735),
.Y(n_19886)
);

NAND2x1p5_ASAP7_75t_L g19887 ( 
.A(n_19685),
.B(n_3846),
.Y(n_19887)
);

NAND2xp33_ASAP7_75t_L g19888 ( 
.A(n_19739),
.B(n_3847),
.Y(n_19888)
);

INVx1_ASAP7_75t_L g19889 ( 
.A(n_19654),
.Y(n_19889)
);

INVx2_ASAP7_75t_SL g19890 ( 
.A(n_19660),
.Y(n_19890)
);

INVx1_ASAP7_75t_L g19891 ( 
.A(n_19660),
.Y(n_19891)
);

BUFx2_ASAP7_75t_L g19892 ( 
.A(n_19744),
.Y(n_19892)
);

OAI22xp33_ASAP7_75t_L g19893 ( 
.A1(n_19674),
.A2(n_3849),
.B1(n_3847),
.B2(n_3848),
.Y(n_19893)
);

INVx1_ASAP7_75t_L g19894 ( 
.A(n_19647),
.Y(n_19894)
);

NAND2xp5_ASAP7_75t_L g19895 ( 
.A(n_19602),
.B(n_3848),
.Y(n_19895)
);

NOR2x1_ASAP7_75t_L g19896 ( 
.A(n_19746),
.B(n_3850),
.Y(n_19896)
);

AO21x1_ASAP7_75t_L g19897 ( 
.A1(n_19734),
.A2(n_19702),
.B(n_19689),
.Y(n_19897)
);

NAND3xp33_ASAP7_75t_L g19898 ( 
.A(n_19716),
.B(n_3850),
.C(n_3851),
.Y(n_19898)
);

NAND3xp33_ASAP7_75t_L g19899 ( 
.A(n_19720),
.B(n_3851),
.C(n_3852),
.Y(n_19899)
);

NAND2xp5_ASAP7_75t_L g19900 ( 
.A(n_19764),
.B(n_19765),
.Y(n_19900)
);

NAND2xp5_ASAP7_75t_L g19901 ( 
.A(n_19766),
.B(n_3852),
.Y(n_19901)
);

INVx1_ASAP7_75t_SL g19902 ( 
.A(n_19682),
.Y(n_19902)
);

BUFx12f_ASAP7_75t_L g19903 ( 
.A(n_19863),
.Y(n_19903)
);

NAND2xp5_ASAP7_75t_L g19904 ( 
.A(n_19781),
.B(n_19675),
.Y(n_19904)
);

AOI22xp33_ASAP7_75t_L g19905 ( 
.A1(n_19809),
.A2(n_19653),
.B1(n_19670),
.B2(n_19708),
.Y(n_19905)
);

OAI211xp5_ASAP7_75t_L g19906 ( 
.A1(n_19814),
.A2(n_19750),
.B(n_19704),
.C(n_19756),
.Y(n_19906)
);

INVx1_ASAP7_75t_L g19907 ( 
.A(n_19837),
.Y(n_19907)
);

NAND2xp5_ASAP7_75t_L g19908 ( 
.A(n_19818),
.B(n_19633),
.Y(n_19908)
);

OAI21xp5_ASAP7_75t_SL g19909 ( 
.A1(n_19861),
.A2(n_19840),
.B(n_19862),
.Y(n_19909)
);

OAI22xp33_ASAP7_75t_L g19910 ( 
.A1(n_19877),
.A2(n_19757),
.B1(n_19637),
.B2(n_19635),
.Y(n_19910)
);

AND2x4_ASAP7_75t_L g19911 ( 
.A(n_19790),
.B(n_19629),
.Y(n_19911)
);

AOI321xp33_ASAP7_75t_L g19912 ( 
.A1(n_19804),
.A2(n_19699),
.A3(n_19687),
.B1(n_19741),
.B2(n_19644),
.C(n_19652),
.Y(n_19912)
);

OAI22xp33_ASAP7_75t_L g19913 ( 
.A1(n_19779),
.A2(n_19636),
.B1(n_19656),
.B2(n_19645),
.Y(n_19913)
);

AND2x4_ASAP7_75t_L g19914 ( 
.A(n_19829),
.B(n_19658),
.Y(n_19914)
);

NAND4xp75_ASAP7_75t_L g19915 ( 
.A(n_19897),
.B(n_19886),
.C(n_19780),
.D(n_19782),
.Y(n_19915)
);

AOI222xp33_ASAP7_75t_L g19916 ( 
.A1(n_19834),
.A2(n_19755),
.B1(n_19662),
.B2(n_19663),
.C1(n_19671),
.C2(n_19666),
.Y(n_19916)
);

A2O1A1Ixp33_ASAP7_75t_L g19917 ( 
.A1(n_19842),
.A2(n_19641),
.B(n_19672),
.C(n_19661),
.Y(n_19917)
);

O2A1O1Ixp33_ASAP7_75t_L g19918 ( 
.A1(n_19795),
.A2(n_19677),
.B(n_19614),
.C(n_19710),
.Y(n_19918)
);

OAI22xp5_ASAP7_75t_L g19919 ( 
.A1(n_19854),
.A2(n_19710),
.B1(n_19718),
.B2(n_19701),
.Y(n_19919)
);

AOI211xp5_ASAP7_75t_L g19920 ( 
.A1(n_19865),
.A2(n_19718),
.B(n_19701),
.C(n_19728),
.Y(n_19920)
);

NAND2xp5_ASAP7_75t_L g19921 ( 
.A(n_19896),
.B(n_19728),
.Y(n_19921)
);

AOI221x1_ASAP7_75t_L g19922 ( 
.A1(n_19794),
.A2(n_19768),
.B1(n_19880),
.B2(n_19889),
.C(n_19876),
.Y(n_19922)
);

OAI322xp33_ASAP7_75t_L g19923 ( 
.A1(n_19778),
.A2(n_3858),
.A3(n_3857),
.B1(n_3855),
.B2(n_3853),
.C1(n_3854),
.C2(n_3856),
.Y(n_19923)
);

NAND3x1_ASAP7_75t_L g19924 ( 
.A(n_19799),
.B(n_3854),
.C(n_3856),
.Y(n_19924)
);

NOR2x1_ASAP7_75t_L g19925 ( 
.A(n_19891),
.B(n_3857),
.Y(n_19925)
);

AOI211xp5_ASAP7_75t_L g19926 ( 
.A1(n_19867),
.A2(n_3860),
.B(n_3858),
.C(n_3859),
.Y(n_19926)
);

AOI221xp5_ASAP7_75t_L g19927 ( 
.A1(n_19797),
.A2(n_3861),
.B1(n_3859),
.B2(n_3860),
.C(n_3862),
.Y(n_19927)
);

INVx2_ASAP7_75t_SL g19928 ( 
.A(n_19887),
.Y(n_19928)
);

NAND2xp5_ASAP7_75t_SL g19929 ( 
.A(n_19833),
.B(n_3861),
.Y(n_19929)
);

NAND2xp5_ASAP7_75t_L g19930 ( 
.A(n_19882),
.B(n_3862),
.Y(n_19930)
);

NOR2xp33_ASAP7_75t_R g19931 ( 
.A(n_19890),
.B(n_3863),
.Y(n_19931)
);

NOR4xp25_ASAP7_75t_L g19932 ( 
.A(n_19883),
.B(n_3866),
.C(n_3864),
.D(n_3865),
.Y(n_19932)
);

AOI321xp33_ASAP7_75t_L g19933 ( 
.A1(n_19825),
.A2(n_3867),
.A3(n_3869),
.B1(n_3864),
.B2(n_3866),
.C(n_3868),
.Y(n_19933)
);

AND2x2_ASAP7_75t_L g19934 ( 
.A(n_19791),
.B(n_3867),
.Y(n_19934)
);

OAI321xp33_ASAP7_75t_L g19935 ( 
.A1(n_19820),
.A2(n_19793),
.A3(n_19771),
.B1(n_19808),
.B2(n_19792),
.C(n_19895),
.Y(n_19935)
);

OAI21xp5_ASAP7_75t_L g19936 ( 
.A1(n_19821),
.A2(n_3868),
.B(n_3870),
.Y(n_19936)
);

NAND2xp5_ASAP7_75t_L g19937 ( 
.A(n_19801),
.B(n_3870),
.Y(n_19937)
);

NAND2xp5_ASAP7_75t_SL g19938 ( 
.A(n_19884),
.B(n_3871),
.Y(n_19938)
);

OAI211xp5_ASAP7_75t_L g19939 ( 
.A1(n_19830),
.A2(n_3873),
.B(n_3871),
.C(n_3872),
.Y(n_19939)
);

NOR2xp33_ASAP7_75t_L g19940 ( 
.A(n_19803),
.B(n_3872),
.Y(n_19940)
);

OAI22xp33_ASAP7_75t_L g19941 ( 
.A1(n_19813),
.A2(n_3875),
.B1(n_3873),
.B2(n_3874),
.Y(n_19941)
);

AOI211xp5_ASAP7_75t_L g19942 ( 
.A1(n_19888),
.A2(n_3878),
.B(n_3876),
.C(n_3877),
.Y(n_19942)
);

HB1xp67_ASAP7_75t_L g19943 ( 
.A(n_19843),
.Y(n_19943)
);

NOR2xp67_ASAP7_75t_L g19944 ( 
.A(n_19856),
.B(n_3876),
.Y(n_19944)
);

NAND2xp5_ASAP7_75t_L g19945 ( 
.A(n_19806),
.B(n_3877),
.Y(n_19945)
);

INVx1_ASAP7_75t_SL g19946 ( 
.A(n_19879),
.Y(n_19946)
);

NOR2x1p5_ASAP7_75t_L g19947 ( 
.A(n_19807),
.B(n_3878),
.Y(n_19947)
);

AOI22xp5_ASAP7_75t_L g19948 ( 
.A1(n_19827),
.A2(n_3881),
.B1(n_3879),
.B2(n_3880),
.Y(n_19948)
);

NAND2xp5_ASAP7_75t_SL g19949 ( 
.A(n_19884),
.B(n_3879),
.Y(n_19949)
);

AND2x4_ASAP7_75t_L g19950 ( 
.A(n_19800),
.B(n_3880),
.Y(n_19950)
);

OAI221xp5_ASAP7_75t_SL g19951 ( 
.A1(n_19875),
.A2(n_3883),
.B1(n_3881),
.B2(n_3882),
.C(n_3884),
.Y(n_19951)
);

OAI22xp33_ASAP7_75t_L g19952 ( 
.A1(n_19847),
.A2(n_3884),
.B1(n_3882),
.B2(n_3883),
.Y(n_19952)
);

OAI211xp5_ASAP7_75t_L g19953 ( 
.A1(n_19777),
.A2(n_3887),
.B(n_3885),
.C(n_3886),
.Y(n_19953)
);

NAND2xp5_ASAP7_75t_L g19954 ( 
.A(n_19866),
.B(n_3885),
.Y(n_19954)
);

AOI221xp5_ASAP7_75t_L g19955 ( 
.A1(n_19775),
.A2(n_3888),
.B1(n_3886),
.B2(n_3887),
.C(n_3889),
.Y(n_19955)
);

A2O1A1Ixp33_ASAP7_75t_SL g19956 ( 
.A1(n_19823),
.A2(n_3890),
.B(n_3888),
.C(n_3889),
.Y(n_19956)
);

NAND4xp25_ASAP7_75t_L g19957 ( 
.A(n_19859),
.B(n_19892),
.C(n_19819),
.D(n_19826),
.Y(n_19957)
);

NAND3xp33_ASAP7_75t_L g19958 ( 
.A(n_19884),
.B(n_3890),
.C(n_3891),
.Y(n_19958)
);

INVx1_ASAP7_75t_L g19959 ( 
.A(n_19873),
.Y(n_19959)
);

AOI222xp33_ASAP7_75t_L g19960 ( 
.A1(n_19845),
.A2(n_3893),
.B1(n_3895),
.B2(n_3891),
.C1(n_3892),
.C2(n_3894),
.Y(n_19960)
);

NAND3xp33_ASAP7_75t_L g19961 ( 
.A(n_19851),
.B(n_3892),
.C(n_3896),
.Y(n_19961)
);

AOI22xp5_ASAP7_75t_L g19962 ( 
.A1(n_19849),
.A2(n_3899),
.B1(n_3897),
.B2(n_3898),
.Y(n_19962)
);

AOI22xp33_ASAP7_75t_L g19963 ( 
.A1(n_19788),
.A2(n_19787),
.B1(n_19784),
.B2(n_19785),
.Y(n_19963)
);

NAND3xp33_ASAP7_75t_SL g19964 ( 
.A(n_19902),
.B(n_3897),
.C(n_3898),
.Y(n_19964)
);

NAND2xp5_ASAP7_75t_L g19965 ( 
.A(n_19881),
.B(n_3899),
.Y(n_19965)
);

NOR3xp33_ASAP7_75t_L g19966 ( 
.A(n_19798),
.B(n_3900),
.C(n_3901),
.Y(n_19966)
);

OR2x2_ASAP7_75t_L g19967 ( 
.A(n_19796),
.B(n_3900),
.Y(n_19967)
);

XOR2xp5_ASAP7_75t_L g19968 ( 
.A(n_19783),
.B(n_3901),
.Y(n_19968)
);

INVx1_ASAP7_75t_L g19969 ( 
.A(n_19789),
.Y(n_19969)
);

AOI221xp5_ASAP7_75t_L g19970 ( 
.A1(n_19770),
.A2(n_3904),
.B1(n_3902),
.B2(n_3903),
.C(n_3905),
.Y(n_19970)
);

AOI221xp5_ASAP7_75t_L g19971 ( 
.A1(n_19772),
.A2(n_3905),
.B1(n_3902),
.B2(n_3903),
.C(n_3906),
.Y(n_19971)
);

NAND4xp75_ASAP7_75t_L g19972 ( 
.A(n_19774),
.B(n_3908),
.C(n_3906),
.D(n_3907),
.Y(n_19972)
);

INVx1_ASAP7_75t_SL g19973 ( 
.A(n_19860),
.Y(n_19973)
);

NAND2xp5_ASAP7_75t_L g19974 ( 
.A(n_19841),
.B(n_3907),
.Y(n_19974)
);

NOR2x1p5_ASAP7_75t_L g19975 ( 
.A(n_19817),
.B(n_19776),
.Y(n_19975)
);

AOI222xp33_ASAP7_75t_L g19976 ( 
.A1(n_19901),
.A2(n_3910),
.B1(n_3912),
.B2(n_3908),
.C1(n_3909),
.C2(n_3911),
.Y(n_19976)
);

INVx1_ASAP7_75t_L g19977 ( 
.A(n_19802),
.Y(n_19977)
);

OR2x2_ASAP7_75t_L g19978 ( 
.A(n_19805),
.B(n_3910),
.Y(n_19978)
);

OAI22xp33_ASAP7_75t_L g19979 ( 
.A1(n_19872),
.A2(n_3914),
.B1(n_3912),
.B2(n_3913),
.Y(n_19979)
);

AOI21xp5_ASAP7_75t_L g19980 ( 
.A1(n_19812),
.A2(n_3913),
.B(n_3914),
.Y(n_19980)
);

AOI33xp33_ASAP7_75t_L g19981 ( 
.A1(n_19894),
.A2(n_3917),
.A3(n_3919),
.B1(n_3915),
.B2(n_3916),
.B3(n_3918),
.Y(n_19981)
);

AOI22xp33_ASAP7_75t_L g19982 ( 
.A1(n_19815),
.A2(n_3917),
.B1(n_3915),
.B2(n_3916),
.Y(n_19982)
);

AOI221x1_ASAP7_75t_L g19983 ( 
.A1(n_19822),
.A2(n_3921),
.B1(n_3918),
.B2(n_3920),
.C(n_3922),
.Y(n_19983)
);

NAND3xp33_ASAP7_75t_SL g19984 ( 
.A(n_19848),
.B(n_3920),
.C(n_3921),
.Y(n_19984)
);

AOI22xp33_ASAP7_75t_L g19985 ( 
.A1(n_19815),
.A2(n_19869),
.B1(n_19868),
.B2(n_19824),
.Y(n_19985)
);

NAND2xp33_ASAP7_75t_SL g19986 ( 
.A(n_19878),
.B(n_3923),
.Y(n_19986)
);

AOI21xp33_ASAP7_75t_SL g19987 ( 
.A1(n_19811),
.A2(n_3923),
.B(n_3924),
.Y(n_19987)
);

OAI221xp5_ASAP7_75t_L g19988 ( 
.A1(n_19870),
.A2(n_3927),
.B1(n_3925),
.B2(n_3926),
.C(n_3928),
.Y(n_19988)
);

INVx1_ASAP7_75t_L g19989 ( 
.A(n_19810),
.Y(n_19989)
);

OAI21xp5_ASAP7_75t_L g19990 ( 
.A1(n_19835),
.A2(n_3926),
.B(n_3927),
.Y(n_19990)
);

NOR3xp33_ASAP7_75t_L g19991 ( 
.A(n_19874),
.B(n_3928),
.C(n_3929),
.Y(n_19991)
);

INVx1_ASAP7_75t_SL g19992 ( 
.A(n_19816),
.Y(n_19992)
);

NAND3xp33_ASAP7_75t_L g19993 ( 
.A(n_19852),
.B(n_3929),
.C(n_3930),
.Y(n_19993)
);

NAND4xp25_ASAP7_75t_L g19994 ( 
.A(n_19850),
.B(n_3932),
.C(n_3930),
.D(n_3931),
.Y(n_19994)
);

OR5x1_ASAP7_75t_L g19995 ( 
.A(n_19906),
.B(n_19885),
.C(n_19857),
.D(n_19900),
.E(n_19836),
.Y(n_19995)
);

AND4x1_ASAP7_75t_L g19996 ( 
.A(n_19922),
.B(n_19864),
.C(n_19858),
.D(n_19831),
.Y(n_19996)
);

OR2x2_ASAP7_75t_L g19997 ( 
.A(n_19930),
.B(n_19838),
.Y(n_19997)
);

AND2x4_ASAP7_75t_L g19998 ( 
.A(n_19944),
.B(n_19871),
.Y(n_19998)
);

OA21x2_ASAP7_75t_L g19999 ( 
.A1(n_19915),
.A2(n_19855),
.B(n_19839),
.Y(n_19999)
);

NOR2xp33_ASAP7_75t_L g20000 ( 
.A(n_19940),
.B(n_19846),
.Y(n_20000)
);

INVxp67_ASAP7_75t_SL g20001 ( 
.A(n_19925),
.Y(n_20001)
);

NAND2xp5_ASAP7_75t_L g20002 ( 
.A(n_19942),
.B(n_19769),
.Y(n_20002)
);

NAND3xp33_ASAP7_75t_L g20003 ( 
.A(n_19912),
.B(n_19844),
.C(n_19828),
.Y(n_20003)
);

NOR2x1_ASAP7_75t_L g20004 ( 
.A(n_19969),
.B(n_19786),
.Y(n_20004)
);

CKINVDCx5p33_ASAP7_75t_R g20005 ( 
.A(n_19903),
.Y(n_20005)
);

OAI22xp5_ASAP7_75t_L g20006 ( 
.A1(n_19962),
.A2(n_19899),
.B1(n_19898),
.B2(n_19832),
.Y(n_20006)
);

AND2x2_ASAP7_75t_L g20007 ( 
.A(n_19934),
.B(n_19773),
.Y(n_20007)
);

NAND3xp33_ASAP7_75t_L g20008 ( 
.A(n_19963),
.B(n_19893),
.C(n_19853),
.Y(n_20008)
);

NAND4xp75_ASAP7_75t_L g20009 ( 
.A(n_19928),
.B(n_3933),
.C(n_3931),
.D(n_3932),
.Y(n_20009)
);

AND2x2_ASAP7_75t_L g20010 ( 
.A(n_19947),
.B(n_3933),
.Y(n_20010)
);

NOR4xp75_ASAP7_75t_SL g20011 ( 
.A(n_19921),
.B(n_3936),
.C(n_3934),
.D(n_3935),
.Y(n_20011)
);

AND2x2_ASAP7_75t_L g20012 ( 
.A(n_19907),
.B(n_3935),
.Y(n_20012)
);

NOR3xp33_ASAP7_75t_L g20013 ( 
.A(n_19910),
.B(n_3936),
.C(n_3937),
.Y(n_20013)
);

NOR2x1_ASAP7_75t_L g20014 ( 
.A(n_19954),
.B(n_3938),
.Y(n_20014)
);

NAND2xp5_ASAP7_75t_L g20015 ( 
.A(n_19960),
.B(n_3939),
.Y(n_20015)
);

XOR2x2_ASAP7_75t_L g20016 ( 
.A(n_19924),
.B(n_3939),
.Y(n_20016)
);

NAND2xp5_ASAP7_75t_L g20017 ( 
.A(n_19931),
.B(n_3940),
.Y(n_20017)
);

NOR2xp33_ASAP7_75t_L g20018 ( 
.A(n_19992),
.B(n_3941),
.Y(n_20018)
);

INVx1_ASAP7_75t_L g20019 ( 
.A(n_19967),
.Y(n_20019)
);

NOR2x1_ASAP7_75t_L g20020 ( 
.A(n_19984),
.B(n_3942),
.Y(n_20020)
);

A2O1A1Ixp33_ASAP7_75t_L g20021 ( 
.A1(n_19987),
.A2(n_3945),
.B(n_3943),
.C(n_3944),
.Y(n_20021)
);

INVx2_ASAP7_75t_L g20022 ( 
.A(n_19972),
.Y(n_20022)
);

INVx2_ASAP7_75t_SL g20023 ( 
.A(n_19978),
.Y(n_20023)
);

NAND3xp33_ASAP7_75t_SL g20024 ( 
.A(n_19918),
.B(n_3943),
.C(n_3944),
.Y(n_20024)
);

NAND3x2_ASAP7_75t_L g20025 ( 
.A(n_19911),
.B(n_19914),
.C(n_19959),
.Y(n_20025)
);

XNOR2xp5_ASAP7_75t_L g20026 ( 
.A(n_19975),
.B(n_3945),
.Y(n_20026)
);

OAI21xp5_ASAP7_75t_L g20027 ( 
.A1(n_19917),
.A2(n_19936),
.B(n_19985),
.Y(n_20027)
);

AND2x4_ASAP7_75t_L g20028 ( 
.A(n_19943),
.B(n_3946),
.Y(n_20028)
);

NAND4xp25_ASAP7_75t_L g20029 ( 
.A(n_19905),
.B(n_19916),
.C(n_19927),
.D(n_19955),
.Y(n_20029)
);

INVx1_ASAP7_75t_L g20030 ( 
.A(n_19919),
.Y(n_20030)
);

NAND3xp33_ASAP7_75t_L g20031 ( 
.A(n_19909),
.B(n_3946),
.C(n_3947),
.Y(n_20031)
);

NAND4xp75_ASAP7_75t_L g20032 ( 
.A(n_19904),
.B(n_3949),
.C(n_3947),
.D(n_3948),
.Y(n_20032)
);

NOR2xp67_ASAP7_75t_L g20033 ( 
.A(n_19957),
.B(n_3948),
.Y(n_20033)
);

A2O1A1Ixp33_ASAP7_75t_L g20034 ( 
.A1(n_19980),
.A2(n_3951),
.B(n_3949),
.C(n_3950),
.Y(n_20034)
);

CKINVDCx16_ASAP7_75t_R g20035 ( 
.A(n_19914),
.Y(n_20035)
);

NAND3xp33_ASAP7_75t_SL g20036 ( 
.A(n_19920),
.B(n_3950),
.C(n_3952),
.Y(n_20036)
);

BUFx2_ASAP7_75t_L g20037 ( 
.A(n_19990),
.Y(n_20037)
);

NAND2xp5_ASAP7_75t_L g20038 ( 
.A(n_19926),
.B(n_19941),
.Y(n_20038)
);

NOR2x1_ASAP7_75t_L g20039 ( 
.A(n_19964),
.B(n_3952),
.Y(n_20039)
);

NOR3xp33_ASAP7_75t_L g20040 ( 
.A(n_19913),
.B(n_3953),
.C(n_3954),
.Y(n_20040)
);

NOR3x2_ASAP7_75t_L g20041 ( 
.A(n_19986),
.B(n_3953),
.C(n_3954),
.Y(n_20041)
);

OAI221xp5_ASAP7_75t_L g20042 ( 
.A1(n_19956),
.A2(n_3957),
.B1(n_3955),
.B2(n_3956),
.C(n_3958),
.Y(n_20042)
);

NOR3x1_ASAP7_75t_L g20043 ( 
.A(n_19953),
.B(n_3955),
.C(n_3956),
.Y(n_20043)
);

AND2x4_ASAP7_75t_L g20044 ( 
.A(n_19911),
.B(n_19974),
.Y(n_20044)
);

AOI221x1_ASAP7_75t_L g20045 ( 
.A1(n_19908),
.A2(n_3960),
.B1(n_3958),
.B2(n_3959),
.C(n_3961),
.Y(n_20045)
);

OAI211xp5_ASAP7_75t_SL g20046 ( 
.A1(n_19946),
.A2(n_3962),
.B(n_3959),
.C(n_3961),
.Y(n_20046)
);

NAND4xp75_ASAP7_75t_L g20047 ( 
.A(n_19989),
.B(n_3964),
.C(n_3962),
.D(n_3963),
.Y(n_20047)
);

OR2x2_ASAP7_75t_L g20048 ( 
.A(n_19932),
.B(n_3964),
.Y(n_20048)
);

OAI22xp5_ASAP7_75t_L g20049 ( 
.A1(n_19961),
.A2(n_3967),
.B1(n_3965),
.B2(n_3966),
.Y(n_20049)
);

INVx1_ASAP7_75t_L g20050 ( 
.A(n_19937),
.Y(n_20050)
);

NOR2x1_ASAP7_75t_L g20051 ( 
.A(n_19993),
.B(n_19938),
.Y(n_20051)
);

NAND3xp33_ASAP7_75t_L g20052 ( 
.A(n_19977),
.B(n_3965),
.C(n_3966),
.Y(n_20052)
);

O2A1O1Ixp33_ASAP7_75t_L g20053 ( 
.A1(n_19935),
.A2(n_3969),
.B(n_3967),
.C(n_3968),
.Y(n_20053)
);

OAI21xp5_ASAP7_75t_L g20054 ( 
.A1(n_19929),
.A2(n_3968),
.B(n_3969),
.Y(n_20054)
);

OAI211xp5_ASAP7_75t_SL g20055 ( 
.A1(n_19973),
.A2(n_3972),
.B(n_3970),
.C(n_3971),
.Y(n_20055)
);

AND2x2_ASAP7_75t_L g20056 ( 
.A(n_19991),
.B(n_3970),
.Y(n_20056)
);

OR2x2_ASAP7_75t_L g20057 ( 
.A(n_19951),
.B(n_3972),
.Y(n_20057)
);

NAND3xp33_ASAP7_75t_L g20058 ( 
.A(n_19933),
.B(n_3973),
.C(n_3974),
.Y(n_20058)
);

INVx1_ASAP7_75t_L g20059 ( 
.A(n_19945),
.Y(n_20059)
);

NAND4xp75_ASAP7_75t_L g20060 ( 
.A(n_19983),
.B(n_3975),
.C(n_3973),
.D(n_3974),
.Y(n_20060)
);

NAND4xp25_ASAP7_75t_L g20061 ( 
.A(n_19976),
.B(n_3977),
.C(n_3975),
.D(n_3976),
.Y(n_20061)
);

NOR2x1_ASAP7_75t_L g20062 ( 
.A(n_19949),
.B(n_3976),
.Y(n_20062)
);

NAND4xp75_ASAP7_75t_L g20063 ( 
.A(n_19970),
.B(n_3979),
.C(n_3977),
.D(n_3978),
.Y(n_20063)
);

AND2x2_ASAP7_75t_L g20064 ( 
.A(n_19966),
.B(n_3978),
.Y(n_20064)
);

OAI221xp5_ASAP7_75t_L g20065 ( 
.A1(n_19988),
.A2(n_3981),
.B1(n_3979),
.B2(n_3980),
.C(n_3982),
.Y(n_20065)
);

NOR2x1_ASAP7_75t_L g20066 ( 
.A(n_19979),
.B(n_3980),
.Y(n_20066)
);

INVx1_ASAP7_75t_L g20067 ( 
.A(n_19965),
.Y(n_20067)
);

INVx2_ASAP7_75t_L g20068 ( 
.A(n_19950),
.Y(n_20068)
);

OR2x2_ASAP7_75t_L g20069 ( 
.A(n_19994),
.B(n_3981),
.Y(n_20069)
);

NAND3xp33_ASAP7_75t_L g20070 ( 
.A(n_19958),
.B(n_3983),
.C(n_3985),
.Y(n_20070)
);

NOR2xp33_ASAP7_75t_L g20071 ( 
.A(n_19939),
.B(n_19923),
.Y(n_20071)
);

AO22x2_ASAP7_75t_L g20072 ( 
.A1(n_19968),
.A2(n_19950),
.B1(n_19952),
.B2(n_19981),
.Y(n_20072)
);

AND2x2_ASAP7_75t_L g20073 ( 
.A(n_19948),
.B(n_3985),
.Y(n_20073)
);

NAND3xp33_ASAP7_75t_L g20074 ( 
.A(n_19971),
.B(n_3986),
.C(n_3987),
.Y(n_20074)
);

AND2x2_ASAP7_75t_L g20075 ( 
.A(n_19982),
.B(n_3986),
.Y(n_20075)
);

INVx1_ASAP7_75t_L g20076 ( 
.A(n_19924),
.Y(n_20076)
);

HB1xp67_ASAP7_75t_L g20077 ( 
.A(n_19925),
.Y(n_20077)
);

OAI21xp5_ASAP7_75t_L g20078 ( 
.A1(n_19944),
.A2(n_3987),
.B(n_3988),
.Y(n_20078)
);

OAI22xp5_ASAP7_75t_L g20079 ( 
.A1(n_19930),
.A2(n_3991),
.B1(n_3989),
.B2(n_3990),
.Y(n_20079)
);

NOR2x1_ASAP7_75t_L g20080 ( 
.A(n_19925),
.B(n_3989),
.Y(n_20080)
);

NOR2x1p5_ASAP7_75t_L g20081 ( 
.A(n_19915),
.B(n_3990),
.Y(n_20081)
);

NAND2xp5_ASAP7_75t_L g20082 ( 
.A(n_19925),
.B(n_3991),
.Y(n_20082)
);

NOR3xp33_ASAP7_75t_L g20083 ( 
.A(n_19906),
.B(n_3992),
.C(n_3993),
.Y(n_20083)
);

INVx1_ASAP7_75t_L g20084 ( 
.A(n_19924),
.Y(n_20084)
);

INVx1_ASAP7_75t_L g20085 ( 
.A(n_19924),
.Y(n_20085)
);

NAND3xp33_ASAP7_75t_SL g20086 ( 
.A(n_19992),
.B(n_3992),
.C(n_3993),
.Y(n_20086)
);

NOR2xp67_ASAP7_75t_L g20087 ( 
.A(n_19919),
.B(n_3994),
.Y(n_20087)
);

OR2x2_ASAP7_75t_L g20088 ( 
.A(n_19930),
.B(n_3994),
.Y(n_20088)
);

OAI22x1_ASAP7_75t_L g20089 ( 
.A1(n_19947),
.A2(n_3997),
.B1(n_3995),
.B2(n_3996),
.Y(n_20089)
);

HB1xp67_ASAP7_75t_L g20090 ( 
.A(n_19925),
.Y(n_20090)
);

AND2x2_ASAP7_75t_L g20091 ( 
.A(n_19934),
.B(n_3995),
.Y(n_20091)
);

NOR3xp33_ASAP7_75t_L g20092 ( 
.A(n_19906),
.B(n_3996),
.C(n_3997),
.Y(n_20092)
);

INVx1_ASAP7_75t_L g20093 ( 
.A(n_19924),
.Y(n_20093)
);

INVx1_ASAP7_75t_SL g20094 ( 
.A(n_20012),
.Y(n_20094)
);

AOI21xp5_ASAP7_75t_L g20095 ( 
.A1(n_20001),
.A2(n_3998),
.B(n_3999),
.Y(n_20095)
);

AOI211xp5_ASAP7_75t_L g20096 ( 
.A1(n_20087),
.A2(n_4000),
.B(n_3998),
.C(n_3999),
.Y(n_20096)
);

OR3x2_ASAP7_75t_L g20097 ( 
.A(n_20029),
.B(n_4000),
.C(n_4001),
.Y(n_20097)
);

AOI22xp5_ASAP7_75t_L g20098 ( 
.A1(n_20005),
.A2(n_4003),
.B1(n_4001),
.B2(n_4002),
.Y(n_20098)
);

OAI211xp5_ASAP7_75t_L g20099 ( 
.A1(n_20025),
.A2(n_4005),
.B(n_4003),
.C(n_4004),
.Y(n_20099)
);

NAND4xp75_ASAP7_75t_L g20100 ( 
.A(n_20004),
.B(n_4006),
.C(n_4004),
.D(n_4005),
.Y(n_20100)
);

AOI21xp33_ASAP7_75t_SL g20101 ( 
.A1(n_20035),
.A2(n_4006),
.B(n_4007),
.Y(n_20101)
);

INVx1_ASAP7_75t_L g20102 ( 
.A(n_20091),
.Y(n_20102)
);

XNOR2xp5_ASAP7_75t_L g20103 ( 
.A(n_20041),
.B(n_4008),
.Y(n_20103)
);

AOI21xp5_ASAP7_75t_L g20104 ( 
.A1(n_20030),
.A2(n_4008),
.B(n_4009),
.Y(n_20104)
);

NOR3xp33_ASAP7_75t_L g20105 ( 
.A(n_20003),
.B(n_4009),
.C(n_4010),
.Y(n_20105)
);

AOI221xp5_ASAP7_75t_L g20106 ( 
.A1(n_20042),
.A2(n_4012),
.B1(n_4010),
.B2(n_4011),
.C(n_4013),
.Y(n_20106)
);

AND2x4_ASAP7_75t_L g20107 ( 
.A(n_20062),
.B(n_4011),
.Y(n_20107)
);

NAND2xp5_ASAP7_75t_L g20108 ( 
.A(n_20033),
.B(n_4012),
.Y(n_20108)
);

NOR3xp33_ASAP7_75t_L g20109 ( 
.A(n_20027),
.B(n_4013),
.C(n_4015),
.Y(n_20109)
);

BUFx2_ASAP7_75t_L g20110 ( 
.A(n_20078),
.Y(n_20110)
);

AND2x4_ASAP7_75t_L g20111 ( 
.A(n_20080),
.B(n_4016),
.Y(n_20111)
);

NAND3xp33_ASAP7_75t_L g20112 ( 
.A(n_19996),
.B(n_4016),
.C(n_4017),
.Y(n_20112)
);

OR2x2_ASAP7_75t_L g20113 ( 
.A(n_20036),
.B(n_4018),
.Y(n_20113)
);

NAND2xp5_ASAP7_75t_L g20114 ( 
.A(n_20010),
.B(n_4018),
.Y(n_20114)
);

AND2x2_ASAP7_75t_L g20115 ( 
.A(n_20073),
.B(n_4019),
.Y(n_20115)
);

NOR3xp33_ASAP7_75t_SL g20116 ( 
.A(n_20008),
.B(n_20084),
.C(n_20076),
.Y(n_20116)
);

NOR2x1_ASAP7_75t_L g20117 ( 
.A(n_20081),
.B(n_20085),
.Y(n_20117)
);

OAI22xp5_ASAP7_75t_L g20118 ( 
.A1(n_20058),
.A2(n_4021),
.B1(n_4019),
.B2(n_4020),
.Y(n_20118)
);

AOI21xp5_ASAP7_75t_L g20119 ( 
.A1(n_20077),
.A2(n_4020),
.B(n_4021),
.Y(n_20119)
);

O2A1O1Ixp33_ASAP7_75t_L g20120 ( 
.A1(n_20090),
.A2(n_4024),
.B(n_4022),
.C(n_4023),
.Y(n_20120)
);

AND2x2_ASAP7_75t_SL g20121 ( 
.A(n_20022),
.B(n_4022),
.Y(n_20121)
);

INVx1_ASAP7_75t_L g20122 ( 
.A(n_20082),
.Y(n_20122)
);

AND2x4_ASAP7_75t_L g20123 ( 
.A(n_20014),
.B(n_4023),
.Y(n_20123)
);

AOI22xp5_ASAP7_75t_L g20124 ( 
.A1(n_20024),
.A2(n_4026),
.B1(n_4024),
.B2(n_4025),
.Y(n_20124)
);

NAND4xp25_ASAP7_75t_L g20125 ( 
.A(n_20017),
.B(n_20071),
.C(n_20054),
.D(n_20000),
.Y(n_20125)
);

NOR3xp33_ASAP7_75t_L g20126 ( 
.A(n_20093),
.B(n_4025),
.C(n_4026),
.Y(n_20126)
);

OR2x2_ASAP7_75t_L g20127 ( 
.A(n_20086),
.B(n_4027),
.Y(n_20127)
);

OAI21xp33_ASAP7_75t_SL g20128 ( 
.A1(n_20061),
.A2(n_4028),
.B(n_4029),
.Y(n_20128)
);

NOR3xp33_ASAP7_75t_SL g20129 ( 
.A(n_20019),
.B(n_20059),
.C(n_20050),
.Y(n_20129)
);

NAND3xp33_ASAP7_75t_L g20130 ( 
.A(n_19999),
.B(n_4028),
.C(n_4029),
.Y(n_20130)
);

AOI221xp5_ASAP7_75t_L g20131 ( 
.A1(n_20074),
.A2(n_4032),
.B1(n_4030),
.B2(n_4031),
.C(n_4033),
.Y(n_20131)
);

AND2x2_ASAP7_75t_L g20132 ( 
.A(n_20075),
.B(n_4030),
.Y(n_20132)
);

NOR2xp33_ASAP7_75t_L g20133 ( 
.A(n_20069),
.B(n_20048),
.Y(n_20133)
);

NOR2x1p5_ASAP7_75t_L g20134 ( 
.A(n_20015),
.B(n_4032),
.Y(n_20134)
);

NAND4xp25_ASAP7_75t_L g20135 ( 
.A(n_20043),
.B(n_20070),
.C(n_20038),
.D(n_20007),
.Y(n_20135)
);

OAI322xp33_ASAP7_75t_L g20136 ( 
.A1(n_20057),
.A2(n_4038),
.A3(n_4037),
.B1(n_4035),
.B2(n_4033),
.C1(n_4034),
.C2(n_4036),
.Y(n_20136)
);

XNOR2x1_ASAP7_75t_L g20137 ( 
.A(n_20016),
.B(n_4034),
.Y(n_20137)
);

NAND2xp5_ASAP7_75t_L g20138 ( 
.A(n_20083),
.B(n_4036),
.Y(n_20138)
);

NAND4xp75_ASAP7_75t_L g20139 ( 
.A(n_19999),
.B(n_4039),
.C(n_4037),
.D(n_4038),
.Y(n_20139)
);

NOR2x1_ASAP7_75t_L g20140 ( 
.A(n_20060),
.B(n_4039),
.Y(n_20140)
);

AOI222xp33_ASAP7_75t_L g20141 ( 
.A1(n_20056),
.A2(n_4042),
.B1(n_4044),
.B2(n_4040),
.C1(n_4041),
.C2(n_4043),
.Y(n_20141)
);

NOR2x1_ASAP7_75t_L g20142 ( 
.A(n_20068),
.B(n_4040),
.Y(n_20142)
);

NOR2x1_ASAP7_75t_L g20143 ( 
.A(n_20039),
.B(n_4041),
.Y(n_20143)
);

XNOR2x1_ASAP7_75t_L g20144 ( 
.A(n_20020),
.B(n_4042),
.Y(n_20144)
);

NOR2x1_ASAP7_75t_L g20145 ( 
.A(n_19998),
.B(n_4043),
.Y(n_20145)
);

AOI21xp5_ASAP7_75t_L g20146 ( 
.A1(n_20002),
.A2(n_4044),
.B(n_4045),
.Y(n_20146)
);

INVx1_ASAP7_75t_L g20147 ( 
.A(n_20064),
.Y(n_20147)
);

AOI22xp5_ASAP7_75t_L g20148 ( 
.A1(n_20092),
.A2(n_4047),
.B1(n_4045),
.B2(n_4046),
.Y(n_20148)
);

AOI32xp33_ASAP7_75t_L g20149 ( 
.A1(n_20066),
.A2(n_4048),
.A3(n_4046),
.B1(n_4047),
.B2(n_4049),
.Y(n_20149)
);

NAND3xp33_ASAP7_75t_SL g20150 ( 
.A(n_20037),
.B(n_4048),
.C(n_4049),
.Y(n_20150)
);

INVxp67_ASAP7_75t_L g20151 ( 
.A(n_20018),
.Y(n_20151)
);

O2A1O1Ixp33_ASAP7_75t_L g20152 ( 
.A1(n_20023),
.A2(n_4052),
.B(n_4050),
.C(n_4051),
.Y(n_20152)
);

NAND3xp33_ASAP7_75t_L g20153 ( 
.A(n_20067),
.B(n_4050),
.C(n_4051),
.Y(n_20153)
);

AND2x4_ASAP7_75t_L g20154 ( 
.A(n_20051),
.B(n_4052),
.Y(n_20154)
);

AOI21xp33_ASAP7_75t_SL g20155 ( 
.A1(n_20089),
.A2(n_4053),
.B(n_4054),
.Y(n_20155)
);

NOR3xp33_ASAP7_75t_L g20156 ( 
.A(n_20044),
.B(n_4053),
.C(n_4054),
.Y(n_20156)
);

NAND2xp5_ASAP7_75t_L g20157 ( 
.A(n_20021),
.B(n_4055),
.Y(n_20157)
);

AOI22xp5_ASAP7_75t_L g20158 ( 
.A1(n_20055),
.A2(n_4058),
.B1(n_4055),
.B2(n_4056),
.Y(n_20158)
);

AOI22xp33_ASAP7_75t_SL g20159 ( 
.A1(n_20065),
.A2(n_4059),
.B1(n_4056),
.B2(n_4058),
.Y(n_20159)
);

OR3x1_ASAP7_75t_L g20160 ( 
.A(n_20046),
.B(n_4062),
.C(n_4061),
.Y(n_20160)
);

OAI221xp5_ASAP7_75t_SL g20161 ( 
.A1(n_20034),
.A2(n_4062),
.B1(n_4060),
.B2(n_4061),
.C(n_4063),
.Y(n_20161)
);

AND2x4_ASAP7_75t_L g20162 ( 
.A(n_19998),
.B(n_4060),
.Y(n_20162)
);

OAI21xp5_ASAP7_75t_SL g20163 ( 
.A1(n_20006),
.A2(n_4064),
.B(n_4065),
.Y(n_20163)
);

NOR2x1p5_ASAP7_75t_L g20164 ( 
.A(n_20063),
.B(n_19997),
.Y(n_20164)
);

NAND2xp5_ASAP7_75t_SL g20165 ( 
.A(n_20011),
.B(n_4064),
.Y(n_20165)
);

INVx1_ASAP7_75t_L g20166 ( 
.A(n_20026),
.Y(n_20166)
);

OR2x2_ASAP7_75t_L g20167 ( 
.A(n_20049),
.B(n_4065),
.Y(n_20167)
);

AND2x4_ASAP7_75t_L g20168 ( 
.A(n_20044),
.B(n_4066),
.Y(n_20168)
);

OAI21xp5_ASAP7_75t_L g20169 ( 
.A1(n_20053),
.A2(n_4066),
.B(n_4067),
.Y(n_20169)
);

AOI21xp33_ASAP7_75t_L g20170 ( 
.A1(n_20072),
.A2(n_4067),
.B(n_4068),
.Y(n_20170)
);

AND4x1_ASAP7_75t_L g20171 ( 
.A(n_20040),
.B(n_4070),
.C(n_4071),
.D(n_4069),
.Y(n_20171)
);

NAND4xp75_ASAP7_75t_L g20172 ( 
.A(n_20045),
.B(n_4070),
.C(n_4068),
.D(n_4069),
.Y(n_20172)
);

AOI22xp5_ASAP7_75t_L g20173 ( 
.A1(n_20013),
.A2(n_4073),
.B1(n_4071),
.B2(n_4072),
.Y(n_20173)
);

INVx1_ASAP7_75t_L g20174 ( 
.A(n_20088),
.Y(n_20174)
);

AND2x4_ASAP7_75t_L g20175 ( 
.A(n_20031),
.B(n_4072),
.Y(n_20175)
);

OR2x2_ASAP7_75t_L g20176 ( 
.A(n_20052),
.B(n_4073),
.Y(n_20176)
);

NOR2xp33_ASAP7_75t_L g20177 ( 
.A(n_20079),
.B(n_4074),
.Y(n_20177)
);

OR2x2_ASAP7_75t_L g20178 ( 
.A(n_20032),
.B(n_4074),
.Y(n_20178)
);

AOI21xp5_ASAP7_75t_L g20179 ( 
.A1(n_20072),
.A2(n_4075),
.B(n_4076),
.Y(n_20179)
);

NOR3xp33_ASAP7_75t_L g20180 ( 
.A(n_19995),
.B(n_20009),
.C(n_20047),
.Y(n_20180)
);

OAI221xp5_ASAP7_75t_L g20181 ( 
.A1(n_20028),
.A2(n_4077),
.B1(n_4075),
.B2(n_4076),
.C(n_4078),
.Y(n_20181)
);

AND3x4_ASAP7_75t_L g20182 ( 
.A(n_20028),
.B(n_4078),
.C(n_4079),
.Y(n_20182)
);

NAND4xp25_ASAP7_75t_L g20183 ( 
.A(n_20087),
.B(n_4081),
.C(n_4079),
.D(n_4080),
.Y(n_20183)
);

NOR3x1_ASAP7_75t_L g20184 ( 
.A(n_20008),
.B(n_4080),
.C(n_4081),
.Y(n_20184)
);

INVx1_ASAP7_75t_L g20185 ( 
.A(n_20091),
.Y(n_20185)
);

AND2x4_ASAP7_75t_L g20186 ( 
.A(n_20087),
.B(n_4082),
.Y(n_20186)
);

OAI321xp33_ASAP7_75t_L g20187 ( 
.A1(n_20012),
.A2(n_4084),
.A3(n_4086),
.B1(n_4082),
.B2(n_4083),
.C(n_4085),
.Y(n_20187)
);

NAND4xp75_ASAP7_75t_L g20188 ( 
.A(n_20004),
.B(n_4086),
.C(n_4083),
.D(n_4084),
.Y(n_20188)
);

NAND3xp33_ASAP7_75t_SL g20189 ( 
.A(n_20005),
.B(n_4087),
.C(n_4088),
.Y(n_20189)
);

AND2x2_ASAP7_75t_L g20190 ( 
.A(n_20012),
.B(n_4087),
.Y(n_20190)
);

NAND3xp33_ASAP7_75t_SL g20191 ( 
.A(n_20005),
.B(n_4089),
.C(n_4090),
.Y(n_20191)
);

OR2x2_ASAP7_75t_L g20192 ( 
.A(n_20036),
.B(n_4089),
.Y(n_20192)
);

NAND4xp75_ASAP7_75t_L g20193 ( 
.A(n_20004),
.B(n_4092),
.C(n_4090),
.D(n_4091),
.Y(n_20193)
);

NAND3xp33_ASAP7_75t_SL g20194 ( 
.A(n_20005),
.B(n_4091),
.C(n_4093),
.Y(n_20194)
);

AOI221xp5_ASAP7_75t_L g20195 ( 
.A1(n_20042),
.A2(n_4095),
.B1(n_4093),
.B2(n_4094),
.C(n_4096),
.Y(n_20195)
);

INVx1_ASAP7_75t_L g20196 ( 
.A(n_20091),
.Y(n_20196)
);

XNOR2x1_ASAP7_75t_L g20197 ( 
.A(n_20005),
.B(n_4096),
.Y(n_20197)
);

OAI211xp5_ASAP7_75t_SL g20198 ( 
.A1(n_20030),
.A2(n_4099),
.B(n_4097),
.C(n_4098),
.Y(n_20198)
);

NAND4xp75_ASAP7_75t_L g20199 ( 
.A(n_20004),
.B(n_4099),
.C(n_4097),
.D(n_4098),
.Y(n_20199)
);

AND2x2_ASAP7_75t_L g20200 ( 
.A(n_20012),
.B(n_4100),
.Y(n_20200)
);

AND2x2_ASAP7_75t_L g20201 ( 
.A(n_20012),
.B(n_4100),
.Y(n_20201)
);

NOR2x1p5_ASAP7_75t_L g20202 ( 
.A(n_20015),
.B(n_4101),
.Y(n_20202)
);

INVxp67_ASAP7_75t_L g20203 ( 
.A(n_20091),
.Y(n_20203)
);

NAND3xp33_ASAP7_75t_L g20204 ( 
.A(n_19996),
.B(n_4101),
.C(n_4102),
.Y(n_20204)
);

NAND2xp5_ASAP7_75t_L g20205 ( 
.A(n_20091),
.B(n_4102),
.Y(n_20205)
);

AND2x2_ASAP7_75t_L g20206 ( 
.A(n_20012),
.B(n_4103),
.Y(n_20206)
);

INVx1_ASAP7_75t_L g20207 ( 
.A(n_20091),
.Y(n_20207)
);

NAND4xp75_ASAP7_75t_L g20208 ( 
.A(n_20004),
.B(n_4105),
.C(n_4103),
.D(n_4104),
.Y(n_20208)
);

NOR2x1p5_ASAP7_75t_L g20209 ( 
.A(n_20015),
.B(n_4104),
.Y(n_20209)
);

XOR2x1_ASAP7_75t_L g20210 ( 
.A(n_20081),
.B(n_4105),
.Y(n_20210)
);

INVx1_ASAP7_75t_L g20211 ( 
.A(n_20091),
.Y(n_20211)
);

OAI221xp5_ASAP7_75t_L g20212 ( 
.A1(n_20034),
.A2(n_4108),
.B1(n_4106),
.B2(n_4107),
.C(n_4109),
.Y(n_20212)
);

INVxp67_ASAP7_75t_L g20213 ( 
.A(n_20091),
.Y(n_20213)
);

NAND2xp5_ASAP7_75t_SL g20214 ( 
.A(n_20011),
.B(n_4106),
.Y(n_20214)
);

NAND2xp5_ASAP7_75t_L g20215 ( 
.A(n_20091),
.B(n_4107),
.Y(n_20215)
);

INVx1_ASAP7_75t_SL g20216 ( 
.A(n_20137),
.Y(n_20216)
);

HB1xp67_ASAP7_75t_L g20217 ( 
.A(n_20123),
.Y(n_20217)
);

CKINVDCx5p33_ASAP7_75t_R g20218 ( 
.A(n_20116),
.Y(n_20218)
);

AND2x4_ASAP7_75t_SL g20219 ( 
.A(n_20107),
.B(n_4108),
.Y(n_20219)
);

BUFx6f_ASAP7_75t_L g20220 ( 
.A(n_20102),
.Y(n_20220)
);

INVx1_ASAP7_75t_L g20221 ( 
.A(n_20165),
.Y(n_20221)
);

INVx1_ASAP7_75t_L g20222 ( 
.A(n_20214),
.Y(n_20222)
);

CKINVDCx5p33_ASAP7_75t_R g20223 ( 
.A(n_20129),
.Y(n_20223)
);

BUFx6f_ASAP7_75t_L g20224 ( 
.A(n_20185),
.Y(n_20224)
);

BUFx2_ASAP7_75t_L g20225 ( 
.A(n_20123),
.Y(n_20225)
);

CKINVDCx5p33_ASAP7_75t_R g20226 ( 
.A(n_20094),
.Y(n_20226)
);

BUFx2_ASAP7_75t_L g20227 ( 
.A(n_20111),
.Y(n_20227)
);

INVx1_ASAP7_75t_L g20228 ( 
.A(n_20186),
.Y(n_20228)
);

INVx2_ASAP7_75t_L g20229 ( 
.A(n_20197),
.Y(n_20229)
);

NOR3xp33_ASAP7_75t_L g20230 ( 
.A(n_20135),
.B(n_4109),
.C(n_4110),
.Y(n_20230)
);

INVx3_ASAP7_75t_SL g20231 ( 
.A(n_20144),
.Y(n_20231)
);

INVx1_ASAP7_75t_L g20232 ( 
.A(n_20186),
.Y(n_20232)
);

CKINVDCx5p33_ASAP7_75t_R g20233 ( 
.A(n_20196),
.Y(n_20233)
);

CKINVDCx5p33_ASAP7_75t_R g20234 ( 
.A(n_20207),
.Y(n_20234)
);

CKINVDCx5p33_ASAP7_75t_R g20235 ( 
.A(n_20211),
.Y(n_20235)
);

BUFx6f_ASAP7_75t_L g20236 ( 
.A(n_20122),
.Y(n_20236)
);

INVx1_ASAP7_75t_SL g20237 ( 
.A(n_20210),
.Y(n_20237)
);

HB1xp67_ASAP7_75t_L g20238 ( 
.A(n_20142),
.Y(n_20238)
);

OAI22xp5_ASAP7_75t_L g20239 ( 
.A1(n_20097),
.A2(n_4112),
.B1(n_4113),
.B2(n_4111),
.Y(n_20239)
);

OAI22xp33_ASAP7_75t_L g20240 ( 
.A1(n_20124),
.A2(n_4118),
.B1(n_4126),
.B2(n_4110),
.Y(n_20240)
);

AND2x2_ASAP7_75t_L g20241 ( 
.A(n_20134),
.B(n_20202),
.Y(n_20241)
);

INVx1_ASAP7_75t_SL g20242 ( 
.A(n_20114),
.Y(n_20242)
);

HB1xp67_ASAP7_75t_L g20243 ( 
.A(n_20145),
.Y(n_20243)
);

INVx2_ASAP7_75t_L g20244 ( 
.A(n_20139),
.Y(n_20244)
);

CKINVDCx5p33_ASAP7_75t_R g20245 ( 
.A(n_20203),
.Y(n_20245)
);

BUFx2_ASAP7_75t_L g20246 ( 
.A(n_20111),
.Y(n_20246)
);

CKINVDCx6p67_ASAP7_75t_R g20247 ( 
.A(n_20110),
.Y(n_20247)
);

AOI32xp33_ASAP7_75t_L g20248 ( 
.A1(n_20140),
.A2(n_4113),
.A3(n_4111),
.B1(n_4112),
.B2(n_4114),
.Y(n_20248)
);

AND2x4_ASAP7_75t_L g20249 ( 
.A(n_20143),
.B(n_4114),
.Y(n_20249)
);

NOR2xp33_ASAP7_75t_R g20250 ( 
.A(n_20103),
.B(n_4115),
.Y(n_20250)
);

NOR3xp33_ASAP7_75t_L g20251 ( 
.A(n_20125),
.B(n_4116),
.C(n_4117),
.Y(n_20251)
);

BUFx2_ASAP7_75t_L g20252 ( 
.A(n_20107),
.Y(n_20252)
);

OAI22xp5_ASAP7_75t_L g20253 ( 
.A1(n_20112),
.A2(n_4119),
.B1(n_4120),
.B2(n_4117),
.Y(n_20253)
);

NOR2xp33_ASAP7_75t_L g20254 ( 
.A(n_20128),
.B(n_4116),
.Y(n_20254)
);

BUFx2_ASAP7_75t_L g20255 ( 
.A(n_20115),
.Y(n_20255)
);

BUFx2_ASAP7_75t_L g20256 ( 
.A(n_20132),
.Y(n_20256)
);

CKINVDCx5p33_ASAP7_75t_R g20257 ( 
.A(n_20213),
.Y(n_20257)
);

INVx1_ASAP7_75t_L g20258 ( 
.A(n_20108),
.Y(n_20258)
);

CKINVDCx16_ASAP7_75t_R g20259 ( 
.A(n_20117),
.Y(n_20259)
);

BUFx4f_ASAP7_75t_SL g20260 ( 
.A(n_20166),
.Y(n_20260)
);

INVx1_ASAP7_75t_L g20261 ( 
.A(n_20178),
.Y(n_20261)
);

BUFx12f_ASAP7_75t_L g20262 ( 
.A(n_20164),
.Y(n_20262)
);

HB1xp67_ASAP7_75t_L g20263 ( 
.A(n_20130),
.Y(n_20263)
);

INVx1_ASAP7_75t_SL g20264 ( 
.A(n_20113),
.Y(n_20264)
);

INVx1_ASAP7_75t_L g20265 ( 
.A(n_20138),
.Y(n_20265)
);

OAI21xp33_ASAP7_75t_SL g20266 ( 
.A1(n_20172),
.A2(n_4119),
.B(n_4120),
.Y(n_20266)
);

NAND2xp5_ASAP7_75t_SL g20267 ( 
.A(n_20204),
.B(n_4121),
.Y(n_20267)
);

BUFx2_ASAP7_75t_L g20268 ( 
.A(n_20169),
.Y(n_20268)
);

CKINVDCx5p33_ASAP7_75t_R g20269 ( 
.A(n_20133),
.Y(n_20269)
);

INVx2_ASAP7_75t_L g20270 ( 
.A(n_20121),
.Y(n_20270)
);

BUFx10_ASAP7_75t_L g20271 ( 
.A(n_20147),
.Y(n_20271)
);

BUFx12f_ASAP7_75t_L g20272 ( 
.A(n_20209),
.Y(n_20272)
);

INVxp67_ASAP7_75t_L g20273 ( 
.A(n_20192),
.Y(n_20273)
);

INVx1_ASAP7_75t_SL g20274 ( 
.A(n_20205),
.Y(n_20274)
);

CKINVDCx5p33_ASAP7_75t_R g20275 ( 
.A(n_20151),
.Y(n_20275)
);

HB1xp67_ASAP7_75t_L g20276 ( 
.A(n_20182),
.Y(n_20276)
);

CKINVDCx5p33_ASAP7_75t_R g20277 ( 
.A(n_20174),
.Y(n_20277)
);

XNOR2xp5_ASAP7_75t_L g20278 ( 
.A(n_20160),
.B(n_4121),
.Y(n_20278)
);

AO22x2_ASAP7_75t_L g20279 ( 
.A1(n_20180),
.A2(n_4130),
.B1(n_4138),
.B2(n_4122),
.Y(n_20279)
);

OA21x2_ASAP7_75t_L g20280 ( 
.A1(n_20157),
.A2(n_4123),
.B(n_4124),
.Y(n_20280)
);

BUFx2_ASAP7_75t_L g20281 ( 
.A(n_20175),
.Y(n_20281)
);

AOI22xp33_ASAP7_75t_L g20282 ( 
.A1(n_20175),
.A2(n_4125),
.B1(n_4123),
.B2(n_4124),
.Y(n_20282)
);

AOI21xp5_ASAP7_75t_L g20283 ( 
.A1(n_20177),
.A2(n_4125),
.B(n_4126),
.Y(n_20283)
);

CKINVDCx5p33_ASAP7_75t_R g20284 ( 
.A(n_20118),
.Y(n_20284)
);

CKINVDCx5p33_ASAP7_75t_R g20285 ( 
.A(n_20127),
.Y(n_20285)
);

INVx1_ASAP7_75t_L g20286 ( 
.A(n_20176),
.Y(n_20286)
);

INVx1_ASAP7_75t_L g20287 ( 
.A(n_20184),
.Y(n_20287)
);

INVx1_ASAP7_75t_SL g20288 ( 
.A(n_20215),
.Y(n_20288)
);

AOI221xp5_ASAP7_75t_SL g20289 ( 
.A1(n_20155),
.A2(n_20195),
.B1(n_20106),
.B2(n_20167),
.C(n_20212),
.Y(n_20289)
);

INVx1_ASAP7_75t_L g20290 ( 
.A(n_20105),
.Y(n_20290)
);

INVx1_ASAP7_75t_L g20291 ( 
.A(n_20171),
.Y(n_20291)
);

INVx2_ASAP7_75t_SL g20292 ( 
.A(n_20154),
.Y(n_20292)
);

CKINVDCx5p33_ASAP7_75t_R g20293 ( 
.A(n_20159),
.Y(n_20293)
);

AOI221xp5_ASAP7_75t_L g20294 ( 
.A1(n_20161),
.A2(n_4129),
.B1(n_4127),
.B2(n_4128),
.C(n_4130),
.Y(n_20294)
);

BUFx4f_ASAP7_75t_SL g20295 ( 
.A(n_20154),
.Y(n_20295)
);

NOR2xp67_ASAP7_75t_L g20296 ( 
.A(n_20183),
.B(n_4127),
.Y(n_20296)
);

CKINVDCx5p33_ASAP7_75t_R g20297 ( 
.A(n_20158),
.Y(n_20297)
);

HB1xp67_ASAP7_75t_L g20298 ( 
.A(n_20096),
.Y(n_20298)
);

CKINVDCx5p33_ASAP7_75t_R g20299 ( 
.A(n_20173),
.Y(n_20299)
);

CKINVDCx20_ASAP7_75t_R g20300 ( 
.A(n_20148),
.Y(n_20300)
);

INVx1_ASAP7_75t_L g20301 ( 
.A(n_20099),
.Y(n_20301)
);

OAI221xp5_ASAP7_75t_L g20302 ( 
.A1(n_20149),
.A2(n_4131),
.B1(n_4128),
.B2(n_4129),
.C(n_4132),
.Y(n_20302)
);

HB1xp67_ASAP7_75t_L g20303 ( 
.A(n_20179),
.Y(n_20303)
);

O2A1O1Ixp33_ASAP7_75t_SL g20304 ( 
.A1(n_20131),
.A2(n_4134),
.B(n_4135),
.C(n_4133),
.Y(n_20304)
);

CKINVDCx5p33_ASAP7_75t_R g20305 ( 
.A(n_20189),
.Y(n_20305)
);

CKINVDCx16_ASAP7_75t_R g20306 ( 
.A(n_20191),
.Y(n_20306)
);

HB1xp67_ASAP7_75t_L g20307 ( 
.A(n_20100),
.Y(n_20307)
);

AND2x2_ASAP7_75t_L g20308 ( 
.A(n_20109),
.B(n_4132),
.Y(n_20308)
);

INVx1_ASAP7_75t_L g20309 ( 
.A(n_20194),
.Y(n_20309)
);

XOR2xp5_ASAP7_75t_L g20310 ( 
.A(n_20150),
.B(n_4134),
.Y(n_20310)
);

HB1xp67_ASAP7_75t_L g20311 ( 
.A(n_20188),
.Y(n_20311)
);

NOR2xp67_ASAP7_75t_L g20312 ( 
.A(n_20104),
.B(n_4133),
.Y(n_20312)
);

NOR2xp33_ASAP7_75t_L g20313 ( 
.A(n_20198),
.B(n_4135),
.Y(n_20313)
);

INVx2_ASAP7_75t_L g20314 ( 
.A(n_20193),
.Y(n_20314)
);

INVx2_ASAP7_75t_L g20315 ( 
.A(n_20199),
.Y(n_20315)
);

INVx1_ASAP7_75t_SL g20316 ( 
.A(n_20190),
.Y(n_20316)
);

O2A1O1Ixp33_ASAP7_75t_L g20317 ( 
.A1(n_20152),
.A2(n_4139),
.B(n_4140),
.C(n_4137),
.Y(n_20317)
);

CKINVDCx5p33_ASAP7_75t_R g20318 ( 
.A(n_20146),
.Y(n_20318)
);

CKINVDCx5p33_ASAP7_75t_R g20319 ( 
.A(n_20095),
.Y(n_20319)
);

BUFx2_ASAP7_75t_L g20320 ( 
.A(n_20153),
.Y(n_20320)
);

CKINVDCx16_ASAP7_75t_R g20321 ( 
.A(n_20098),
.Y(n_20321)
);

INVx1_ASAP7_75t_SL g20322 ( 
.A(n_20200),
.Y(n_20322)
);

CKINVDCx5p33_ASAP7_75t_R g20323 ( 
.A(n_20119),
.Y(n_20323)
);

HB1xp67_ASAP7_75t_L g20324 ( 
.A(n_20208),
.Y(n_20324)
);

CKINVDCx20_ASAP7_75t_R g20325 ( 
.A(n_20170),
.Y(n_20325)
);

NOR2xp67_ASAP7_75t_L g20326 ( 
.A(n_20101),
.B(n_4136),
.Y(n_20326)
);

NOR2x1_ASAP7_75t_L g20327 ( 
.A(n_20163),
.B(n_4137),
.Y(n_20327)
);

HB1xp67_ASAP7_75t_L g20328 ( 
.A(n_20126),
.Y(n_20328)
);

INVx1_ASAP7_75t_L g20329 ( 
.A(n_20136),
.Y(n_20329)
);

HB1xp67_ASAP7_75t_L g20330 ( 
.A(n_20156),
.Y(n_20330)
);

AOI22xp5_ASAP7_75t_L g20331 ( 
.A1(n_20141),
.A2(n_4141),
.B1(n_4136),
.B2(n_4139),
.Y(n_20331)
);

INVx1_ASAP7_75t_L g20332 ( 
.A(n_20120),
.Y(n_20332)
);

CKINVDCx5p33_ASAP7_75t_R g20333 ( 
.A(n_20162),
.Y(n_20333)
);

CKINVDCx5p33_ASAP7_75t_R g20334 ( 
.A(n_20162),
.Y(n_20334)
);

CKINVDCx20_ASAP7_75t_R g20335 ( 
.A(n_20201),
.Y(n_20335)
);

BUFx2_ASAP7_75t_L g20336 ( 
.A(n_20206),
.Y(n_20336)
);

HB1xp67_ASAP7_75t_L g20337 ( 
.A(n_20181),
.Y(n_20337)
);

CKINVDCx5p33_ASAP7_75t_R g20338 ( 
.A(n_20168),
.Y(n_20338)
);

BUFx2_ASAP7_75t_L g20339 ( 
.A(n_20168),
.Y(n_20339)
);

XNOR2xp5_ASAP7_75t_L g20340 ( 
.A(n_20187),
.B(n_4142),
.Y(n_20340)
);

CKINVDCx20_ASAP7_75t_R g20341 ( 
.A(n_20116),
.Y(n_20341)
);

INVx1_ASAP7_75t_L g20342 ( 
.A(n_20165),
.Y(n_20342)
);

NAND2xp33_ASAP7_75t_R g20343 ( 
.A(n_20116),
.B(n_4144),
.Y(n_20343)
);

HB1xp67_ASAP7_75t_L g20344 ( 
.A(n_20123),
.Y(n_20344)
);

HB1xp67_ASAP7_75t_L g20345 ( 
.A(n_20123),
.Y(n_20345)
);

NAND2xp5_ASAP7_75t_L g20346 ( 
.A(n_20123),
.B(n_4143),
.Y(n_20346)
);

OR2x6_ASAP7_75t_L g20347 ( 
.A(n_20117),
.B(n_4144),
.Y(n_20347)
);

CKINVDCx5p33_ASAP7_75t_R g20348 ( 
.A(n_20116),
.Y(n_20348)
);

NOR2xp33_ASAP7_75t_L g20349 ( 
.A(n_20128),
.B(n_4145),
.Y(n_20349)
);

INVx3_ASAP7_75t_SL g20350 ( 
.A(n_20094),
.Y(n_20350)
);

OR2x2_ASAP7_75t_L g20351 ( 
.A(n_20183),
.B(n_4145),
.Y(n_20351)
);

CKINVDCx5p33_ASAP7_75t_R g20352 ( 
.A(n_20116),
.Y(n_20352)
);

NAND2xp33_ASAP7_75t_R g20353 ( 
.A(n_20116),
.B(n_4147),
.Y(n_20353)
);

BUFx12f_ASAP7_75t_L g20354 ( 
.A(n_20164),
.Y(n_20354)
);

AOI31xp33_ASAP7_75t_L g20355 ( 
.A1(n_20221),
.A2(n_4150),
.A3(n_4151),
.B(n_4148),
.Y(n_20355)
);

INVx1_ASAP7_75t_L g20356 ( 
.A(n_20219),
.Y(n_20356)
);

NAND4xp25_ASAP7_75t_L g20357 ( 
.A(n_20343),
.B(n_4151),
.C(n_4146),
.D(n_4150),
.Y(n_20357)
);

AO22x2_ASAP7_75t_L g20358 ( 
.A1(n_20292),
.A2(n_4154),
.B1(n_4152),
.B2(n_4153),
.Y(n_20358)
);

INVx3_ASAP7_75t_SL g20359 ( 
.A(n_20338),
.Y(n_20359)
);

INVx1_ASAP7_75t_L g20360 ( 
.A(n_20249),
.Y(n_20360)
);

NOR2x1_ASAP7_75t_L g20361 ( 
.A(n_20339),
.B(n_4152),
.Y(n_20361)
);

OA22x2_ASAP7_75t_L g20362 ( 
.A1(n_20331),
.A2(n_4156),
.B1(n_4154),
.B2(n_4155),
.Y(n_20362)
);

NAND5xp2_ASAP7_75t_L g20363 ( 
.A(n_20289),
.B(n_4157),
.C(n_4155),
.D(n_4156),
.E(n_4158),
.Y(n_20363)
);

AOI221xp5_ASAP7_75t_L g20364 ( 
.A1(n_20304),
.A2(n_4160),
.B1(n_4157),
.B2(n_4159),
.C(n_4161),
.Y(n_20364)
);

INVx1_ASAP7_75t_L g20365 ( 
.A(n_20249),
.Y(n_20365)
);

AOI22xp5_ASAP7_75t_L g20366 ( 
.A1(n_20341),
.A2(n_4161),
.B1(n_4159),
.B2(n_4160),
.Y(n_20366)
);

AO22x2_ASAP7_75t_L g20367 ( 
.A1(n_20222),
.A2(n_4164),
.B1(n_4162),
.B2(n_4163),
.Y(n_20367)
);

OAI21xp5_ASAP7_75t_L g20368 ( 
.A1(n_20278),
.A2(n_20349),
.B(n_20254),
.Y(n_20368)
);

INVx1_ASAP7_75t_L g20369 ( 
.A(n_20346),
.Y(n_20369)
);

A2O1A1Ixp33_ASAP7_75t_SL g20370 ( 
.A1(n_20342),
.A2(n_4164),
.B(n_4162),
.C(n_4163),
.Y(n_20370)
);

NAND2xp5_ASAP7_75t_L g20371 ( 
.A(n_20326),
.B(n_4165),
.Y(n_20371)
);

OAI22xp5_ASAP7_75t_L g20372 ( 
.A1(n_20302),
.A2(n_4167),
.B1(n_4165),
.B2(n_4166),
.Y(n_20372)
);

INVx2_ASAP7_75t_L g20373 ( 
.A(n_20347),
.Y(n_20373)
);

INVx4_ASAP7_75t_L g20374 ( 
.A(n_20295),
.Y(n_20374)
);

AOI22xp5_ASAP7_75t_L g20375 ( 
.A1(n_20353),
.A2(n_4169),
.B1(n_4167),
.B2(n_4168),
.Y(n_20375)
);

NAND2xp5_ASAP7_75t_L g20376 ( 
.A(n_20296),
.B(n_20312),
.Y(n_20376)
);

CKINVDCx5p33_ASAP7_75t_R g20377 ( 
.A(n_20218),
.Y(n_20377)
);

OAI22xp5_ASAP7_75t_L g20378 ( 
.A1(n_20348),
.A2(n_4170),
.B1(n_4168),
.B2(n_4169),
.Y(n_20378)
);

NAND5xp2_ASAP7_75t_L g20379 ( 
.A(n_20291),
.B(n_4172),
.C(n_4170),
.D(n_4171),
.E(n_4173),
.Y(n_20379)
);

NOR3xp33_ASAP7_75t_L g20380 ( 
.A(n_20259),
.B(n_4171),
.C(n_4173),
.Y(n_20380)
);

INVx1_ASAP7_75t_L g20381 ( 
.A(n_20351),
.Y(n_20381)
);

INVx1_ASAP7_75t_SL g20382 ( 
.A(n_20250),
.Y(n_20382)
);

AND3x1_ASAP7_75t_L g20383 ( 
.A(n_20244),
.B(n_4183),
.C(n_4174),
.Y(n_20383)
);

INVx2_ASAP7_75t_SL g20384 ( 
.A(n_20327),
.Y(n_20384)
);

AOI22xp5_ASAP7_75t_L g20385 ( 
.A1(n_20352),
.A2(n_20239),
.B1(n_20247),
.B2(n_20223),
.Y(n_20385)
);

INVx1_ASAP7_75t_L g20386 ( 
.A(n_20310),
.Y(n_20386)
);

OR2x2_ASAP7_75t_L g20387 ( 
.A(n_20253),
.B(n_4174),
.Y(n_20387)
);

INVx1_ASAP7_75t_L g20388 ( 
.A(n_20340),
.Y(n_20388)
);

AOI211xp5_ASAP7_75t_L g20389 ( 
.A1(n_20350),
.A2(n_4178),
.B(n_4175),
.C(n_4176),
.Y(n_20389)
);

INVx1_ASAP7_75t_L g20390 ( 
.A(n_20280),
.Y(n_20390)
);

NAND4xp75_ASAP7_75t_L g20391 ( 
.A(n_20228),
.B(n_4179),
.C(n_4175),
.D(n_4178),
.Y(n_20391)
);

OA21x2_ASAP7_75t_L g20392 ( 
.A1(n_20232),
.A2(n_4179),
.B(n_4180),
.Y(n_20392)
);

AOI22xp5_ASAP7_75t_L g20393 ( 
.A1(n_20226),
.A2(n_4182),
.B1(n_4180),
.B2(n_4181),
.Y(n_20393)
);

NAND5xp2_ASAP7_75t_L g20394 ( 
.A(n_20313),
.B(n_4184),
.C(n_4181),
.D(n_4183),
.E(n_4185),
.Y(n_20394)
);

NAND2xp5_ASAP7_75t_L g20395 ( 
.A(n_20283),
.B(n_4184),
.Y(n_20395)
);

XNOR2x1_ASAP7_75t_L g20396 ( 
.A(n_20233),
.B(n_4185),
.Y(n_20396)
);

OAI22x1_ASAP7_75t_L g20397 ( 
.A1(n_20333),
.A2(n_4188),
.B1(n_4189),
.B2(n_4187),
.Y(n_20397)
);

NAND2xp5_ASAP7_75t_L g20398 ( 
.A(n_20248),
.B(n_4186),
.Y(n_20398)
);

INVx1_ASAP7_75t_L g20399 ( 
.A(n_20280),
.Y(n_20399)
);

AOI311xp33_ASAP7_75t_L g20400 ( 
.A1(n_20266),
.A2(n_4190),
.A3(n_4188),
.B(n_4189),
.C(n_4191),
.Y(n_20400)
);

NOR2x1_ASAP7_75t_L g20401 ( 
.A(n_20227),
.B(n_4190),
.Y(n_20401)
);

INVx2_ASAP7_75t_L g20402 ( 
.A(n_20347),
.Y(n_20402)
);

INVxp67_ASAP7_75t_SL g20403 ( 
.A(n_20243),
.Y(n_20403)
);

OAI22xp5_ASAP7_75t_L g20404 ( 
.A1(n_20294),
.A2(n_4193),
.B1(n_4191),
.B2(n_4192),
.Y(n_20404)
);

OAI221xp5_ASAP7_75t_L g20405 ( 
.A1(n_20317),
.A2(n_4194),
.B1(n_4192),
.B2(n_4193),
.C(n_4195),
.Y(n_20405)
);

INVx1_ASAP7_75t_L g20406 ( 
.A(n_20308),
.Y(n_20406)
);

XNOR2xp5_ASAP7_75t_L g20407 ( 
.A(n_20245),
.B(n_4195),
.Y(n_20407)
);

OAI211xp5_ASAP7_75t_SL g20408 ( 
.A1(n_20273),
.A2(n_4198),
.B(n_4199),
.C(n_4197),
.Y(n_20408)
);

INVx1_ASAP7_75t_L g20409 ( 
.A(n_20267),
.Y(n_20409)
);

AOI21xp5_ASAP7_75t_L g20410 ( 
.A1(n_20238),
.A2(n_4196),
.B(n_4198),
.Y(n_20410)
);

INVxp67_ASAP7_75t_L g20411 ( 
.A(n_20303),
.Y(n_20411)
);

INVx2_ASAP7_75t_L g20412 ( 
.A(n_20279),
.Y(n_20412)
);

INVx1_ASAP7_75t_L g20413 ( 
.A(n_20276),
.Y(n_20413)
);

AOI22xp5_ASAP7_75t_L g20414 ( 
.A1(n_20234),
.A2(n_4200),
.B1(n_4196),
.B2(n_4199),
.Y(n_20414)
);

BUFx2_ASAP7_75t_L g20415 ( 
.A(n_20262),
.Y(n_20415)
);

HB1xp67_ASAP7_75t_L g20416 ( 
.A(n_20217),
.Y(n_20416)
);

XOR2xp5_ASAP7_75t_L g20417 ( 
.A(n_20257),
.B(n_4201),
.Y(n_20417)
);

AOI22xp33_ASAP7_75t_L g20418 ( 
.A1(n_20220),
.A2(n_4202),
.B1(n_4200),
.B2(n_4201),
.Y(n_20418)
);

XNOR2x1_ASAP7_75t_L g20419 ( 
.A(n_20235),
.B(n_4202),
.Y(n_20419)
);

INVx1_ASAP7_75t_L g20420 ( 
.A(n_20344),
.Y(n_20420)
);

INVx1_ASAP7_75t_L g20421 ( 
.A(n_20345),
.Y(n_20421)
);

AOI22xp5_ASAP7_75t_L g20422 ( 
.A1(n_20325),
.A2(n_4205),
.B1(n_4203),
.B2(n_4204),
.Y(n_20422)
);

INVxp33_ASAP7_75t_L g20423 ( 
.A(n_20220),
.Y(n_20423)
);

OAI22x1_ASAP7_75t_L g20424 ( 
.A1(n_20334),
.A2(n_4206),
.B1(n_4207),
.B2(n_4204),
.Y(n_20424)
);

INVx1_ASAP7_75t_L g20425 ( 
.A(n_20336),
.Y(n_20425)
);

NAND2xp5_ASAP7_75t_L g20426 ( 
.A(n_20240),
.B(n_4203),
.Y(n_20426)
);

OR5x1_ASAP7_75t_L g20427 ( 
.A(n_20260),
.B(n_4208),
.C(n_4206),
.D(n_4207),
.E(n_4209),
.Y(n_20427)
);

AOI211xp5_ASAP7_75t_SL g20428 ( 
.A1(n_20263),
.A2(n_4211),
.B(n_4212),
.C(n_4210),
.Y(n_20428)
);

XNOR2xp5_ASAP7_75t_L g20429 ( 
.A(n_20277),
.B(n_4209),
.Y(n_20429)
);

HB1xp67_ASAP7_75t_L g20430 ( 
.A(n_20246),
.Y(n_20430)
);

INVx1_ASAP7_75t_L g20431 ( 
.A(n_20307),
.Y(n_20431)
);

NAND2xp5_ASAP7_75t_L g20432 ( 
.A(n_20316),
.B(n_20322),
.Y(n_20432)
);

AOI221xp5_ASAP7_75t_L g20433 ( 
.A1(n_20372),
.A2(n_20224),
.B1(n_20220),
.B2(n_20301),
.C(n_20329),
.Y(n_20433)
);

INVx1_ASAP7_75t_L g20434 ( 
.A(n_20371),
.Y(n_20434)
);

NAND4xp75_ASAP7_75t_L g20435 ( 
.A(n_20425),
.B(n_20261),
.C(n_20286),
.D(n_20258),
.Y(n_20435)
);

OAI22xp5_ASAP7_75t_L g20436 ( 
.A1(n_20375),
.A2(n_20335),
.B1(n_20306),
.B2(n_20224),
.Y(n_20436)
);

OAI21xp5_ASAP7_75t_L g20437 ( 
.A1(n_20423),
.A2(n_20324),
.B(n_20311),
.Y(n_20437)
);

NAND2xp5_ASAP7_75t_SL g20438 ( 
.A(n_20420),
.B(n_20224),
.Y(n_20438)
);

INVx1_ASAP7_75t_L g20439 ( 
.A(n_20395),
.Y(n_20439)
);

INVx4_ASAP7_75t_L g20440 ( 
.A(n_20359),
.Y(n_20440)
);

NAND2xp5_ASAP7_75t_L g20441 ( 
.A(n_20364),
.B(n_20270),
.Y(n_20441)
);

AOI32xp33_ASAP7_75t_L g20442 ( 
.A1(n_20415),
.A2(n_20237),
.A3(n_20287),
.B1(n_20309),
.B2(n_20314),
.Y(n_20442)
);

NOR2x1p5_ASAP7_75t_L g20443 ( 
.A(n_20403),
.B(n_20315),
.Y(n_20443)
);

OA21x2_ASAP7_75t_L g20444 ( 
.A1(n_20390),
.A2(n_20399),
.B(n_20368),
.Y(n_20444)
);

XNOR2xp5_ASAP7_75t_L g20445 ( 
.A(n_20377),
.B(n_20275),
.Y(n_20445)
);

AOI211xp5_ASAP7_75t_SL g20446 ( 
.A1(n_20430),
.A2(n_20328),
.B(n_20265),
.C(n_20337),
.Y(n_20446)
);

OAI221xp5_ASAP7_75t_L g20447 ( 
.A1(n_20405),
.A2(n_20225),
.B1(n_20231),
.B2(n_20252),
.C(n_20332),
.Y(n_20447)
);

AOI322xp5_ASAP7_75t_L g20448 ( 
.A1(n_20416),
.A2(n_20264),
.A3(n_20290),
.B1(n_20216),
.B2(n_20330),
.C1(n_20298),
.C2(n_20274),
.Y(n_20448)
);

OAI22xp5_ASAP7_75t_L g20449 ( 
.A1(n_20411),
.A2(n_20305),
.B1(n_20293),
.B2(n_20300),
.Y(n_20449)
);

NAND5xp2_ASAP7_75t_L g20450 ( 
.A(n_20385),
.B(n_20241),
.C(n_20255),
.D(n_20256),
.E(n_20268),
.Y(n_20450)
);

INVx2_ASAP7_75t_L g20451 ( 
.A(n_20396),
.Y(n_20451)
);

NAND3xp33_ASAP7_75t_L g20452 ( 
.A(n_20421),
.B(n_20236),
.C(n_20269),
.Y(n_20452)
);

O2A1O1Ixp33_ASAP7_75t_L g20453 ( 
.A1(n_20432),
.A2(n_20229),
.B(n_20288),
.C(n_20281),
.Y(n_20453)
);

AOI21xp33_ASAP7_75t_L g20454 ( 
.A1(n_20431),
.A2(n_20413),
.B(n_20412),
.Y(n_20454)
);

XNOR2xp5_ASAP7_75t_L g20455 ( 
.A(n_20427),
.B(n_20297),
.Y(n_20455)
);

AOI221xp5_ASAP7_75t_L g20456 ( 
.A1(n_20404),
.A2(n_20236),
.B1(n_20320),
.B2(n_20242),
.C(n_20323),
.Y(n_20456)
);

NAND4xp25_ASAP7_75t_L g20457 ( 
.A(n_20374),
.B(n_20230),
.C(n_20271),
.D(n_20354),
.Y(n_20457)
);

INVx1_ASAP7_75t_L g20458 ( 
.A(n_20387),
.Y(n_20458)
);

AOI211x1_ASAP7_75t_L g20459 ( 
.A1(n_20426),
.A2(n_20271),
.B(n_20321),
.C(n_20319),
.Y(n_20459)
);

AOI221x1_ASAP7_75t_L g20460 ( 
.A1(n_20360),
.A2(n_20236),
.B1(n_20272),
.B2(n_20285),
.C(n_20251),
.Y(n_20460)
);

NAND4xp25_ASAP7_75t_L g20461 ( 
.A(n_20400),
.B(n_20282),
.C(n_20284),
.D(n_20299),
.Y(n_20461)
);

OR2x2_ASAP7_75t_L g20462 ( 
.A(n_20394),
.B(n_20318),
.Y(n_20462)
);

OAI221xp5_ASAP7_75t_L g20463 ( 
.A1(n_20398),
.A2(n_20279),
.B1(n_4212),
.B2(n_4210),
.C(n_4211),
.Y(n_20463)
);

INVx1_ASAP7_75t_L g20464 ( 
.A(n_20362),
.Y(n_20464)
);

AOI221x1_ASAP7_75t_L g20465 ( 
.A1(n_20365),
.A2(n_4215),
.B1(n_4213),
.B2(n_4214),
.C(n_4216),
.Y(n_20465)
);

INVx1_ASAP7_75t_L g20466 ( 
.A(n_20376),
.Y(n_20466)
);

OAI22xp33_ASAP7_75t_L g20467 ( 
.A1(n_20357),
.A2(n_4216),
.B1(n_4213),
.B2(n_4214),
.Y(n_20467)
);

XNOR2x2_ASAP7_75t_L g20468 ( 
.A(n_20382),
.B(n_4217),
.Y(n_20468)
);

BUFx12f_ASAP7_75t_L g20469 ( 
.A(n_20384),
.Y(n_20469)
);

NOR2xp33_ASAP7_75t_L g20470 ( 
.A(n_20373),
.B(n_4217),
.Y(n_20470)
);

INVx1_ASAP7_75t_L g20471 ( 
.A(n_20356),
.Y(n_20471)
);

AND3x4_ASAP7_75t_L g20472 ( 
.A(n_20402),
.B(n_20401),
.C(n_20361),
.Y(n_20472)
);

OAI21xp33_ASAP7_75t_L g20473 ( 
.A1(n_20388),
.A2(n_4218),
.B(n_4219),
.Y(n_20473)
);

AND3x4_ASAP7_75t_L g20474 ( 
.A(n_20409),
.B(n_4218),
.C(n_4219),
.Y(n_20474)
);

OAI221xp5_ASAP7_75t_L g20475 ( 
.A1(n_20370),
.A2(n_4222),
.B1(n_4220),
.B2(n_4221),
.C(n_4223),
.Y(n_20475)
);

A2O1A1Ixp33_ASAP7_75t_SL g20476 ( 
.A1(n_20381),
.A2(n_20386),
.B(n_20369),
.C(n_20406),
.Y(n_20476)
);

INVx1_ASAP7_75t_L g20477 ( 
.A(n_20419),
.Y(n_20477)
);

AOI21xp33_ASAP7_75t_L g20478 ( 
.A1(n_20408),
.A2(n_4220),
.B(n_4221),
.Y(n_20478)
);

OR2x2_ASAP7_75t_L g20479 ( 
.A(n_20363),
.B(n_4224),
.Y(n_20479)
);

INVx3_ASAP7_75t_L g20480 ( 
.A(n_20383),
.Y(n_20480)
);

INVx1_ASAP7_75t_L g20481 ( 
.A(n_20379),
.Y(n_20481)
);

AOI322xp5_ASAP7_75t_L g20482 ( 
.A1(n_20380),
.A2(n_4228),
.A3(n_4227),
.B1(n_4225),
.B2(n_4222),
.C1(n_4224),
.C2(n_4226),
.Y(n_20482)
);

BUFx2_ASAP7_75t_L g20483 ( 
.A(n_20392),
.Y(n_20483)
);

OR2x2_ASAP7_75t_L g20484 ( 
.A(n_20410),
.B(n_4226),
.Y(n_20484)
);

AOI22xp33_ASAP7_75t_SL g20485 ( 
.A1(n_20378),
.A2(n_4228),
.B1(n_4225),
.B2(n_4227),
.Y(n_20485)
);

AOI21xp5_ASAP7_75t_L g20486 ( 
.A1(n_20389),
.A2(n_4231),
.B(n_4230),
.Y(n_20486)
);

AOI22xp5_ASAP7_75t_L g20487 ( 
.A1(n_20391),
.A2(n_4237),
.B1(n_4245),
.B2(n_4229),
.Y(n_20487)
);

OAI22xp5_ASAP7_75t_L g20488 ( 
.A1(n_20366),
.A2(n_4231),
.B1(n_4229),
.B2(n_4230),
.Y(n_20488)
);

HB1xp67_ASAP7_75t_L g20489 ( 
.A(n_20468),
.Y(n_20489)
);

OR2x2_ASAP7_75t_L g20490 ( 
.A(n_20479),
.B(n_20355),
.Y(n_20490)
);

INVx2_ASAP7_75t_L g20491 ( 
.A(n_20474),
.Y(n_20491)
);

INVx1_ASAP7_75t_L g20492 ( 
.A(n_20483),
.Y(n_20492)
);

OAI21xp5_ASAP7_75t_L g20493 ( 
.A1(n_20452),
.A2(n_20428),
.B(n_20429),
.Y(n_20493)
);

INVx1_ASAP7_75t_L g20494 ( 
.A(n_20484),
.Y(n_20494)
);

INVx2_ASAP7_75t_L g20495 ( 
.A(n_20463),
.Y(n_20495)
);

BUFx2_ASAP7_75t_L g20496 ( 
.A(n_20469),
.Y(n_20496)
);

XNOR2xp5_ASAP7_75t_L g20497 ( 
.A(n_20445),
.B(n_20417),
.Y(n_20497)
);

AND2x4_ASAP7_75t_SL g20498 ( 
.A(n_20440),
.B(n_20393),
.Y(n_20498)
);

CKINVDCx20_ASAP7_75t_R g20499 ( 
.A(n_20449),
.Y(n_20499)
);

AOI22xp5_ASAP7_75t_L g20500 ( 
.A1(n_20438),
.A2(n_20407),
.B1(n_20422),
.B2(n_20414),
.Y(n_20500)
);

INVx1_ASAP7_75t_L g20501 ( 
.A(n_20455),
.Y(n_20501)
);

OR5x1_ASAP7_75t_L g20502 ( 
.A(n_20457),
.B(n_20424),
.C(n_20397),
.D(n_20392),
.E(n_20358),
.Y(n_20502)
);

INVx1_ASAP7_75t_L g20503 ( 
.A(n_20480),
.Y(n_20503)
);

OAI22xp5_ASAP7_75t_SL g20504 ( 
.A1(n_20472),
.A2(n_20464),
.B1(n_20471),
.B2(n_20459),
.Y(n_20504)
);

INVx2_ASAP7_75t_L g20505 ( 
.A(n_20443),
.Y(n_20505)
);

INVx1_ASAP7_75t_L g20506 ( 
.A(n_20481),
.Y(n_20506)
);

INVx3_ASAP7_75t_L g20507 ( 
.A(n_20440),
.Y(n_20507)
);

BUFx2_ASAP7_75t_L g20508 ( 
.A(n_20444),
.Y(n_20508)
);

INVx1_ASAP7_75t_L g20509 ( 
.A(n_20444),
.Y(n_20509)
);

INVx1_ASAP7_75t_SL g20510 ( 
.A(n_20462),
.Y(n_20510)
);

OAI221xp5_ASAP7_75t_L g20511 ( 
.A1(n_20442),
.A2(n_20418),
.B1(n_20367),
.B2(n_20358),
.C(n_4234),
.Y(n_20511)
);

NOR4xp25_ASAP7_75t_L g20512 ( 
.A(n_20453),
.B(n_20367),
.C(n_4234),
.D(n_4232),
.Y(n_20512)
);

NAND2xp5_ASAP7_75t_L g20513 ( 
.A(n_20486),
.B(n_4233),
.Y(n_20513)
);

NAND3xp33_ASAP7_75t_L g20514 ( 
.A(n_20446),
.B(n_4232),
.C(n_4233),
.Y(n_20514)
);

INVx1_ASAP7_75t_L g20515 ( 
.A(n_20435),
.Y(n_20515)
);

AO22x2_ASAP7_75t_L g20516 ( 
.A1(n_20436),
.A2(n_4237),
.B1(n_4235),
.B2(n_4236),
.Y(n_20516)
);

AO22x2_ASAP7_75t_L g20517 ( 
.A1(n_20460),
.A2(n_4239),
.B1(n_4236),
.B2(n_4238),
.Y(n_20517)
);

INVx1_ASAP7_75t_L g20518 ( 
.A(n_20441),
.Y(n_20518)
);

INVx1_ASAP7_75t_L g20519 ( 
.A(n_20458),
.Y(n_20519)
);

OAI22xp5_ASAP7_75t_L g20520 ( 
.A1(n_20485),
.A2(n_20487),
.B1(n_20475),
.B2(n_20488),
.Y(n_20520)
);

INVx1_ASAP7_75t_L g20521 ( 
.A(n_20434),
.Y(n_20521)
);

HB1xp67_ASAP7_75t_L g20522 ( 
.A(n_20437),
.Y(n_20522)
);

INVx2_ASAP7_75t_L g20523 ( 
.A(n_20451),
.Y(n_20523)
);

AND3x1_ASAP7_75t_L g20524 ( 
.A(n_20450),
.B(n_4238),
.C(n_4239),
.Y(n_20524)
);

OR5x1_ASAP7_75t_L g20525 ( 
.A(n_20461),
.B(n_20448),
.C(n_20454),
.D(n_20476),
.E(n_20433),
.Y(n_20525)
);

AO22x1_ASAP7_75t_L g20526 ( 
.A1(n_20466),
.A2(n_4242),
.B1(n_4240),
.B2(n_4241),
.Y(n_20526)
);

OAI22xp5_ASAP7_75t_SL g20527 ( 
.A1(n_20447),
.A2(n_4242),
.B1(n_4240),
.B2(n_4241),
.Y(n_20527)
);

XNOR2xp5_ASAP7_75t_L g20528 ( 
.A(n_20456),
.B(n_4243),
.Y(n_20528)
);

OAI21xp5_ASAP7_75t_L g20529 ( 
.A1(n_20477),
.A2(n_4243),
.B(n_4244),
.Y(n_20529)
);

INVx1_ASAP7_75t_L g20530 ( 
.A(n_20439),
.Y(n_20530)
);

AOI21xp5_ASAP7_75t_L g20531 ( 
.A1(n_20478),
.A2(n_4244),
.B(n_4246),
.Y(n_20531)
);

INVx2_ASAP7_75t_L g20532 ( 
.A(n_20470),
.Y(n_20532)
);

INVx1_ASAP7_75t_L g20533 ( 
.A(n_20467),
.Y(n_20533)
);

INVx2_ASAP7_75t_L g20534 ( 
.A(n_20482),
.Y(n_20534)
);

INVx2_ASAP7_75t_L g20535 ( 
.A(n_20473),
.Y(n_20535)
);

AOI31xp33_ASAP7_75t_L g20536 ( 
.A1(n_20465),
.A2(n_4254),
.A3(n_4262),
.B(n_4246),
.Y(n_20536)
);

AOI22xp5_ASAP7_75t_L g20537 ( 
.A1(n_20524),
.A2(n_20499),
.B1(n_20504),
.B2(n_20515),
.Y(n_20537)
);

OAI211xp5_ASAP7_75t_L g20538 ( 
.A1(n_20496),
.A2(n_4249),
.B(n_4247),
.C(n_4248),
.Y(n_20538)
);

NAND2xp5_ASAP7_75t_L g20539 ( 
.A(n_20512),
.B(n_4248),
.Y(n_20539)
);

OAI22xp5_ASAP7_75t_L g20540 ( 
.A1(n_20528),
.A2(n_4251),
.B1(n_4249),
.B2(n_4250),
.Y(n_20540)
);

OAI22x1_ASAP7_75t_L g20541 ( 
.A1(n_20500),
.A2(n_4252),
.B1(n_4250),
.B2(n_4251),
.Y(n_20541)
);

AOI22x1_ASAP7_75t_L g20542 ( 
.A1(n_20508),
.A2(n_4261),
.B1(n_4270),
.B2(n_4252),
.Y(n_20542)
);

INVx1_ASAP7_75t_L g20543 ( 
.A(n_20509),
.Y(n_20543)
);

OAI21x1_ASAP7_75t_SL g20544 ( 
.A1(n_20493),
.A2(n_20531),
.B(n_20491),
.Y(n_20544)
);

OAI22x1_ASAP7_75t_L g20545 ( 
.A1(n_20492),
.A2(n_4256),
.B1(n_4253),
.B2(n_4255),
.Y(n_20545)
);

NAND2xp5_ASAP7_75t_L g20546 ( 
.A(n_20522),
.B(n_4253),
.Y(n_20546)
);

INVx1_ASAP7_75t_L g20547 ( 
.A(n_20513),
.Y(n_20547)
);

OAI22xp5_ASAP7_75t_SL g20548 ( 
.A1(n_20525),
.A2(n_4257),
.B1(n_4255),
.B2(n_4256),
.Y(n_20548)
);

INVx2_ASAP7_75t_L g20549 ( 
.A(n_20502),
.Y(n_20549)
);

OAI22xp5_ASAP7_75t_L g20550 ( 
.A1(n_20501),
.A2(n_4259),
.B1(n_4257),
.B2(n_4258),
.Y(n_20550)
);

NAND2xp33_ASAP7_75t_SL g20551 ( 
.A(n_20490),
.B(n_4258),
.Y(n_20551)
);

XNOR2xp5_ASAP7_75t_L g20552 ( 
.A(n_20497),
.B(n_4260),
.Y(n_20552)
);

OAI22xp5_ASAP7_75t_L g20553 ( 
.A1(n_20507),
.A2(n_4263),
.B1(n_4259),
.B2(n_4261),
.Y(n_20553)
);

AOI21xp5_ASAP7_75t_L g20554 ( 
.A1(n_20519),
.A2(n_4263),
.B(n_4264),
.Y(n_20554)
);

INVx1_ASAP7_75t_L g20555 ( 
.A(n_20511),
.Y(n_20555)
);

OA22x2_ASAP7_75t_L g20556 ( 
.A1(n_20505),
.A2(n_4267),
.B1(n_4265),
.B2(n_4266),
.Y(n_20556)
);

INVx1_ASAP7_75t_L g20557 ( 
.A(n_20489),
.Y(n_20557)
);

AOI21x1_ASAP7_75t_L g20558 ( 
.A1(n_20494),
.A2(n_4265),
.B(n_4266),
.Y(n_20558)
);

INVx1_ASAP7_75t_L g20559 ( 
.A(n_20523),
.Y(n_20559)
);

OAI22x1_ASAP7_75t_L g20560 ( 
.A1(n_20518),
.A2(n_4269),
.B1(n_4267),
.B2(n_4268),
.Y(n_20560)
);

INVx1_ASAP7_75t_L g20561 ( 
.A(n_20520),
.Y(n_20561)
);

INVx2_ASAP7_75t_L g20562 ( 
.A(n_20516),
.Y(n_20562)
);

OAI22xp5_ASAP7_75t_L g20563 ( 
.A1(n_20503),
.A2(n_4271),
.B1(n_4268),
.B2(n_4269),
.Y(n_20563)
);

INVx2_ASAP7_75t_L g20564 ( 
.A(n_20514),
.Y(n_20564)
);

OAI22xp5_ASAP7_75t_L g20565 ( 
.A1(n_20510),
.A2(n_4274),
.B1(n_4272),
.B2(n_4273),
.Y(n_20565)
);

AOI22x1_ASAP7_75t_L g20566 ( 
.A1(n_20521),
.A2(n_4280),
.B1(n_4288),
.B2(n_4272),
.Y(n_20566)
);

NAND2xp5_ASAP7_75t_L g20567 ( 
.A(n_20532),
.B(n_4273),
.Y(n_20567)
);

INVx1_ASAP7_75t_L g20568 ( 
.A(n_20498),
.Y(n_20568)
);

OAI22xp33_ASAP7_75t_L g20569 ( 
.A1(n_20536),
.A2(n_4276),
.B1(n_4274),
.B2(n_4275),
.Y(n_20569)
);

AOI311xp33_ASAP7_75t_L g20570 ( 
.A1(n_20506),
.A2(n_4277),
.A3(n_4275),
.B(n_4276),
.C(n_4278),
.Y(n_20570)
);

OAI22xp5_ASAP7_75t_L g20571 ( 
.A1(n_20530),
.A2(n_4280),
.B1(n_4277),
.B2(n_4279),
.Y(n_20571)
);

OAI22xp5_ASAP7_75t_SL g20572 ( 
.A1(n_20533),
.A2(n_20534),
.B1(n_20495),
.B2(n_20535),
.Y(n_20572)
);

OAI22xp5_ASAP7_75t_L g20573 ( 
.A1(n_20527),
.A2(n_4283),
.B1(n_4281),
.B2(n_4282),
.Y(n_20573)
);

NAND4xp25_ASAP7_75t_SL g20574 ( 
.A(n_20539),
.B(n_20529),
.C(n_20517),
.D(n_20526),
.Y(n_20574)
);

INVx1_ASAP7_75t_L g20575 ( 
.A(n_20548),
.Y(n_20575)
);

OAI22xp5_ASAP7_75t_SL g20576 ( 
.A1(n_20572),
.A2(n_20517),
.B1(n_4283),
.B2(n_4284),
.Y(n_20576)
);

OAI22x1_ASAP7_75t_L g20577 ( 
.A1(n_20537),
.A2(n_4285),
.B1(n_4281),
.B2(n_4282),
.Y(n_20577)
);

NAND4xp25_ASAP7_75t_L g20578 ( 
.A(n_20559),
.B(n_4287),
.C(n_4285),
.D(n_4286),
.Y(n_20578)
);

AOI211xp5_ASAP7_75t_L g20579 ( 
.A1(n_20557),
.A2(n_4289),
.B(n_4287),
.C(n_4288),
.Y(n_20579)
);

AOI22xp5_ASAP7_75t_L g20580 ( 
.A1(n_20568),
.A2(n_4291),
.B1(n_4289),
.B2(n_4290),
.Y(n_20580)
);

A2O1A1Ixp33_ASAP7_75t_L g20581 ( 
.A1(n_20543),
.A2(n_4292),
.B(n_4290),
.C(n_4291),
.Y(n_20581)
);

AND3x2_ASAP7_75t_L g20582 ( 
.A(n_20549),
.B(n_4292),
.C(n_4293),
.Y(n_20582)
);

AOI21xp33_ASAP7_75t_L g20583 ( 
.A1(n_20561),
.A2(n_20562),
.B(n_20547),
.Y(n_20583)
);

AOI22xp33_ASAP7_75t_L g20584 ( 
.A1(n_20564),
.A2(n_4296),
.B1(n_4294),
.B2(n_4295),
.Y(n_20584)
);

AOI22xp5_ASAP7_75t_L g20585 ( 
.A1(n_20551),
.A2(n_4296),
.B1(n_4294),
.B2(n_4295),
.Y(n_20585)
);

AOI22xp33_ASAP7_75t_L g20586 ( 
.A1(n_20555),
.A2(n_4300),
.B1(n_4297),
.B2(n_4298),
.Y(n_20586)
);

OAI22xp5_ASAP7_75t_SL g20587 ( 
.A1(n_20544),
.A2(n_4301),
.B1(n_4302),
.B2(n_4298),
.Y(n_20587)
);

OAI22xp5_ASAP7_75t_L g20588 ( 
.A1(n_20569),
.A2(n_4302),
.B1(n_4297),
.B2(n_4301),
.Y(n_20588)
);

OAI22xp5_ASAP7_75t_L g20589 ( 
.A1(n_20573),
.A2(n_20540),
.B1(n_20554),
.B2(n_20542),
.Y(n_20589)
);

NOR4xp25_ASAP7_75t_L g20590 ( 
.A(n_20570),
.B(n_4305),
.C(n_4303),
.D(n_4304),
.Y(n_20590)
);

AOI222xp33_ASAP7_75t_L g20591 ( 
.A1(n_20550),
.A2(n_4305),
.B1(n_4308),
.B2(n_4303),
.C1(n_4304),
.C2(n_4306),
.Y(n_20591)
);

INVx1_ASAP7_75t_L g20592 ( 
.A(n_20552),
.Y(n_20592)
);

OR5x1_ASAP7_75t_L g20593 ( 
.A(n_20538),
.B(n_4309),
.C(n_4306),
.D(n_4308),
.E(n_4310),
.Y(n_20593)
);

NAND2xp5_ASAP7_75t_L g20594 ( 
.A(n_20565),
.B(n_4309),
.Y(n_20594)
);

AOI22xp5_ASAP7_75t_L g20595 ( 
.A1(n_20553),
.A2(n_4312),
.B1(n_4310),
.B2(n_4311),
.Y(n_20595)
);

NAND4xp25_ASAP7_75t_L g20596 ( 
.A(n_20563),
.B(n_4313),
.C(n_4311),
.D(n_4312),
.Y(n_20596)
);

INVx1_ASAP7_75t_L g20597 ( 
.A(n_20575),
.Y(n_20597)
);

AOI21xp5_ASAP7_75t_L g20598 ( 
.A1(n_20583),
.A2(n_20541),
.B(n_20571),
.Y(n_20598)
);

AOI21xp33_ASAP7_75t_L g20599 ( 
.A1(n_20592),
.A2(n_20589),
.B(n_20594),
.Y(n_20599)
);

OAI22xp5_ASAP7_75t_L g20600 ( 
.A1(n_20576),
.A2(n_20595),
.B1(n_20588),
.B2(n_20585),
.Y(n_20600)
);

NAND2xp5_ASAP7_75t_L g20601 ( 
.A(n_20590),
.B(n_20566),
.Y(n_20601)
);

AOI21xp5_ASAP7_75t_L g20602 ( 
.A1(n_20574),
.A2(n_20545),
.B(n_20560),
.Y(n_20602)
);

AOI21xp5_ASAP7_75t_L g20603 ( 
.A1(n_20596),
.A2(n_20556),
.B(n_20546),
.Y(n_20603)
);

INVx1_ASAP7_75t_L g20604 ( 
.A(n_20582),
.Y(n_20604)
);

XNOR2x1_ASAP7_75t_L g20605 ( 
.A(n_20593),
.B(n_20558),
.Y(n_20605)
);

AOI22xp5_ASAP7_75t_L g20606 ( 
.A1(n_20591),
.A2(n_20567),
.B1(n_4315),
.B2(n_4313),
.Y(n_20606)
);

OAI21xp33_ASAP7_75t_L g20607 ( 
.A1(n_20581),
.A2(n_4314),
.B(n_4316),
.Y(n_20607)
);

XNOR2x1_ASAP7_75t_L g20608 ( 
.A(n_20577),
.B(n_20580),
.Y(n_20608)
);

OAI21xp5_ASAP7_75t_L g20609 ( 
.A1(n_20579),
.A2(n_4314),
.B(n_4316),
.Y(n_20609)
);

INVx1_ASAP7_75t_L g20610 ( 
.A(n_20587),
.Y(n_20610)
);

OAI22xp5_ASAP7_75t_SL g20611 ( 
.A1(n_20586),
.A2(n_4319),
.B1(n_4317),
.B2(n_4318),
.Y(n_20611)
);

AOI21xp5_ASAP7_75t_L g20612 ( 
.A1(n_20584),
.A2(n_4319),
.B(n_4320),
.Y(n_20612)
);

INVx2_ASAP7_75t_L g20613 ( 
.A(n_20578),
.Y(n_20613)
);

OAI22x1_ASAP7_75t_L g20614 ( 
.A1(n_20575),
.A2(n_4323),
.B1(n_4321),
.B2(n_4322),
.Y(n_20614)
);

AOI22xp5_ASAP7_75t_L g20615 ( 
.A1(n_20576),
.A2(n_4323),
.B1(n_4321),
.B2(n_4322),
.Y(n_20615)
);

AOI221xp5_ASAP7_75t_L g20616 ( 
.A1(n_20599),
.A2(n_20597),
.B1(n_20600),
.B2(n_20602),
.C(n_20598),
.Y(n_20616)
);

AOI22xp5_ASAP7_75t_L g20617 ( 
.A1(n_20613),
.A2(n_4326),
.B1(n_4324),
.B2(n_4325),
.Y(n_20617)
);

OAI211xp5_ASAP7_75t_L g20618 ( 
.A1(n_20604),
.A2(n_4326),
.B(n_4324),
.C(n_4325),
.Y(n_20618)
);

AND2x2_ASAP7_75t_L g20619 ( 
.A(n_20610),
.B(n_4327),
.Y(n_20619)
);

AOI21xp5_ASAP7_75t_L g20620 ( 
.A1(n_20608),
.A2(n_4329),
.B(n_4328),
.Y(n_20620)
);

AOI22xp5_ASAP7_75t_L g20621 ( 
.A1(n_20607),
.A2(n_4329),
.B1(n_4327),
.B2(n_4328),
.Y(n_20621)
);

NAND2x1p5_ASAP7_75t_L g20622 ( 
.A(n_20605),
.B(n_4330),
.Y(n_20622)
);

OAI21xp5_ASAP7_75t_L g20623 ( 
.A1(n_20603),
.A2(n_20601),
.B(n_20606),
.Y(n_20623)
);

OAI21xp5_ASAP7_75t_SL g20624 ( 
.A1(n_20612),
.A2(n_4330),
.B(n_4331),
.Y(n_20624)
);

AOI21xp5_ASAP7_75t_L g20625 ( 
.A1(n_20609),
.A2(n_4333),
.B(n_4332),
.Y(n_20625)
);

AOI22xp5_ASAP7_75t_L g20626 ( 
.A1(n_20611),
.A2(n_4333),
.B1(n_4331),
.B2(n_4332),
.Y(n_20626)
);

AOI21xp5_ASAP7_75t_L g20627 ( 
.A1(n_20615),
.A2(n_4336),
.B(n_4335),
.Y(n_20627)
);

XNOR2xp5_ASAP7_75t_L g20628 ( 
.A(n_20616),
.B(n_20614),
.Y(n_20628)
);

NAND4xp25_ASAP7_75t_L g20629 ( 
.A(n_20623),
.B(n_4336),
.C(n_4334),
.D(n_4335),
.Y(n_20629)
);

XNOR2xp5_ASAP7_75t_L g20630 ( 
.A(n_20627),
.B(n_4334),
.Y(n_20630)
);

AOI22xp33_ASAP7_75t_L g20631 ( 
.A1(n_20625),
.A2(n_4339),
.B1(n_4337),
.B2(n_4338),
.Y(n_20631)
);

O2A1O1Ixp33_ASAP7_75t_L g20632 ( 
.A1(n_20624),
.A2(n_4339),
.B(n_4337),
.C(n_4338),
.Y(n_20632)
);

OR2x6_ASAP7_75t_L g20633 ( 
.A(n_20628),
.B(n_20622),
.Y(n_20633)
);

OR2x6_ASAP7_75t_L g20634 ( 
.A(n_20632),
.B(n_20630),
.Y(n_20634)
);

AOI22xp33_ASAP7_75t_SL g20635 ( 
.A1(n_20633),
.A2(n_20620),
.B1(n_20618),
.B2(n_20631),
.Y(n_20635)
);

AOI22xp33_ASAP7_75t_SL g20636 ( 
.A1(n_20634),
.A2(n_20626),
.B1(n_20619),
.B2(n_20621),
.Y(n_20636)
);

AOI21xp5_ASAP7_75t_L g20637 ( 
.A1(n_20636),
.A2(n_20629),
.B(n_20617),
.Y(n_20637)
);

NAND2xp5_ASAP7_75t_L g20638 ( 
.A(n_20635),
.B(n_4340),
.Y(n_20638)
);

INVx1_ASAP7_75t_L g20639 ( 
.A(n_20637),
.Y(n_20639)
);

NAND2x1_ASAP7_75t_SL g20640 ( 
.A(n_20639),
.B(n_20638),
.Y(n_20640)
);

OAI21x1_ASAP7_75t_L g20641 ( 
.A1(n_20639),
.A2(n_4340),
.B(n_4341),
.Y(n_20641)
);

AOI22xp5_ASAP7_75t_L g20642 ( 
.A1(n_20640),
.A2(n_4343),
.B1(n_4341),
.B2(n_4342),
.Y(n_20642)
);

AOI21xp5_ASAP7_75t_L g20643 ( 
.A1(n_20642),
.A2(n_20641),
.B(n_4342),
.Y(n_20643)
);

AOI211xp5_ASAP7_75t_L g20644 ( 
.A1(n_20643),
.A2(n_4345),
.B(n_4343),
.C(n_4344),
.Y(n_20644)
);


endmodule