module fake_jpeg_10768_n_589 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_589);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_60),
.B(n_82),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g174 ( 
.A(n_64),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_67),
.B(n_103),
.Y(n_150)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_77),
.Y(n_197)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_25),
.B(n_16),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_84),
.Y(n_161)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_89),
.Y(n_172)
);

BUFx2_ASAP7_75t_R g90 ( 
.A(n_19),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_90),
.Y(n_139)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_40),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_106),
.Y(n_124)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_96),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_40),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_36),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_20),
.B(n_2),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_31),
.B(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_117),
.Y(n_141)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_112),
.B(n_115),
.Y(n_181)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_33),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_118),
.Y(n_134)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_119),
.B(n_4),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_53),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_42),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_32),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_122),
.B(n_131),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_58),
.A2(n_50),
.B1(n_53),
.B2(n_52),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_127),
.A2(n_129),
.B1(n_153),
.B2(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_128),
.B(n_160),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_76),
.A2(n_85),
.B1(n_102),
.B2(n_113),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_57),
.B(n_52),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_133),
.B(n_144),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_35),
.B1(n_51),
.B2(n_49),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_143),
.A2(n_22),
.B1(n_27),
.B2(n_36),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_185),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_100),
.A2(n_53),
.B1(n_46),
.B2(n_44),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_118),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_64),
.B(n_32),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_35),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_59),
.B(n_49),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_68),
.A2(n_46),
.B1(n_44),
.B2(n_42),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_173),
.A2(n_196),
.B1(n_41),
.B2(n_27),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_61),
.B(n_51),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_62),
.B(n_48),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_65),
.B(n_48),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_116),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_93),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_78),
.A2(n_88),
.B1(n_86),
.B2(n_77),
.Y(n_196)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_134),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_200),
.Y(n_302)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_202),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_204),
.Y(n_304)
);

CKINVDCx12_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_205),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_73),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_207),
.B(n_226),
.Y(n_295)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_211),
.Y(n_297)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_212),
.Y(n_315)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_83),
.B1(n_79),
.B2(n_95),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_214),
.A2(n_228),
.B1(n_265),
.B2(n_179),
.Y(n_292)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_215),
.Y(n_298)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_216),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_217),
.B(n_241),
.Y(n_308)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

BUFx2_ASAP7_75t_SL g290 ( 
.A(n_218),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_224),
.B(n_227),
.Y(n_273)
);

CKINVDCx9p33_ASAP7_75t_R g225 ( 
.A(n_139),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_120),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_22),
.Y(n_227)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

CKINVDCx12_ASAP7_75t_R g234 ( 
.A(n_181),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_234),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_141),
.B(n_124),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_240),
.Y(n_279)
);

INVx4_ASAP7_75t_SL g237 ( 
.A(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_149),
.A2(n_98),
.B1(n_109),
.B2(n_161),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_239),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_162),
.B(n_47),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_137),
.B(n_114),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_145),
.B(n_45),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_242),
.B(n_245),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_181),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_243),
.B(n_244),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_173),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_43),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_266),
.B1(n_225),
.B2(n_154),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_41),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_252),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_127),
.A2(n_89),
.B(n_5),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_261),
.B(n_136),
.Y(n_274)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_135),
.Y(n_249)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_167),
.Y(n_251)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_163),
.B(n_89),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_156),
.B(n_4),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_161),
.C(n_172),
.Y(n_300)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_123),
.Y(n_255)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

BUFx12_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_123),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_122),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_171),
.B1(n_169),
.B2(n_140),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_153),
.A2(n_129),
.B(n_178),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_136),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_264),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_156),
.B(n_5),
.Y(n_265)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_168),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_268),
.A2(n_320),
.B(n_293),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_283),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_281),
.B(n_251),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_210),
.A2(n_171),
.B1(n_192),
.B2(n_154),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_210),
.A2(n_261),
.B1(n_221),
.B2(n_260),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_284),
.A2(n_287),
.B1(n_292),
.B2(n_299),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_248),
.A2(n_132),
.B1(n_168),
.B2(n_179),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_228),
.A2(n_132),
.B1(n_140),
.B2(n_126),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_300),
.B(n_207),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_246),
.A2(n_148),
.B1(n_175),
.B2(n_126),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_241),
.B1(n_202),
.B2(n_262),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_206),
.A2(n_169),
.B1(n_180),
.B2(n_167),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_314),
.B1(n_317),
.B2(n_322),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_203),
.A2(n_246),
.B1(n_198),
.B2(n_239),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_198),
.A2(n_180),
.B1(n_176),
.B2(n_149),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_200),
.A2(n_186),
.B(n_176),
.C(n_8),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_254),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_323),
.A2(n_330),
.B1(n_354),
.B2(n_287),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_351),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_280),
.B(n_235),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_329),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_223),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_326),
.B(n_340),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_327),
.A2(n_290),
.B1(n_282),
.B2(n_229),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_226),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_346),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_274),
.A2(n_266),
.B1(n_256),
.B2(n_213),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx6_ASAP7_75t_SL g334 ( 
.A(n_302),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_334),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_338),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_362),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_201),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_273),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_285),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_344),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_308),
.B(n_208),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_212),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_347),
.Y(n_382)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_267),
.Y(n_348)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_310),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_350),
.Y(n_395)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_300),
.C(n_309),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_295),
.B(n_298),
.C(n_317),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_352),
.B(n_318),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_253),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_360),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_283),
.A2(n_250),
.B1(n_249),
.B2(n_238),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_267),
.B(n_264),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_357),
.Y(n_402)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_356),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_304),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_270),
.B(n_219),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_270),
.B(n_186),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_359),
.B(n_361),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_296),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_277),
.B(n_218),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_272),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_364),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_233),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_278),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_365),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_339),
.A2(n_333),
.B1(n_338),
.B2(n_353),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_378),
.B1(n_380),
.B2(n_387),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_377),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_339),
.A2(n_283),
.B1(n_303),
.B2(n_281),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_343),
.A2(n_283),
.B1(n_320),
.B2(n_305),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_379),
.A2(n_222),
.B1(n_231),
.B2(n_276),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_352),
.A2(n_305),
.B1(n_286),
.B2(n_277),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_328),
.A2(n_286),
.B1(n_275),
.B2(n_306),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_326),
.A2(n_275),
.B1(n_306),
.B2(n_269),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_388),
.A2(n_398),
.B1(n_401),
.B2(n_387),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_334),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_389),
.B(n_349),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_324),
.C(n_348),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_341),
.A2(n_293),
.B(n_319),
.C(n_318),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_361),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_341),
.A2(n_319),
.B(n_297),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_397),
.B(n_400),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_341),
.A2(n_297),
.B(n_294),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_346),
.A2(n_301),
.B(n_289),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_271),
.B1(n_230),
.B2(n_199),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_377),
.A2(n_344),
.B1(n_330),
.B2(n_351),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_404),
.A2(n_428),
.B1(n_430),
.B2(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_405),
.Y(n_443)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

MAJx2_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_367),
.C(n_380),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_385),
.B(n_325),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_408),
.B(n_415),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_409),
.B(n_411),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_360),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_412),
.A2(n_433),
.B(n_434),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_390),
.B(n_331),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_427),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_365),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_402),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_384),
.Y(n_457)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_340),
.Y(n_418)
);

AO22x1_ASAP7_75t_L g460 ( 
.A1(n_418),
.A2(n_431),
.B1(n_429),
.B2(n_412),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_363),
.Y(n_420)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_378),
.A2(n_362),
.B1(n_332),
.B2(n_345),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_425),
.B1(n_438),
.B2(n_395),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_394),
.A2(n_347),
.B(n_356),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_426),
.B(n_429),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_350),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_423),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_396),
.A2(n_329),
.B1(n_282),
.B2(n_289),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_397),
.A2(n_294),
.B(n_321),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_329),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_383),
.A2(n_255),
.B(n_329),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_379),
.A2(n_291),
.B1(n_276),
.B2(n_237),
.Y(n_430)
);

OR2x4_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_257),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_370),
.A2(n_291),
.B1(n_257),
.B2(n_9),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_15),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_400),
.A2(n_7),
.B(n_8),
.Y(n_434)
);

CKINVDCx12_ASAP7_75t_R g435 ( 
.A(n_399),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_435),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_384),
.Y(n_436)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_9),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_399),
.Y(n_445)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_445),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_419),
.A2(n_383),
.B1(n_371),
.B2(n_372),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_444),
.A2(n_433),
.B1(n_428),
.B2(n_430),
.Y(n_483)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_465),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_407),
.B(n_391),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_468),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_457),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_410),
.A2(n_368),
.B(n_395),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_458),
.A2(n_410),
.B(n_405),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_416),
.A2(n_368),
.B1(n_371),
.B2(n_386),
.Y(n_459)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_459),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_L g495 ( 
.A1(n_460),
.A2(n_382),
.B(n_374),
.C(n_381),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_420),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_461),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_414),
.Y(n_470)
);

AOI21xp33_ASAP7_75t_L g463 ( 
.A1(n_404),
.A2(n_367),
.B(n_366),
.Y(n_463)
);

AOI21xp33_ASAP7_75t_L g493 ( 
.A1(n_463),
.A2(n_366),
.B(n_433),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_413),
.B(n_386),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_411),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_391),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_418),
.B(n_366),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_452),
.C(n_450),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_487),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_440),
.A2(n_419),
.B1(n_424),
.B2(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_440),
.A2(n_419),
.B1(n_424),
.B2(n_423),
.Y(n_472)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_456),
.A2(n_408),
.B1(n_438),
.B2(n_437),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_475),
.A2(n_460),
.B(n_442),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_449),
.B(n_409),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_476),
.B(n_439),
.Y(n_511)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_427),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_480),
.Y(n_497)
);

XOR2x2_ASAP7_75t_SL g480 ( 
.A(n_469),
.B(n_444),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_415),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_481),
.B(n_489),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_483),
.A2(n_488),
.B1(n_494),
.B2(n_464),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_456),
.A2(n_434),
.B1(n_431),
.B2(n_433),
.Y(n_484)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_484),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_433),
.B1(n_401),
.B2(n_431),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_422),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_443),
.B(n_373),
.C(n_426),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_441),
.C(n_458),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_493),
.B(n_489),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_455),
.A2(n_398),
.B1(n_381),
.B2(n_432),
.Y(n_494)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_500),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_501),
.B(n_506),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_441),
.C(n_442),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_464),
.C(n_446),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_507),
.B(n_509),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_482),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_511),
.Y(n_523)
);

XOR2x2_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_446),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_514),
.Y(n_519)
);

OAI22x1_ASAP7_75t_SL g513 ( 
.A1(n_488),
.A2(n_451),
.B1(n_453),
.B2(n_461),
.Y(n_513)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_477),
.B(n_465),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_474),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_495),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_451),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_490),
.C(n_481),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_486),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_492),
.B1(n_467),
.B2(n_448),
.Y(n_528)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_520),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_522),
.A2(n_534),
.B1(n_497),
.B2(n_369),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_491),
.C(n_490),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_528),
.Y(n_540)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_510),
.Y(n_527)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_527),
.Y(n_547)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_529),
.B(n_530),
.Y(n_549)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_496),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_499),
.A2(n_485),
.B1(n_483),
.B2(n_494),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_533),
.A2(n_485),
.B1(n_504),
.B2(n_525),
.Y(n_542)
);

XNOR2x1_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_484),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_500),
.A2(n_472),
.B(n_471),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_535),
.A2(n_445),
.B(n_448),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_508),
.B(n_506),
.C(n_498),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_515),
.C(n_508),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_538),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_521),
.A2(n_503),
.B(n_504),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_502),
.C(n_515),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_545),
.Y(n_556)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_542),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_525),
.A2(n_502),
.B1(n_513),
.B2(n_512),
.Y(n_543)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_543),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_544),
.A2(n_520),
.B(n_535),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_497),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_523),
.A2(n_447),
.B1(n_466),
.B2(n_373),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_546),
.B(n_550),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_548),
.B(n_522),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_369),
.C(n_382),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_531),
.A2(n_526),
.B(n_519),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_551),
.B(n_532),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_532),
.C(n_530),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_558),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_557),
.A2(n_552),
.B(n_556),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_540),
.B(n_519),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_539),
.A2(n_526),
.B(n_527),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_560),
.B(n_561),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_562),
.B(n_550),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_537),
.B(n_534),
.C(n_374),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_544),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_565),
.A2(n_554),
.B1(n_561),
.B2(n_13),
.Y(n_578)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_567),
.A2(n_572),
.B(n_549),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_563),
.B(n_545),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_548),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_555),
.B(n_542),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_569),
.B(n_570),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_547),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_545),
.C(n_543),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_560),
.Y(n_575)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_574),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_575),
.B(n_576),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_566),
.Y(n_576)
);

NOR2x1_ASAP7_75t_L g582 ( 
.A(n_577),
.B(n_578),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_573),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_580),
.B(n_564),
.C(n_573),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_581),
.B(n_564),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_583),
.B(n_584),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_579),
.C(n_582),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_586),
.B(n_10),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_11),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_589)
);


endmodule