module fake_jpeg_10160_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx2_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_21),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_17),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_14),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_19),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_60),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_1),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_48),
.C(n_11),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_69),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_73),
.B1(n_74),
.B2(n_15),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_48),
.C(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_26),
.B(n_24),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_45),
.B1(n_19),
.B2(n_23),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_45),
.B1(n_15),
.B2(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_25),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_23),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_55),
.B(n_54),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_57),
.B(n_62),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22x1_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_57),
.B1(n_15),
.B2(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_80),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_54),
.C(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_88),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_15),
.B(n_20),
.C(n_3),
.D(n_4),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_99),
.B(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_66),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_108),
.B1(n_91),
.B2(n_92),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_81),
.C(n_77),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_102),
.C(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_64),
.C(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_87),
.C(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_96),
.B1(n_85),
.B2(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_117),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_96),
.B1(n_99),
.B2(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_114),
.B(n_47),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_76),
.B(n_74),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_26),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_8),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_103),
.C(n_20),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_2),
.B(n_4),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_110),
.C(n_24),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_121),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_7),
.B(n_10),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_7),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_2),
.A3(n_5),
.B1(n_118),
.B2(n_121),
.C1(n_62),
.C2(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_131),
.B(n_125),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_133),
.Y(n_135)
);


endmodule