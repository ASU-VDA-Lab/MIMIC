module fake_netlist_6_832_n_829 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_829);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_829;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_611;
wire n_491;
wire n_772;
wire n_656;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_91),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_7),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_81),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_25),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_35),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_25),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_68),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_50),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_74),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_100),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_16),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_5),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_57),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_77),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_79),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_78),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_31),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_114),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_90),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_53),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_8),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_52),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_71),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_26),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_38),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_19),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_41),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_44),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_148),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_6),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_66),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_22),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_160),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_12),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_73),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_0),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_165),
.B(n_0),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_1),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_166),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_28),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_30),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_164),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_1),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_2),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_32),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_2),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_3),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_3),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

BUFx8_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_33),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_173),
.B(n_4),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_205),
.B(n_208),
.Y(n_267)
);

BUFx8_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_173),
.B(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_212),
.B(n_6),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_211),
.B(n_34),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_226),
.B1(n_171),
.B2(n_172),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_236),
.A2(n_216),
.B1(n_175),
.B2(n_190),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_246),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_200),
.B1(n_227),
.B2(n_222),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_235),
.A2(n_223),
.B1(n_215),
.B2(n_214),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

AO22x2_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_162),
.Y(n_285)
);

OR2x6_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_9),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_213),
.B1(n_210),
.B2(n_207),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_163),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_170),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_237),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_251),
.B1(n_248),
.B2(n_258),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_230),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_240),
.B(n_174),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_203),
.B1(n_201),
.B2(n_199),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_177),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_179),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_230),
.B(n_272),
.Y(n_300)
);

AOI22x1_ASAP7_75t_L g301 ( 
.A1(n_239),
.A2(n_274),
.B1(n_252),
.B2(n_264),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_192),
.B1(n_195),
.B2(n_194),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_240),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_239),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_197),
.B1(n_193),
.B2(n_191),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_182),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_239),
.A2(n_187),
.B1(n_184),
.B2(n_14),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_276),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_238),
.B(n_36),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_274),
.B1(n_264),
.B2(n_270),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_252),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_231),
.B(n_37),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_244),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_264),
.B(n_17),
.Y(n_315)
);

AO22x2_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_250),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_257),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_318)
);

AO22x2_ASAP7_75t_L g319 ( 
.A1(n_256),
.A2(n_27),
.B1(n_42),
.B2(n_43),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g320 ( 
.A1(n_257),
.A2(n_27),
.B1(n_45),
.B2(n_46),
.Y(n_320)
);

AO22x2_ASAP7_75t_L g321 ( 
.A1(n_256),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_321)
);

OR2x6_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_51),
.Y(n_322)
);

NAND3x1_ASAP7_75t_L g323 ( 
.A(n_263),
.B(n_54),
.C(n_55),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_231),
.B(n_233),
.Y(n_324)
);

OR2x6_ASAP7_75t_L g325 ( 
.A(n_229),
.B(n_58),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_229),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_300),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_242),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_315),
.B(n_263),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_242),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_279),
.B(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_243),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_289),
.B(n_243),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_243),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_305),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_311),
.A2(n_261),
.B(n_241),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_243),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_324),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_278),
.B(n_59),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_290),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_60),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_293),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_284),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_308),
.B(n_277),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_302),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_294),
.B(n_241),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

XNOR2x2_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_261),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_287),
.A2(n_241),
.B(n_275),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_275),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_280),
.B(n_263),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_282),
.B(n_249),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_280),
.B(n_247),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_317),
.B(n_231),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_231),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_322),
.B(n_231),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_286),
.B(n_241),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_249),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_286),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_318),
.B(n_247),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_306),
.B(n_233),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_299),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_330),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_336),
.B(n_247),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_336),
.A2(n_241),
.B(n_254),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_247),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_348),
.B(n_228),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_247),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_333),
.B(n_233),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_365),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_329),
.B(n_253),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_352),
.B(n_253),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_363),
.A2(n_260),
.B(n_253),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_332),
.Y(n_422)
);

AND2x2_ASAP7_75t_SL g423 ( 
.A(n_360),
.B(n_377),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_361),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_328),
.B(n_253),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_360),
.B(n_253),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_361),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_356),
.A2(n_241),
.B(n_254),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_396),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_345),
.B(n_260),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_346),
.B(n_260),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_357),
.A2(n_249),
.B(n_254),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_260),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_338),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_358),
.B(n_260),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_393),
.B(n_228),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_386),
.B(n_228),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_381),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_387),
.B(n_228),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_389),
.B(n_232),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_354),
.B(n_268),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_397),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_232),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_232),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_378),
.B(n_232),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_349),
.B(n_350),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_380),
.B(n_232),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_370),
.B(n_249),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_370),
.B(n_249),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_334),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_394),
.A2(n_254),
.B(n_262),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_371),
.B(n_366),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_369),
.B(n_254),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_372),
.B(n_233),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g465 ( 
.A(n_331),
.B(n_62),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_384),
.A2(n_262),
.B(n_233),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_375),
.B(n_262),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_337),
.B(n_268),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_388),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_392),
.B(n_63),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_423),
.B(n_364),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_423),
.B(n_331),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_445),
.Y(n_475)
);

BUFx4f_ASAP7_75t_L g476 ( 
.A(n_465),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_373),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_383),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_431),
.B(n_376),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_376),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_395),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_421),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_413),
.Y(n_487)
);

CKINVDCx6p67_ASAP7_75t_R g488 ( 
.A(n_465),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g489 ( 
.A(n_400),
.B(n_390),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_408),
.B(n_385),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_385),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_416),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_428),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_442),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_417),
.B(n_391),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

INVx6_ASAP7_75t_L g501 ( 
.A(n_470),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g502 ( 
.A(n_413),
.B(n_362),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_461),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_412),
.B(n_382),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_382),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_470),
.B(n_337),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_422),
.B(n_340),
.Y(n_510)
);

BUFx12f_ASAP7_75t_L g511 ( 
.A(n_465),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_471),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_399),
.B(n_410),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_417),
.B(n_268),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_423),
.B(n_340),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_399),
.B(n_364),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_404),
.B(n_364),
.Y(n_522)
);

NAND2x1_ASAP7_75t_L g523 ( 
.A(n_400),
.B(n_64),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_471),
.B(n_410),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_262),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_516),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

BUFx12f_ASAP7_75t_L g531 ( 
.A(n_484),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_410),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_510),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_498),
.B(n_400),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_494),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_514),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_482),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_498),
.B(n_400),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_483),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_521),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_495),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_470),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_479),
.B(n_453),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_496),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_516),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_482),
.Y(n_548)
);

INVx3_ASAP7_75t_SL g549 ( 
.A(n_488),
.Y(n_549)
);

BUFx24_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_516),
.Y(n_551)
);

INVx5_ASAP7_75t_SL g552 ( 
.A(n_516),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_496),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_482),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_524),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_505),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_473),
.Y(n_558)
);

BUFx4f_ASAP7_75t_L g559 ( 
.A(n_492),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_478),
.B(n_469),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_505),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_524),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_505),
.B(n_414),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_480),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_477),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_486),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_505),
.B(n_414),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_501),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_500),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_514),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_504),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

BUFx12f_ASAP7_75t_L g575 ( 
.A(n_531),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_532),
.B(n_545),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_546),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

INVx8_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_534),
.A2(n_518),
.B1(n_502),
.B2(n_476),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_560),
.A2(n_476),
.B1(n_518),
.B2(n_519),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_534),
.A2(n_474),
.B1(n_519),
.B2(n_480),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_564),
.A2(n_472),
.B1(n_525),
.B2(n_511),
.Y(n_583)
);

BUFx12f_ASAP7_75t_L g584 ( 
.A(n_531),
.Y(n_584)
);

OAI22xp33_ASAP7_75t_L g585 ( 
.A1(n_542),
.A2(n_490),
.B1(n_474),
.B2(n_493),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_539),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_570),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_541),
.B(n_493),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_544),
.A2(n_501),
.B1(n_513),
.B2(n_526),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_542),
.A2(n_507),
.B1(n_492),
.B2(n_550),
.Y(n_591)
);

CKINVDCx11_ASAP7_75t_R g592 ( 
.A(n_549),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_549),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_572),
.A2(n_506),
.B1(n_497),
.B2(n_492),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_558),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_571),
.A2(n_507),
.B1(n_492),
.B2(n_448),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_453),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_572),
.A2(n_506),
.B1(n_501),
.B2(n_520),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_558),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_544),
.A2(n_573),
.B1(n_559),
.B2(n_522),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_573),
.A2(n_492),
.B1(n_507),
.B2(n_499),
.Y(n_602)
);

CKINVDCx11_ASAP7_75t_R g603 ( 
.A(n_549),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_SL g604 ( 
.A1(n_571),
.A2(n_507),
.B1(n_403),
.B2(n_520),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_570),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_559),
.A2(n_487),
.B(n_427),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_539),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_574),
.Y(n_609)
);

OAI22xp33_ASAP7_75t_L g610 ( 
.A1(n_559),
.A2(n_503),
.B1(n_458),
.B2(n_449),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_544),
.A2(n_507),
.B1(n_368),
.B2(n_515),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_535),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_529),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_544),
.A2(n_367),
.B(n_454),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_566),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_580),
.A2(n_535),
.B1(n_552),
.B2(n_458),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_595),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_600),
.Y(n_619)
);

BUFx4f_ASAP7_75t_SL g620 ( 
.A(n_575),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_576),
.A2(n_419),
.B1(n_460),
.B2(n_438),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_589),
.B(n_452),
.Y(n_622)
);

OAI21xp33_ASAP7_75t_L g623 ( 
.A1(n_581),
.A2(n_419),
.B(n_460),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_614),
.A2(n_468),
.B(n_403),
.Y(n_624)
);

NAND2x1_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_414),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_588),
.B(n_368),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_581),
.A2(n_460),
.B1(n_438),
.B2(n_433),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_615),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_616),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_606),
.A2(n_414),
.B(n_487),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_611),
.A2(n_468),
.B1(n_450),
.B2(n_569),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_598),
.A2(n_433),
.B1(n_451),
.B2(n_426),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_577),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_582),
.A2(n_552),
.B1(n_569),
.B2(n_449),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_587),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_605),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_591),
.A2(n_552),
.B1(n_569),
.B2(n_449),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_585),
.A2(n_597),
.B1(n_604),
.B2(n_591),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_585),
.A2(n_597),
.B1(n_604),
.B2(n_583),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_583),
.A2(n_552),
.B1(n_569),
.B2(n_427),
.Y(n_641)
);

OAI222xp33_ASAP7_75t_L g642 ( 
.A1(n_599),
.A2(n_509),
.B1(n_567),
.B2(n_446),
.C1(n_418),
.C2(n_401),
.Y(n_642)
);

NOR2x1_ASAP7_75t_L g643 ( 
.A(n_586),
.B(n_529),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_609),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_596),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_592),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_584),
.A2(n_418),
.B1(n_401),
.B2(n_441),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_593),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_594),
.A2(n_436),
.B1(n_439),
.B2(n_540),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_602),
.A2(n_420),
.B(n_429),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_596),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_612),
.A2(n_436),
.B1(n_439),
.B2(n_540),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_613),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_590),
.A2(n_540),
.B1(n_536),
.B2(n_489),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_610),
.A2(n_536),
.B1(n_489),
.B2(n_547),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_601),
.A2(n_451),
.B1(n_426),
.B2(n_420),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_610),
.A2(n_434),
.B1(n_567),
.B2(n_446),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_603),
.A2(n_434),
.B1(n_491),
.B2(n_432),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_613),
.B(n_467),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_613),
.A2(n_434),
.B1(n_432),
.B2(n_444),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_607),
.A2(n_441),
.B1(n_547),
.B2(n_565),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_579),
.A2(n_429),
.B(n_466),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_607),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_579),
.A2(n_444),
.B1(n_447),
.B2(n_443),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_608),
.A2(n_411),
.B(n_425),
.Y(n_665)
);

OAI222xp33_ASAP7_75t_L g666 ( 
.A1(n_608),
.A2(n_553),
.B1(n_543),
.B2(n_533),
.C1(n_455),
.C2(n_523),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_640),
.A2(n_450),
.B1(n_555),
.B2(n_556),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_640),
.A2(n_450),
.B1(n_555),
.B2(n_556),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_624),
.A2(n_551),
.B1(n_562),
.B2(n_565),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_639),
.A2(n_562),
.B1(n_551),
.B2(n_536),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_639),
.A2(n_450),
.B1(n_447),
.B2(n_443),
.Y(n_671)
);

AOI222xp33_ASAP7_75t_L g672 ( 
.A1(n_622),
.A2(n_425),
.B1(n_459),
.B2(n_466),
.C1(n_409),
.C2(n_437),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_623),
.A2(n_406),
.B1(n_409),
.B2(n_440),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_618),
.B(n_574),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_631),
.A2(n_406),
.B1(n_440),
.B2(n_435),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_617),
.A2(n_607),
.B1(n_579),
.B2(n_455),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_658),
.A2(n_607),
.B1(n_557),
.B2(n_563),
.Y(n_677)
);

OAI211xp5_ASAP7_75t_SL g678 ( 
.A1(n_645),
.A2(n_459),
.B(n_437),
.C(n_406),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_L g679 ( 
.A1(n_658),
.A2(n_533),
.B(n_543),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_652),
.A2(n_440),
.B1(n_435),
.B2(n_512),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_621),
.A2(n_568),
.B1(n_563),
.B2(n_530),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_621),
.A2(n_568),
.B1(n_563),
.B2(n_530),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_626),
.A2(n_435),
.B1(n_512),
.B2(n_485),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_627),
.A2(n_568),
.B1(n_530),
.B2(n_554),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_647),
.A2(n_635),
.B1(n_648),
.B2(n_659),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_638),
.A2(n_641),
.B1(n_620),
.B2(n_632),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_620),
.A2(n_481),
.B1(n_485),
.B2(n_527),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_656),
.A2(n_554),
.B1(n_481),
.B2(n_553),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_619),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_654),
.A2(n_561),
.B1(n_548),
.B2(n_539),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_L g691 ( 
.A1(n_650),
.A2(n_632),
.B1(n_656),
.B2(n_665),
.C(n_662),
.Y(n_691)
);

OAI222xp33_ASAP7_75t_L g692 ( 
.A1(n_661),
.A2(n_528),
.B1(n_517),
.B2(n_508),
.C1(n_554),
.C2(n_467),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_655),
.A2(n_630),
.B1(n_649),
.B2(n_651),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_628),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_653),
.A2(n_430),
.B1(n_528),
.B2(n_405),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_664),
.A2(n_430),
.B1(n_405),
.B2(n_407),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_664),
.A2(n_430),
.B1(n_405),
.B2(n_407),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_642),
.B(n_462),
.C(n_463),
.Y(n_698)
);

OAI211xp5_ASAP7_75t_SL g699 ( 
.A1(n_629),
.A2(n_517),
.B(n_508),
.C(n_462),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_660),
.A2(n_430),
.B1(n_407),
.B2(n_548),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_660),
.A2(n_430),
.B1(n_407),
.B2(n_548),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_657),
.A2(n_407),
.B1(n_463),
.B2(n_456),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_633),
.A2(n_634),
.B1(n_636),
.B2(n_637),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_689),
.B(n_657),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_694),
.B(n_644),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_685),
.B(n_646),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_SL g707 ( 
.A(n_669),
.B(n_666),
.C(n_643),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_692),
.B(n_663),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_689),
.B(n_625),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_703),
.B(n_548),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_674),
.B(n_65),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_686),
.B(n_262),
.C(n_548),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_674),
.B(n_693),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_698),
.B(n_561),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_679),
.B(n_561),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_691),
.A2(n_430),
.B1(n_561),
.B2(n_407),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_690),
.B(n_676),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_702),
.B(n_67),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_L g719 ( 
.A1(n_671),
.A2(n_667),
.B1(n_668),
.B2(n_687),
.C(n_679),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_702),
.B(n_688),
.Y(n_720)
);

AOI221xp5_ASAP7_75t_L g721 ( 
.A1(n_678),
.A2(n_457),
.B1(n_456),
.B2(n_561),
.C(n_76),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_675),
.B(n_70),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_670),
.B(n_72),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_672),
.B(n_75),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_700),
.B(n_701),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_699),
.A2(n_407),
.B1(n_457),
.B2(n_83),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_681),
.B(n_80),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_683),
.B(n_82),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_677),
.B(n_84),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_673),
.B(n_85),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_713),
.B(n_704),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_705),
.B(n_680),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_713),
.B(n_682),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_724),
.A2(n_684),
.B1(n_696),
.B2(n_697),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_706),
.B(n_86),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_704),
.B(n_695),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_709),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_717),
.B(n_87),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_721),
.B(n_88),
.C(n_89),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_717),
.B(n_92),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_723),
.B(n_95),
.C(n_96),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_715),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_SL g743 ( 
.A1(n_708),
.A2(n_407),
.B1(n_98),
.B2(n_99),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_727),
.B(n_97),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_727),
.B(n_710),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_712),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_715),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_731),
.B(n_720),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_747),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_742),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_737),
.B(n_720),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_731),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_745),
.B(n_733),
.Y(n_753)
);

XOR2x2_ASAP7_75t_L g754 ( 
.A(n_738),
.B(n_712),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_745),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_745),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_739),
.B(n_729),
.C(n_719),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_733),
.B(n_714),
.Y(n_758)
);

XNOR2xp5_ASAP7_75t_L g759 ( 
.A(n_754),
.B(n_738),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_749),
.Y(n_760)
);

XNOR2x1_ASAP7_75t_L g761 ( 
.A(n_748),
.B(n_740),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_750),
.B(n_751),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_755),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_761),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_753),
.B1(n_758),
.B2(n_757),
.Y(n_765)
);

XNOR2xp5_ASAP7_75t_L g766 ( 
.A(n_759),
.B(n_740),
.Y(n_766)
);

OA22x2_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_752),
.B1(n_756),
.B2(n_763),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_762),
.A2(n_757),
.B1(n_752),
.B2(n_734),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_767),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_765),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_768),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_764),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_770),
.A2(n_766),
.B1(n_736),
.B2(n_735),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_772),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_769),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_774),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_773),
.A2(n_771),
.B1(n_769),
.B2(n_735),
.Y(n_777)
);

AND4x1_ASAP7_75t_L g778 ( 
.A(n_775),
.B(n_741),
.C(n_746),
.D(n_708),
.Y(n_778)
);

OAI22x1_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_744),
.B1(n_718),
.B2(n_711),
.Y(n_779)
);

NOR2x1_ASAP7_75t_L g780 ( 
.A(n_776),
.B(n_744),
.Y(n_780)
);

AOI31xp33_ASAP7_75t_L g781 ( 
.A1(n_777),
.A2(n_743),
.A3(n_744),
.B(n_718),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_777),
.B(n_711),
.Y(n_782)
);

AOI221xp5_ASAP7_75t_L g783 ( 
.A1(n_777),
.A2(n_716),
.B1(n_707),
.B2(n_722),
.C(n_732),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_777),
.B(n_722),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_780),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_779),
.A2(n_784),
.B1(n_782),
.B2(n_783),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_781),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_SL g788 ( 
.A1(n_784),
.A2(n_725),
.B1(n_728),
.B2(n_730),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_779),
.A2(n_725),
.B1(n_726),
.B2(n_106),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_780),
.Y(n_790)
);

OR3x2_ASAP7_75t_L g791 ( 
.A(n_785),
.B(n_104),
.C(n_105),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_787),
.B(n_725),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_786),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.C(n_110),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_790),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_788),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_789),
.Y(n_796)
);

AND4x1_ASAP7_75t_L g797 ( 
.A(n_786),
.B(n_112),
.C(n_115),
.D(n_116),
.Y(n_797)
);

AO22x2_ASAP7_75t_L g798 ( 
.A1(n_787),
.A2(n_725),
.B1(n_119),
.B2(n_120),
.Y(n_798)
);

NOR2x1_ASAP7_75t_L g799 ( 
.A(n_794),
.B(n_117),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_792),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_796),
.B(n_121),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_798),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_798),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_795),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_791),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_797),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_793),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_794),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_794),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_804),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_808),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_SL g812 ( 
.A1(n_802),
.A2(n_128),
.B(n_129),
.C(n_133),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_805),
.A2(n_806),
.B1(n_809),
.B2(n_807),
.Y(n_813)
);

AND4x2_ASAP7_75t_L g814 ( 
.A(n_799),
.B(n_134),
.C(n_135),
.D(n_137),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_808),
.Y(n_815)
);

OAI22x1_ASAP7_75t_L g816 ( 
.A1(n_803),
.A2(n_800),
.B1(n_801),
.B2(n_142),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_815),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_811),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_813),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_816),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_814),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_819),
.A2(n_810),
.B1(n_812),
.B2(n_143),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_817),
.A2(n_138),
.B1(n_141),
.B2(n_144),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_818),
.A2(n_145),
.B1(n_147),
.B2(n_149),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_822),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_825),
.A2(n_821),
.B1(n_820),
.B2(n_823),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_826),
.Y(n_827)
);

AOI221xp5_ASAP7_75t_L g828 ( 
.A1(n_827),
.A2(n_824),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_828)
);

AOI211xp5_ASAP7_75t_L g829 ( 
.A1(n_828),
.A2(n_150),
.B(n_155),
.C(n_156),
.Y(n_829)
);


endmodule