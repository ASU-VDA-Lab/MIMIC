module fake_jpeg_29052_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_62),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_0),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_1),
.Y(n_65)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_53),
.B1(n_49),
.B2(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_75),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_SL g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_20),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_45),
.B1(n_54),
.B2(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_4),
.Y(n_91)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_3),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_6),
.B(n_8),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_5),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_66),
.B(n_26),
.C(n_10),
.D(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_66),
.C(n_27),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_112),
.C(n_19),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_109),
.B1(n_39),
.B2(n_21),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_18),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_112),
.B1(n_92),
.B2(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_72),
.B1(n_80),
.B2(n_24),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_110),
.B1(n_97),
.B2(n_100),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_100),
.A3(n_103),
.B1(n_30),
.B2(n_31),
.C1(n_32),
.C2(n_25),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.C(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_116),
.C(n_126),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

AOI31xp33_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_115),
.A3(n_113),
.B(n_123),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_117),
.Y(n_134)
);


endmodule