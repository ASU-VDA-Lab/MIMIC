module real_aes_16848_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g122 ( .A(n_0), .B(n_123), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_1), .A2(n_34), .B1(n_157), .B2(n_169), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_2), .A2(n_10), .B1(n_535), .B2(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g123 ( .A(n_3), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_4), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_5), .A2(n_11), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_6), .A2(n_842), .B1(n_848), .B2(n_849), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_6), .Y(n_848) );
BUFx2_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
OR2x2_ASAP7_75t_L g137 ( .A(n_7), .B(n_30), .Y(n_137) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_8), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_9), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_12), .B(n_208), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_13), .A2(n_101), .B1(n_205), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_14), .A2(n_31), .B1(n_558), .B2(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_15), .B(n_208), .Y(n_600) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_16), .A2(n_45), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_17), .B(n_297), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_18), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_19), .A2(n_94), .B1(n_846), .B2(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_19), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_20), .A2(n_38), .B1(n_195), .B2(n_213), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_21), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_22), .A2(n_43), .B1(n_195), .B2(n_535), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_23), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_23), .A2(n_82), .B1(n_592), .B2(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_24), .B(n_558), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_25), .B(n_160), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_26), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_27), .B(n_218), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_28), .Y(n_204) );
AOI22x1_ASAP7_75t_L g874 ( .A1(n_29), .A2(n_875), .B1(n_876), .B2(n_878), .Y(n_874) );
INVx1_ASAP7_75t_L g878 ( .A(n_29), .Y(n_878) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_30), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_32), .A2(n_85), .B1(n_157), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_33), .A2(n_37), .B1(n_157), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_35), .A2(n_48), .B1(n_535), .B2(n_537), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_36), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_39), .B(n_208), .Y(n_258) );
INVx2_ASAP7_75t_L g128 ( .A(n_40), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_41), .B(n_209), .Y(n_292) );
INVx1_ASAP7_75t_L g117 ( .A(n_42), .Y(n_117) );
BUFx3_ASAP7_75t_L g136 ( .A(n_42), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_44), .B(n_177), .Y(n_299) );
AND2x2_ASAP7_75t_L g197 ( .A(n_46), .B(n_177), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_47), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_49), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_50), .B(n_213), .Y(n_212) );
XNOR2x1_ASAP7_75t_L g138 ( .A(n_51), .B(n_139), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_51), .A2(n_78), .B1(n_870), .B2(n_871), .Y(n_869) );
INVx1_ASAP7_75t_SL g870 ( .A(n_51), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_52), .A2(n_70), .B1(n_213), .B2(n_537), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_53), .A2(n_73), .B1(n_157), .B2(n_548), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_54), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_55), .A2(n_162), .B(n_187), .C(n_188), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_56), .A2(n_98), .B1(n_535), .B2(n_546), .Y(n_609) );
INVx1_ASAP7_75t_L g153 ( .A(n_57), .Y(n_153) );
AND2x4_ASAP7_75t_L g174 ( .A(n_58), .B(n_175), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_59), .A2(n_60), .B1(n_195), .B2(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_61), .B(n_218), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_62), .A2(n_106), .B1(n_124), .B2(n_887), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_63), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_64), .B(n_177), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_65), .B(n_195), .Y(n_261) );
INVx1_ASAP7_75t_L g175 ( .A(n_66), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_67), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_68), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_69), .B(n_218), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_71), .B(n_157), .Y(n_156) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_72), .B(n_169), .C(n_209), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_74), .B(n_157), .Y(n_239) );
INVx2_ASAP7_75t_L g164 ( .A(n_75), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_76), .B(n_208), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_77), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g871 ( .A(n_78), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_79), .B(n_215), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_80), .A2(n_97), .B1(n_187), .B2(n_195), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_81), .Y(n_574) );
INVx1_ASAP7_75t_L g877 ( .A(n_82), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_83), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g843 ( .A(n_83), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_84), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_86), .A2(n_91), .B1(n_160), .B2(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_87), .B(n_208), .Y(n_207) );
NAND2xp33_ASAP7_75t_SL g231 ( .A(n_88), .B(n_214), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_89), .B(n_206), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_90), .B(n_218), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_92), .Y(n_552) );
INVx1_ASAP7_75t_L g121 ( .A(n_93), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_93), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g846 ( .A(n_94), .Y(n_846) );
NAND2xp33_ASAP7_75t_L g603 ( .A(n_95), .B(n_208), .Y(n_603) );
NAND2xp33_ASAP7_75t_L g240 ( .A(n_96), .B(n_214), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_99), .B(n_177), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g227 ( .A(n_100), .B(n_214), .C(n_226), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_102), .B(n_157), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_103), .B(n_160), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_104), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx8_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx8_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx12f_ASAP7_75t_L g887 ( .A(n_110), .Y(n_887) );
BUFx12f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
AND3x2_ASAP7_75t_L g857 ( .A(n_116), .B(n_120), .C(n_858), .Y(n_857) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g866 ( .A(n_117), .Y(n_866) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_860), .Y(n_124) );
OAI21xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B(n_854), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_127), .Y(n_883) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g862 ( .A(n_128), .B(n_863), .Y(n_862) );
A2O1A1O1Ixp25_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_138), .B(n_520), .C(n_841), .D(n_850), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx2_ASAP7_75t_L g885 ( .A(n_131), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
NOR2x1_ASAP7_75t_R g522 ( .A(n_132), .B(n_523), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g853 ( .A(n_133), .B(n_135), .Y(n_853) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx2_ASAP7_75t_L g523 ( .A(n_135), .Y(n_523) );
NOR2x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g858 ( .A(n_137), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_138), .A2(n_521), .B1(n_885), .B2(n_886), .Y(n_884) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g872 ( .A(n_140), .Y(n_872) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_141), .B(n_415), .Y(n_140) );
NOR2x1_ASAP7_75t_L g141 ( .A(n_142), .B(n_350), .Y(n_141) );
NAND3xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_273), .C(n_323), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_198), .B(n_233), .C(n_250), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g489 ( .A(n_145), .B(n_408), .Y(n_489) );
OR2x2_ASAP7_75t_L g500 ( .A(n_145), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_146), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g391 ( .A(n_146), .B(n_280), .Y(n_391) );
AND2x2_ASAP7_75t_L g512 ( .A(n_146), .B(n_322), .Y(n_512) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_178), .Y(n_146) );
INVx2_ASAP7_75t_L g342 ( .A(n_147), .Y(n_342) );
AND2x2_ASAP7_75t_L g357 ( .A(n_147), .B(n_309), .Y(n_357) );
AND2x2_ASAP7_75t_L g366 ( .A(n_147), .B(n_235), .Y(n_366) );
AND2x2_ASAP7_75t_L g435 ( .A(n_147), .B(n_321), .Y(n_435) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g248 ( .A(n_148), .Y(n_248) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_154), .B(n_176), .Y(n_148) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_149), .A2(n_202), .B(n_217), .Y(n_201) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_149), .A2(n_202), .B(n_217), .Y(n_316) );
OAI21xp33_ASAP7_75t_SL g407 ( .A1(n_149), .A2(n_154), .B(n_176), .Y(n_407) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_150), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_150), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
INVx2_ASAP7_75t_L g272 ( .A(n_151), .Y(n_272) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_165), .B(n_173), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_162), .Y(n_155) );
OAI22xp33_ASAP7_75t_L g193 ( .A1(n_157), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_193) );
INVx1_ASAP7_75t_L g537 ( .A(n_157), .Y(n_537) );
INVx1_ASAP7_75t_L g546 ( .A(n_157), .Y(n_546) );
INVx4_ASAP7_75t_L g548 ( .A(n_157), .Y(n_548) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g161 ( .A(n_158), .Y(n_161) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_158), .Y(n_169) );
INVx1_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
INVx1_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
INVx1_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
INVx1_ASAP7_75t_L g269 ( .A(n_158), .Y(n_269) );
INVx1_ASAP7_75t_L g545 ( .A(n_160), .Y(n_545) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_162), .A2(n_229), .B(n_231), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_162), .A2(n_239), .B(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_162), .A2(n_257), .B(n_258), .Y(n_256) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g172 ( .A(n_164), .Y(n_172) );
BUFx8_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
INVx1_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_170), .Y(n_165) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g192 ( .A(n_171), .Y(n_192) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g216 ( .A(n_172), .Y(n_216) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_173), .A2(n_203), .B(n_210), .Y(n_202) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_173), .A2(n_224), .B(n_228), .Y(n_223) );
AND2x4_ASAP7_75t_SL g245 ( .A(n_173), .B(n_219), .Y(n_245) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_173), .A2(n_256), .B(n_259), .Y(n_255) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_173), .A2(n_291), .B(n_294), .Y(n_290) );
BUFx10_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx10_ASAP7_75t_L g184 ( .A(n_174), .Y(n_184) );
INVx1_ASAP7_75t_L g572 ( .A(n_174), .Y(n_572) );
AND2x2_ASAP7_75t_L g406 ( .A(n_178), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g249 ( .A(n_179), .B(n_221), .Y(n_249) );
INVx2_ASAP7_75t_L g278 ( .A(n_179), .Y(n_278) );
AOI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_185), .B(n_197), .Y(n_179) );
NOR2xp67_ASAP7_75t_SL g180 ( .A(n_181), .B(n_183), .Y(n_180) );
INVx2_ASAP7_75t_L g538 ( .A(n_181), .Y(n_538) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_182), .A2(n_184), .A3(n_264), .B(n_270), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g551 ( .A(n_182), .B(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_182), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g532 ( .A(n_183), .Y(n_532) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AO31x2_ASAP7_75t_L g542 ( .A1(n_184), .A2(n_543), .A3(n_550), .B(n_551), .Y(n_542) );
AO31x2_ASAP7_75t_L g555 ( .A1(n_184), .A2(n_556), .A3(n_562), .B(n_563), .Y(n_555) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_184), .A2(n_619), .A3(n_622), .B(n_623), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_191), .Y(n_185) );
INVx1_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx2_ASAP7_75t_SL g588 ( .A(n_190), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_192), .A2(n_265), .B1(n_267), .B2(n_268), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_192), .A2(n_267), .B1(n_534), .B2(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_192), .A2(n_267), .B1(n_557), .B2(n_560), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_192), .A2(n_267), .B1(n_569), .B2(n_570), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_192), .A2(n_267), .B1(n_620), .B2(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g266 ( .A(n_195), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_195), .A2(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g443 ( .A(n_198), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_220), .Y(n_199) );
INVx1_ASAP7_75t_L g463 ( .A(n_200), .Y(n_463) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g301 ( .A(n_201), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g384 ( .A(n_201), .B(n_289), .Y(n_384) );
O2A1O1Ixp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .C(n_209), .Y(n_203) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_208), .A2(n_225), .B(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g297 ( .A(n_208), .Y(n_297) );
INVx3_ASAP7_75t_L g535 ( .A(n_208), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_209), .A2(n_260), .B(n_261), .Y(n_259) );
INVx6_ASAP7_75t_L g267 ( .A(n_209), .Y(n_267) );
O2A1O1Ixp5_ASAP7_75t_L g598 ( .A1(n_209), .A2(n_548), .B(n_599), .C(n_600), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_215), .Y(n_210) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g558 ( .A(n_214), .Y(n_558) );
INVx2_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_216), .A2(n_242), .B1(n_243), .B2(n_244), .Y(n_241) );
INVx2_ASAP7_75t_L g622 ( .A(n_218), .Y(n_622) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_SL g222 ( .A(n_219), .Y(n_222) );
INVx2_ASAP7_75t_L g254 ( .A(n_219), .Y(n_254) );
BUFx3_ASAP7_75t_L g562 ( .A(n_219), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_219), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g596 ( .A(n_219), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_219), .B(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_219), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g310 ( .A(n_220), .B(n_248), .Y(n_310) );
INVxp67_ASAP7_75t_L g459 ( .A(n_220), .Y(n_459) );
OR2x2_ASAP7_75t_L g501 ( .A(n_220), .B(n_235), .Y(n_501) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g282 ( .A(n_221), .Y(n_282) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_232), .Y(n_221) );
INVx1_ASAP7_75t_L g298 ( .A(n_226), .Y(n_298) );
INVx1_ASAP7_75t_SL g549 ( .A(n_226), .Y(n_549) );
INVx1_ASAP7_75t_L g590 ( .A(n_226), .Y(n_590) );
INVx1_ASAP7_75t_L g559 ( .A(n_230), .Y(n_559) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_246), .Y(n_233) );
INVx1_ASAP7_75t_L g356 ( .A(n_234), .Y(n_356) );
AND2x2_ASAP7_75t_L g510 ( .A(n_234), .B(n_406), .Y(n_510) );
BUFx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g281 ( .A(n_235), .Y(n_281) );
INVx4_ASAP7_75t_L g321 ( .A(n_235), .Y(n_321) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_241), .B(n_245), .Y(n_237) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
AND2x2_ASAP7_75t_L g337 ( .A(n_247), .B(n_320), .Y(n_337) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g374 ( .A(n_248), .B(n_322), .Y(n_374) );
INVx2_ASAP7_75t_L g340 ( .A(n_249), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_249), .B(n_345), .Y(n_508) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_252), .B(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g493 ( .A(n_252), .Y(n_493) );
AND2x2_ASAP7_75t_L g507 ( .A(n_252), .B(n_329), .Y(n_507) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_263), .Y(n_252) );
INVx1_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
AND2x2_ASAP7_75t_L g442 ( .A(n_253), .B(n_349), .Y(n_442) );
OR2x2_ASAP7_75t_L g479 ( .A(n_253), .B(n_263), .Y(n_479) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_262), .Y(n_253) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_254), .A2(n_290), .B(n_299), .Y(n_289) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_254), .A2(n_290), .B(n_299), .Y(n_302) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_254), .A2(n_255), .B(n_262), .Y(n_305) );
AND2x2_ASAP7_75t_L g288 ( .A(n_263), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g303 ( .A(n_263), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g349 ( .A(n_263), .Y(n_349) );
OR2x2_ASAP7_75t_L g362 ( .A(n_263), .B(n_302), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_263), .B(n_302), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_267), .A2(n_544), .B1(n_547), .B2(n_549), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_267), .A2(n_587), .B1(n_589), .B2(n_590), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_267), .A2(n_602), .B(n_603), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_267), .A2(n_549), .B1(n_609), .B2(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g561 ( .A(n_269), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
BUFx2_ASAP7_75t_L g550 ( .A(n_272), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_283), .B(n_306), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI31xp33_ASAP7_75t_L g352 ( .A1(n_275), .A2(n_353), .A3(n_355), .B(n_358), .Y(n_352) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
AND2x2_ASAP7_75t_L g365 ( .A(n_276), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g375 ( .A(n_277), .Y(n_375) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_277), .Y(n_381) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
AND2x2_ASAP7_75t_L g338 ( .A(n_278), .B(n_322), .Y(n_338) );
INVx2_ASAP7_75t_L g388 ( .A(n_278), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_279), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g413 ( .A(n_280), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g462 ( .A(n_280), .B(n_463), .Y(n_462) );
AOI33xp33_ASAP7_75t_L g517 ( .A1(n_280), .A2(n_347), .A3(n_357), .B1(n_384), .B2(n_493), .B3(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
INVx1_ASAP7_75t_L g409 ( .A(n_282), .Y(n_409) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_300), .Y(n_284) );
INVx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
AND2x2_ASAP7_75t_L g398 ( .A(n_285), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g360 ( .A(n_286), .Y(n_360) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g428 ( .A(n_287), .B(n_315), .Y(n_428) );
AND2x2_ASAP7_75t_L g378 ( .A(n_288), .B(n_372), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_288), .B(n_396), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_288), .B(n_428), .Y(n_477) );
AND2x2_ASAP7_75t_L g314 ( .A(n_289), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g333 ( .A(n_289), .B(n_328), .Y(n_333) );
INVx1_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
AOI21x1_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_298), .Y(n_294) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g403 ( .A(n_301), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_301), .B(n_496), .Y(n_498) );
AND2x2_ASAP7_75t_L g511 ( .A(n_301), .B(n_327), .Y(n_511) );
AND2x2_ASAP7_75t_L g329 ( .A(n_302), .B(n_315), .Y(n_329) );
INVx2_ASAP7_75t_L g311 ( .A(n_303), .Y(n_311) );
AND2x2_ASAP7_75t_L g425 ( .A(n_303), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g484 ( .A(n_303), .B(n_396), .Y(n_484) );
BUFx2_ASAP7_75t_L g466 ( .A(n_304), .Y(n_466) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
OAI32xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .A3(n_312), .B1(n_317), .B2(n_318), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g414 ( .A(n_309), .Y(n_414) );
AND2x2_ASAP7_75t_L g444 ( .A(n_309), .B(n_366), .Y(n_444) );
AND2x2_ASAP7_75t_L g386 ( .A(n_310), .B(n_387), .Y(n_386) );
AND3x2_ASAP7_75t_L g393 ( .A(n_310), .B(n_320), .C(n_388), .Y(n_393) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_313), .A2(n_335), .B1(n_344), .B2(n_346), .Y(n_343) );
OAI322xp33_ASAP7_75t_L g491 ( .A1(n_313), .A2(n_412), .A3(n_492), .B1(n_493), .B2(n_494), .C1(n_495), .C2(n_498), .Y(n_491) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g513 ( .A(n_314), .B(n_496), .Y(n_513) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_315), .Y(n_332) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_315), .Y(n_372) );
BUFx3_ASAP7_75t_L g396 ( .A(n_315), .Y(n_396) );
INVx1_ASAP7_75t_L g422 ( .A(n_315), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_315), .Y(n_426) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g380 ( .A(n_319), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g431 ( .A(n_320), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_320), .B(n_388), .Y(n_482) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2x1_ASAP7_75t_L g341 ( .A(n_321), .B(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g345 ( .A(n_321), .Y(n_345) );
AND2x2_ASAP7_75t_L g387 ( .A(n_321), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g408 ( .A(n_321), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_322), .B(n_435), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_330), .B(n_334), .C(n_343), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI31xp33_ASAP7_75t_L g485 ( .A1(n_325), .A2(n_486), .A3(n_488), .B(n_489), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
AND2x4_ASAP7_75t_L g438 ( .A(n_326), .B(n_347), .Y(n_438) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_327), .Y(n_370) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_328), .B(n_348), .Y(n_454) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g494 ( .A(n_337), .Y(n_494) );
AND2x2_ASAP7_75t_L g354 ( .A(n_338), .B(n_345), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_339), .A2(n_424), .B1(n_427), .B2(n_429), .Y(n_423) );
OR2x6_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_SL g481 ( .A(n_342), .Y(n_481) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g451 ( .A(n_347), .B(n_396), .Y(n_451) );
INVx2_ASAP7_75t_L g497 ( .A(n_347), .Y(n_497) );
AND2x4_ASAP7_75t_L g505 ( .A(n_347), .B(n_426), .Y(n_505) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_367), .C(n_397), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_363), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_354), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x4_ASAP7_75t_L g418 ( .A(n_356), .B(n_373), .Y(n_418) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_359), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AND2x2_ASAP7_75t_L g449 ( .A(n_361), .B(n_428), .Y(n_449) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_362), .Y(n_369) );
INVx1_ASAP7_75t_L g487 ( .A(n_362), .Y(n_487) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g516 ( .A(n_365), .Y(n_516) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_366), .Y(n_401) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_373), .B(n_376), .C(n_389), .Y(n_367) );
NOR3x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .C(n_371), .Y(n_368) );
NAND2x1_ASAP7_75t_L g437 ( .A(n_371), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2x1p5_ASAP7_75t_SL g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B1(n_382), .B2(n_385), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g470 ( .A(n_381), .Y(n_470) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g465 ( .A(n_384), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g519 ( .A(n_387), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_394), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g473 ( .A(n_394), .Y(n_473) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g400 ( .A(n_396), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_396), .B(n_454), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B(n_402), .Y(n_397) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_400), .B(n_487), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_410), .B2(n_412), .Y(n_402) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g455 ( .A(n_405), .Y(n_455) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g430 ( .A(n_406), .B(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
INVx1_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_471), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_432), .C(n_445), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_423), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g478 ( .A(n_421), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_430), .B(n_458), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B1(n_439), .B2(n_443), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g488 ( .A(n_438), .Y(n_488) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI21xp33_ASAP7_75t_L g460 ( .A1(n_440), .A2(n_461), .B(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_456), .B1(n_460), .B2(n_468), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_450), .Y(n_446) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_455), .Y(n_450) );
INVx1_ASAP7_75t_L g515 ( .A(n_451), .Y(n_515) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g504 ( .A(n_454), .Y(n_504) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx2_ASAP7_75t_L g496 ( .A(n_466), .Y(n_496) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_490), .Y(n_471) );
AOI211xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_476), .C(n_485), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_480), .C(n_483), .Y(n_476) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_499), .C(n_514), .Y(n_490) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B1(n_506), .B2(n_508), .C(n_509), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_509) );
OAI21xp33_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g886 ( .A(n_524), .Y(n_886) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_750), .Y(n_524) );
NOR2x1_ASAP7_75t_L g525 ( .A(n_526), .B(n_689), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g526 ( .A(n_527), .B(n_640), .C(n_659), .D(n_670), .Y(n_526) );
O2A1O1Ixp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_575), .B(n_582), .C(n_613), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_553), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_529), .B(n_705), .C(n_706), .Y(n_704) );
AND2x2_ASAP7_75t_L g786 ( .A(n_529), .B(n_668), .Y(n_786) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_541), .Y(n_529) );
AND2x2_ASAP7_75t_L g630 ( .A(n_530), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_530), .B(n_649), .Y(n_648) );
INVx3_ASAP7_75t_L g665 ( .A(n_530), .Y(n_665) );
AND2x2_ASAP7_75t_L g710 ( .A(n_530), .B(n_555), .Y(n_710) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g579 ( .A(n_531), .Y(n_579) );
AND2x4_ASAP7_75t_L g658 ( .A(n_531), .B(n_649), .Y(n_658) );
AO31x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .A3(n_538), .B(n_539), .Y(n_531) );
AO31x2_ASAP7_75t_L g607 ( .A1(n_532), .A2(n_550), .A3(n_608), .B(n_611), .Y(n_607) );
AO31x2_ASAP7_75t_L g567 ( .A1(n_538), .A2(n_568), .A3(n_571), .B(n_573), .Y(n_567) );
AND2x2_ASAP7_75t_L g580 ( .A(n_541), .B(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g633 ( .A(n_541), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_541), .Y(n_656) );
INVx1_ASAP7_75t_L g667 ( .A(n_541), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_541), .B(n_565), .Y(n_676) );
INVx2_ASAP7_75t_L g683 ( .A(n_541), .Y(n_683) );
INVx4_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g628 ( .A(n_542), .B(n_555), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_542), .B(n_635), .Y(n_701) );
AND2x2_ASAP7_75t_L g709 ( .A(n_542), .B(n_567), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_542), .B(n_756), .Y(n_755) );
BUFx2_ASAP7_75t_L g762 ( .A(n_542), .Y(n_762) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g778 ( .A(n_554), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_565), .Y(n_554) );
INVx1_ASAP7_75t_L g581 ( .A(n_555), .Y(n_581) );
INVx1_ASAP7_75t_L g635 ( .A(n_555), .Y(n_635) );
INVx2_ASAP7_75t_L g669 ( .A(n_555), .Y(n_669) );
OR2x2_ASAP7_75t_L g673 ( .A(n_555), .B(n_567), .Y(n_673) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_555), .Y(n_722) );
AO31x2_ASAP7_75t_L g585 ( .A1(n_562), .A2(n_571), .A3(n_586), .B(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g695 ( .A(n_566), .B(n_579), .Y(n_695) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_567), .Y(n_631) );
INVx2_ASAP7_75t_L g649 ( .A(n_567), .Y(n_649) );
AND2x4_ASAP7_75t_L g668 ( .A(n_567), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g756 ( .A(n_567), .Y(n_756) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g604 ( .A(n_572), .Y(n_604) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g674 ( .A(n_578), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_578), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g737 ( .A(n_579), .Y(n_737) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_593), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_584), .B(n_594), .Y(n_687) );
INVx1_ASAP7_75t_L g785 ( .A(n_584), .Y(n_785) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g625 ( .A(n_585), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g639 ( .A(n_585), .B(n_618), .Y(n_639) );
AND2x4_ASAP7_75t_L g662 ( .A(n_585), .B(n_606), .Y(n_662) );
INVx2_ASAP7_75t_L g679 ( .A(n_585), .Y(n_679) );
AND2x2_ASAP7_75t_L g705 ( .A(n_585), .B(n_607), .Y(n_705) );
INVx1_ASAP7_75t_L g770 ( .A(n_585), .Y(n_770) );
AND2x2_ASAP7_75t_L g730 ( .A(n_593), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_606), .Y(n_593) );
AND2x2_ASAP7_75t_L g696 ( .A(n_594), .B(n_653), .Y(n_696) );
AND2x4_ASAP7_75t_L g712 ( .A(n_594), .B(n_679), .Y(n_712) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g706 ( .A(n_595), .Y(n_706) );
OAI21x1_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_605), .Y(n_595) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_596), .A2(n_597), .B(n_605), .Y(n_627) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_604), .Y(n_597) );
INVx2_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
INVx3_ASAP7_75t_L g644 ( .A(n_606), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_606), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_606), .B(n_773), .Y(n_772) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g678 ( .A(n_607), .B(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g802 ( .A(n_607), .Y(n_802) );
OAI33xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_628), .A3(n_629), .B1(n_630), .B2(n_632), .B3(n_636), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g736 ( .A(n_617), .B(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g645 ( .A(n_618), .B(n_627), .Y(n_645) );
INVx2_ASAP7_75t_L g653 ( .A(n_618), .Y(n_653) );
INVx1_ASAP7_75t_L g661 ( .A(n_618), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_625), .A2(n_681), .B1(n_684), .B2(n_688), .Y(n_680) );
OR2x2_ASAP7_75t_L g820 ( .A(n_625), .B(n_638), .Y(n_820) );
AND2x4_ASAP7_75t_L g724 ( .A(n_626), .B(n_686), .Y(n_724) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_627), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_628), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g688 ( .A(n_628), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_628), .B(n_664), .Y(n_766) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g739 ( .A(n_630), .Y(n_739) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g797 ( .A(n_633), .B(n_665), .Y(n_797) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_633), .B(n_664), .Y(n_815) );
AND2x2_ASAP7_75t_L g839 ( .A(n_633), .B(n_658), .Y(n_839) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g829 ( .A(n_637), .B(n_706), .Y(n_829) );
NOR2x1p5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g763 ( .A(n_638), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g731 ( .A(n_639), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_646), .B1(n_650), .B2(n_654), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
AND2x2_ASAP7_75t_L g738 ( .A(n_643), .B(n_706), .Y(n_738) );
AND2x2_ASAP7_75t_L g775 ( .A(n_643), .B(n_724), .Y(n_775) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g650 ( .A(n_644), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_644), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g816 ( .A(n_644), .B(n_645), .Y(n_816) );
AND2x2_ASAP7_75t_L g677 ( .A(n_645), .B(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g796 ( .A(n_645), .B(n_662), .Y(n_796) );
AND2x2_ASAP7_75t_L g840 ( .A(n_645), .B(n_705), .Y(n_840) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g774 ( .A1(n_650), .A2(n_775), .B1(n_776), .B2(n_779), .C1(n_781), .C2(n_782), .Y(n_774) );
AND2x2_ASAP7_75t_L g697 ( .A(n_651), .B(n_665), .Y(n_697) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g728 ( .A(n_652), .Y(n_728) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_652), .Y(n_773) );
INVx2_ASAP7_75t_L g686 ( .A(n_653), .Y(n_686) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g743 ( .A(n_656), .Y(n_743) );
INVx2_ASAP7_75t_L g749 ( .A(n_657), .Y(n_749) );
INVx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g733 ( .A(n_658), .B(n_722), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x4_ASAP7_75t_L g764 ( .A(n_661), .B(n_712), .Y(n_764) );
INVx2_ASAP7_75t_L g811 ( .A(n_661), .Y(n_811) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g754 ( .A(n_665), .B(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_L g788 ( .A(n_665), .B(n_673), .Y(n_788) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g693 ( .A(n_667), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_668), .B(n_758), .Y(n_757) );
AND2x4_ASAP7_75t_L g800 ( .A(n_668), .B(n_716), .Y(n_800) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B(n_677), .C(n_680), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
OR2x2_ASAP7_75t_L g681 ( .A(n_673), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g717 ( .A(n_673), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_674), .B(n_709), .Y(n_813) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g789 ( .A(n_676), .B(n_758), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_678), .B(n_728), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_678), .A2(n_694), .B1(n_736), .B2(n_738), .Y(n_735) );
AND2x2_ASAP7_75t_L g741 ( .A(n_678), .B(n_706), .Y(n_741) );
AND2x2_ASAP7_75t_L g810 ( .A(n_678), .B(n_811), .Y(n_810) );
O2A1O1Ixp33_ASAP7_75t_L g803 ( .A1(n_681), .A2(n_783), .B(n_804), .C(n_807), .Y(n_803) );
INVx2_ASAP7_75t_L g716 ( .A(n_683), .Y(n_716) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g794 ( .A(n_686), .Y(n_794) );
INVx1_ASAP7_75t_L g719 ( .A(n_687), .Y(n_719) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_688), .A2(n_735), .B1(n_739), .B2(n_740), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_702), .C(n_725), .Y(n_689) );
AO22x1_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_695), .Y(n_828) );
OR2x2_ASAP7_75t_L g835 ( .A(n_695), .B(n_716), .Y(n_835) );
AND2x2_ASAP7_75t_L g747 ( .A(n_696), .B(n_705), .Y(n_747) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g823 ( .A(n_701), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .C(n_713), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g745 ( .A(n_705), .Y(n_745) );
AND2x4_ASAP7_75t_SL g781 ( .A(n_705), .B(n_724), .Y(n_781) );
INVx1_ASAP7_75t_SL g792 ( .A(n_705), .Y(n_792) );
OR2x2_ASAP7_75t_L g744 ( .A(n_706), .B(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
AND2x4_ASAP7_75t_L g721 ( .A(n_709), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g779 ( .A(n_710), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g801 ( .A(n_712), .B(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g826 ( .A(n_712), .B(n_806), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .B1(n_720), .B2(n_723), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
AND2x4_ASAP7_75t_L g761 ( .A(n_717), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g783 ( .A(n_717), .Y(n_783) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g838 ( .A(n_721), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_734), .C(n_742), .Y(n_725) );
AOI21xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g807 ( .A(n_728), .Y(n_807) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI222xp33_ASAP7_75t_L g830 ( .A1(n_733), .A2(n_831), .B1(n_834), .B2(n_836), .C1(n_838), .C2(n_840), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_736), .B(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g759 ( .A(n_737), .Y(n_759) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B(n_746), .C(n_748), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2x1_ASAP7_75t_L g750 ( .A(n_751), .B(n_808), .Y(n_750) );
NAND4xp25_ASAP7_75t_L g751 ( .A(n_752), .B(n_774), .C(n_784), .D(n_795), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_763), .B1(n_765), .B2(n_767), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .C(n_760), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_754), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g780 ( .A(n_756), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_758), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x4_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g805 ( .A(n_770), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g819 ( .A(n_771), .Y(n_819) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_772), .Y(n_837) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_L g832 ( .A(n_781), .Y(n_832) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B(n_787), .C(n_793), .Y(n_784) );
AOI21xp33_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_789), .B(n_790), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_788), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B1(n_798), .B2(n_801), .C(n_803), .Y(n_795) );
INVx1_ASAP7_75t_L g833 ( .A(n_796), .Y(n_833) );
AOI31xp33_ASAP7_75t_L g817 ( .A1(n_799), .A2(n_818), .A3(n_819), .B(n_820), .Y(n_817) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g806 ( .A(n_802), .Y(n_806) );
INVxp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_821), .C(n_830), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B1(n_814), .B2(n_816), .C(n_817), .Y(n_809) );
INVx2_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_SL g818 ( .A(n_816), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_824), .B1(n_827), .B2(n_829), .Y(n_821) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_841), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g849 ( .A(n_842), .Y(n_849) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NOR2xp33_ASAP7_75t_SL g855 ( .A(n_856), .B(n_859), .Y(n_855) );
INVx4_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AND2x6_ASAP7_75t_SL g864 ( .A(n_858), .B(n_865), .Y(n_864) );
OAI21xp33_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_867), .B(n_880), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
INVx5_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_873), .B1(n_874), .B2(n_879), .Y(n_867) );
XNOR2x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .Y(n_868) );
XOR2x2_ASAP7_75t_L g879 ( .A(n_869), .B(n_872), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_884), .Y(n_880) );
CKINVDCx11_ASAP7_75t_R g882 ( .A(n_883), .Y(n_882) );
endmodule