module fake_jpeg_4322_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_288;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_218;
wire n_63;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_28),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_16),
.B1(n_32),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_16),
.B1(n_26),
.B2(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_88),
.B1(n_58),
.B2(n_51),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_29),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_38),
.B1(n_39),
.B2(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_25),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_33),
.B1(n_23),
.B2(n_39),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_96),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_99),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_49),
.B(n_64),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_84),
.B(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_69),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_102),
.B(n_72),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_116),
.B1(n_86),
.B2(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_112),
.Y(n_123)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_114),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_23),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_66),
.B1(n_48),
.B2(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_56),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_88),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_87),
.B(n_91),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_119),
.B1(n_117),
.B2(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_126),
.B1(n_130),
.B2(n_133),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_86),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_132),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_116),
.B(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_140),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_78),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_52),
.C(n_90),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_101),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_92),
.B1(n_58),
.B2(n_60),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_157)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_112),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_155),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_99),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_169),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_171),
.B1(n_122),
.B2(n_134),
.Y(n_179)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_106),
.B1(n_108),
.B2(n_105),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_170),
.C(n_142),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_190),
.C(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_160),
.B1(n_93),
.B2(n_94),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_131),
.B(n_132),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_195),
.B(n_181),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_158),
.A2(n_138),
.B1(n_126),
.B2(n_144),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_188),
.B1(n_166),
.B2(n_171),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_138),
.B1(n_144),
.B2(n_140),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_142),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_128),
.C(n_137),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_120),
.C(n_133),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_194),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_120),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_134),
.B(n_145),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_73),
.B1(n_85),
.B2(n_94),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_196),
.A2(n_147),
.B1(n_156),
.B2(n_155),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_210),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_216),
.B1(n_189),
.B2(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_184),
.B1(n_186),
.B2(n_195),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_174),
.B1(n_187),
.B2(n_178),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_154),
.C(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_211),
.Y(n_234)
);

OAI221xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_165),
.B1(n_159),
.B2(n_150),
.C(n_169),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_205),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_157),
.B(n_74),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_208),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_146),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_28),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_200),
.B(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_217),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_93),
.B1(n_21),
.B2(n_25),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_173),
.C(n_192),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_230),
.C(n_29),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_236),
.B1(n_202),
.B2(n_22),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_212),
.C(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_209),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_238),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_21),
.B1(n_31),
.B2(n_167),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_70),
.B1(n_35),
.B2(n_30),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_35),
.B1(n_63),
.B2(n_22),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_214),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_248),
.B(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_229),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_247),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_20),
.B1(n_17),
.B2(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

XOR2x1_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_29),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_254),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_29),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_255),
.B1(n_22),
.B2(n_20),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_12),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_223),
.A2(n_30),
.B1(n_35),
.B2(n_63),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_227),
.B(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

AO221x1_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_237),
.B1(n_224),
.B2(n_17),
.C(n_22),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_20),
.B1(n_17),
.B2(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_226),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_230),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_268),
.B1(n_260),
.B2(n_3),
.Y(n_279)
);

AOI221xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_241),
.C(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_251),
.C(n_244),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_272),
.C(n_277),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_9),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_250),
.C(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_261),
.C(n_263),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_1),
.C(n_20),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_282),
.B(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_8),
.Y(n_282)
);

AOI211xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_8),
.B(n_2),
.C(n_4),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_1),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_273),
.B(n_6),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_14),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_276),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_291),
.B(n_294),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_293),
.B(n_286),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_281),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_10),
.C(n_12),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_5),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

AOI321xp33_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_298),
.A3(n_13),
.B1(n_14),
.B2(n_289),
.C(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_295),
.B(n_299),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_13),
.Y(n_303)
);


endmodule