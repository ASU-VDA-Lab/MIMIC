module fake_jpeg_5315_n_117 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_117);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_117;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_42),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_15),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_12),
.B1(n_19),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_10),
.B1(n_19),
.B2(n_14),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_12),
.B1(n_32),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_57),
.B1(n_24),
.B2(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_58),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_43),
.B1(n_24),
.B2(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_44),
.B(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_18),
.C(n_22),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_12),
.B1(n_25),
.B2(n_11),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_13),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_33),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_69),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_43),
.B(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_72),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_24),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_80),
.B1(n_73),
.B2(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_72),
.B(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_78),
.B(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_66),
.B1(n_64),
.B2(n_68),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_77),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_98),
.C(n_99),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_82),
.A3(n_77),
.B1(n_76),
.B2(n_75),
.Y(n_96)
);

OAI21x1_ASAP7_75t_R g97 ( 
.A1(n_86),
.A2(n_34),
.B(n_61),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_73),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_87),
.C(n_89),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_93),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_88),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_92),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_102),
.C(n_100),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_41),
.B1(n_30),
.B2(n_34),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_41),
.B1(n_34),
.B2(n_33),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_29),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_13),
.C(n_23),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_21),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_21),
.C(n_20),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_111),
.C(n_23),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_5),
.C(n_6),
.Y(n_115)
);

XNOR2x2_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_8),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_17),
.Y(n_117)
);


endmodule