module fake_aes_4519_n_545 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_545);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_545;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_41), .Y(n_78) );
INVx3_ASAP7_75t_L g79 ( .A(n_75), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_58), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_44), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_13), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_55), .Y(n_83) );
BUFx5_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_9), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_52), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_24), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_29), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_50), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_47), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_54), .Y(n_91) );
INVx3_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_32), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_49), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_43), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_6), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_59), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_42), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_15), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_13), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_33), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_5), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_27), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_1), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_56), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_66), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_36), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_20), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_69), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_38), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_15), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_100), .B(n_0), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_85), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_101), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_97), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_79), .B(n_0), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_79), .B(n_1), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_79), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_85), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_116), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_92), .B(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_97), .Y(n_128) );
BUFx8_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_116), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_104), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_82), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_102), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_92), .B(n_6), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_92), .B(n_7), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_106), .B(n_80), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_120), .Y(n_139) );
OR2x6_ASAP7_75t_L g140 ( .A(n_126), .B(n_82), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_123), .B(n_81), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_123), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_129), .B(n_83), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_124), .B(n_81), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_119), .B(n_83), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_128), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_121), .B(n_90), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_129), .B(n_90), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_133), .B(n_110), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_117), .B(n_114), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_137), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_117), .B(n_115), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_125), .B(n_87), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_134), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_138), .B(n_105), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_142), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_156), .A2(n_127), .B1(n_125), .B2(n_132), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
CKINVDCx11_ASAP7_75t_R g168 ( .A(n_140), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_145), .A2(n_89), .B(n_86), .C(n_115), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_159), .B(n_160), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_159), .B(n_114), .Y(n_171) );
INVxp67_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_160), .B(n_87), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_162), .B(n_95), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_162), .B(n_130), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_156), .A2(n_89), .B1(n_86), .B2(n_111), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_148), .B(n_130), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_154), .B(n_118), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_153), .B(n_88), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
INVxp67_ASAP7_75t_L g187 ( .A(n_154), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_156), .A2(n_98), .B1(n_113), .B2(n_118), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_143), .A2(n_88), .B(n_111), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_156), .A2(n_96), .B1(n_108), .B2(n_93), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_157), .B(n_107), .Y(n_192) );
AND2x6_ASAP7_75t_SL g193 ( .A(n_140), .B(n_94), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_147), .B(n_109), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_144), .B(n_84), .Y(n_196) );
BUFx8_ASAP7_75t_SL g197 ( .A(n_175), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_170), .A2(n_141), .B1(n_147), .B2(n_144), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_167), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_170), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_176), .Y(n_204) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_195), .B(n_141), .Y(n_205) );
OAI21x1_ASAP7_75t_SL g206 ( .A1(n_190), .A2(n_153), .B(n_150), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_170), .B(n_156), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_171), .B(n_156), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_183), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_171), .B(n_173), .Y(n_214) );
OR2x6_ASAP7_75t_L g215 ( .A(n_195), .B(n_141), .Y(n_215) );
INVxp67_ASAP7_75t_L g216 ( .A(n_184), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_190), .A2(n_185), .B(n_194), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_173), .B(n_156), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_167), .B(n_153), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_178), .B(n_153), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_187), .B(n_151), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_194), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_178), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_172), .B(n_147), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_164), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_172), .A2(n_147), .B1(n_141), .B2(n_140), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_214), .A2(n_169), .B(n_161), .C(n_174), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_218), .A2(n_189), .B(n_179), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_212), .A2(n_187), .B(n_174), .C(n_182), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
AOI21x1_ASAP7_75t_L g234 ( .A1(n_206), .A2(n_186), .B(n_189), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_218), .A2(n_189), .B(n_179), .Y(n_235) );
AOI221xp5_ASAP7_75t_L g236 ( .A1(n_216), .A2(n_182), .B1(n_165), .B2(n_152), .C(n_192), .Y(n_236) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_207), .A2(n_80), .A3(n_91), .B(n_112), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_211), .A2(n_196), .B(n_179), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_224), .A2(n_186), .B(n_164), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_206), .A2(n_180), .B(n_181), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_202), .B(n_195), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_207), .A2(n_180), .B(n_181), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_202), .B(n_188), .Y(n_244) );
OAI222xp33_ASAP7_75t_L g245 ( .A1(n_201), .A2(n_188), .B1(n_140), .B2(n_195), .C1(n_177), .C2(n_191), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_204), .A2(n_91), .B(n_112), .Y(n_247) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_204), .A2(n_180), .B(n_139), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_202), .B(n_178), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_202), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_207), .A2(n_181), .B(n_139), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_208), .A2(n_181), .B(n_149), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_213), .A2(n_149), .B(n_146), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_213), .A2(n_84), .B(n_109), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_230), .A2(n_224), .B(n_222), .C(n_219), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_245), .B(n_197), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_256), .B(n_205), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_256), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_251), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_248), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_232), .B(n_210), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_249), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_251), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_230), .B(n_223), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_236), .A2(n_168), .B1(n_205), .B2(n_140), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_248), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_244), .A2(n_205), .B1(n_199), .B2(n_203), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_229), .B1(n_215), .B2(n_198), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_215), .B1(n_209), .B2(n_226), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
OAI33xp33_ASAP7_75t_L g274 ( .A1(n_246), .A2(n_223), .A3(n_203), .B1(n_221), .B2(n_193), .B3(n_217), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_241), .B(n_215), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_215), .B1(n_220), .B2(n_225), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_250), .A2(n_215), .B1(n_158), .B2(n_200), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_250), .A2(n_158), .B1(n_225), .B2(n_210), .Y(n_278) );
OAI221xp5_ASAP7_75t_L g279 ( .A1(n_239), .A2(n_163), .B1(n_220), .B2(n_193), .C(n_103), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_259), .B(n_247), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_262), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_269), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_269), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_269), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_267), .B(n_237), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_270), .B(n_237), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_259), .B(n_247), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_260), .B(n_247), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_273), .B(n_233), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_264), .B(n_237), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_270), .B(n_237), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_271), .B(n_237), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_273), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_268), .Y(n_298) );
OAI221xp5_ASAP7_75t_L g299 ( .A1(n_258), .A2(n_220), .B1(n_163), .B2(n_238), .C(n_234), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_257), .B(n_248), .Y(n_301) );
BUFx2_ASAP7_75t_SL g302 ( .A(n_284), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_286), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_285), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_294), .B(n_266), .Y(n_309) );
INVx5_ASAP7_75t_SL g310 ( .A(n_293), .Y(n_310) );
AOI211xp5_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_279), .B(n_276), .C(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_292), .Y(n_313) );
NAND2xp33_ASAP7_75t_SL g314 ( .A(n_297), .B(n_273), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_294), .B(n_266), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_296), .A2(n_279), .B1(n_272), .B2(n_275), .C(n_261), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_283), .B(n_240), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_296), .B(n_240), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_291), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_288), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_288), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
AND2x4_ASAP7_75t_SL g327 ( .A(n_293), .B(n_273), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_280), .B(n_268), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_280), .B(n_231), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_290), .B(n_231), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_309), .B(n_295), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_323), .B(n_295), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_305), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_313), .B(n_290), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_309), .B(n_291), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_322), .B(n_289), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_322), .B(n_289), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_315), .B(n_301), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_324), .A2(n_99), .B1(n_163), .B2(n_275), .C(n_299), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_323), .B(n_301), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_300), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_311), .A2(n_263), .B(n_255), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_323), .B(n_300), .Y(n_350) );
AOI31xp33_ASAP7_75t_L g351 ( .A1(n_314), .A2(n_297), .A3(n_293), .B(n_265), .Y(n_351) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_320), .B(n_103), .C(n_277), .D(n_278), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_328), .B(n_300), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
AOI21x1_ASAP7_75t_L g355 ( .A1(n_321), .A2(n_255), .B(n_235), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_307), .B(n_293), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_328), .B(n_298), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_330), .B(n_298), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_325), .B(n_298), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_308), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_312), .B(n_298), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_327), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_329), .B(n_298), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_329), .B(n_235), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_330), .B(n_84), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_321), .B(n_84), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_306), .B(n_163), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_317), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_312), .B(n_316), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_316), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_318), .B(n_84), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_317), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_361), .B(n_307), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_357), .B(n_304), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_366), .B(n_319), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_346), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_339), .B(n_319), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_352), .B(n_338), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_334), .B(n_318), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_366), .B(n_317), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_352), .B(n_302), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_346), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_334), .B(n_302), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_363), .A2(n_327), .B1(n_310), .B2(n_84), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_310), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_335), .B(n_310), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_337), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_367), .Y(n_391) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_331), .B(n_327), .Y(n_392) );
AOI322xp5_ASAP7_75t_L g393 ( .A1(n_342), .A2(n_99), .A3(n_8), .B1(n_9), .B2(n_10), .C1(n_7), .C2(n_12), .Y(n_393) );
NOR2xp67_ASAP7_75t_SL g394 ( .A(n_354), .B(n_233), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_357), .B(n_310), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_337), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_342), .B(n_310), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_367), .B(n_84), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_332), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_333), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_333), .Y(n_402) );
OAI21xp33_ASAP7_75t_L g403 ( .A1(n_351), .A2(n_99), .B(n_254), .Y(n_403) );
OR2x6_ASAP7_75t_L g404 ( .A(n_354), .B(n_252), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_347), .B(n_99), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_344), .B(n_8), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_344), .B(n_10), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_337), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_336), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_354), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_336), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_340), .B(n_11), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_353), .B(n_99), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_340), .B(n_11), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_341), .B(n_12), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_348), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_353), .B(n_14), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_356), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_348), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_345), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_345), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_348), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_372), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_368), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_356), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_376), .B(n_341), .Y(n_427) );
AOI32xp33_ASAP7_75t_L g428 ( .A1(n_380), .A2(n_335), .A3(n_373), .B1(n_365), .B2(n_358), .Y(n_428) );
AOI32xp33_ASAP7_75t_L g429 ( .A1(n_380), .A2(n_335), .A3(n_373), .B1(n_365), .B2(n_358), .Y(n_429) );
NOR3xp33_ASAP7_75t_L g430 ( .A(n_412), .B(n_351), .C(n_349), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_414), .A2(n_335), .B1(n_349), .B2(n_365), .C(n_368), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_418), .B(n_364), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_392), .A2(n_359), .B1(n_365), .B2(n_364), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_405), .B(n_371), .Y(n_434) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_403), .B(n_359), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_415), .A2(n_343), .B1(n_362), .B2(n_371), .C(n_369), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_426), .B(n_350), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_393), .B(n_369), .C(n_350), .Y(n_438) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_383), .A2(n_355), .B(n_360), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_406), .A2(n_360), .B(n_374), .C(n_370), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_413), .B(n_360), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_378), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_381), .B(n_374), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_390), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_384), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_375), .B(n_374), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_399), .A2(n_370), .B(n_14), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_392), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_426), .B(n_370), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_395), .B(n_355), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_396), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_383), .A2(n_252), .B(n_253), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_379), .B(n_253), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g454 ( .A1(n_386), .A2(n_254), .B(n_233), .C(n_243), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_391), .B(n_233), .Y(n_455) );
AOI321xp33_ASAP7_75t_L g456 ( .A1(n_391), .A2(n_217), .A3(n_228), .B1(n_22), .B2(n_23), .C(n_25), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_417), .A2(n_243), .B(n_217), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_388), .B(n_17), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_390), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_404), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_396), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_401), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_387), .Y(n_465) );
AOI221x1_ASAP7_75t_L g466 ( .A1(n_425), .A2(n_225), .B1(n_210), .B2(n_200), .C(n_228), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_402), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_388), .B(n_21), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_410), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_409), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_411), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_442), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_445), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_440), .A2(n_407), .B(n_410), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g475 ( .A1(n_430), .A2(n_385), .B1(n_397), .B2(n_377), .C(n_421), .Y(n_475) );
AOI21xp5_ASAP7_75t_SL g476 ( .A1(n_448), .A2(n_404), .B(n_385), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_460), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_461), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_432), .B(n_404), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_469), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_464), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_465), .Y(n_482) );
AOI222xp33_ASAP7_75t_L g483 ( .A1(n_431), .A2(n_420), .B1(n_424), .B2(n_423), .C1(n_382), .C2(n_419), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_435), .A2(n_422), .B(n_419), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_467), .Y(n_485) );
OAI311xp33_ASAP7_75t_L g486 ( .A1(n_439), .A2(n_394), .A3(n_416), .B1(n_408), .C1(n_422), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_470), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_446), .B(n_416), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_471), .Y(n_489) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_433), .B(n_408), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_446), .B(n_389), .Y(n_493) );
XNOR2x1_ASAP7_75t_L g494 ( .A(n_427), .B(n_389), .Y(n_494) );
XNOR2x1_ASAP7_75t_L g495 ( .A(n_437), .B(n_26), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_451), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_444), .B(n_28), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_449), .Y(n_498) );
OAI322xp33_ASAP7_75t_L g499 ( .A1(n_444), .A2(n_225), .A3(n_210), .B1(n_200), .B2(n_35), .C1(n_37), .C2(n_39), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
AOI22x1_ASAP7_75t_L g502 ( .A1(n_483), .A2(n_448), .B1(n_456), .B2(n_462), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_501), .B(n_459), .Y(n_503) );
OAI21xp33_ASAP7_75t_SL g504 ( .A1(n_494), .A2(n_428), .B(n_429), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_482), .B(n_462), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_491), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_472), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_500), .B(n_430), .Y(n_508) );
XOR2x2_ASAP7_75t_L g509 ( .A(n_495), .B(n_438), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_475), .A2(n_440), .B1(n_447), .B2(n_450), .C(n_463), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_473), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_474), .A2(n_486), .B1(n_500), .B2(n_476), .C(n_490), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_477), .A2(n_434), .B1(n_436), .B2(n_441), .C(n_457), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_478), .A2(n_452), .B1(n_458), .B2(n_468), .C(n_454), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_481), .Y(n_515) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_480), .A2(n_453), .B(n_466), .C(n_455), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_492), .B(n_30), .Y(n_517) );
OAI21xp33_ASAP7_75t_L g518 ( .A1(n_488), .A2(n_225), .B(n_210), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_485), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_508), .A2(n_496), .B1(n_487), .B2(n_489), .C1(n_493), .C2(n_498), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_504), .A2(n_510), .B1(n_512), .B2(n_513), .C(n_516), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_506), .Y(n_522) );
NOR4xp75_ASAP7_75t_L g523 ( .A(n_502), .B(n_499), .C(n_495), .D(n_479), .Y(n_523) );
AOI211xp5_ASAP7_75t_SL g524 ( .A1(n_514), .A2(n_497), .B(n_484), .C(n_40), .Y(n_524) );
OAI222xp33_ASAP7_75t_L g525 ( .A1(n_505), .A2(n_484), .B1(n_497), .B2(n_45), .C1(n_46), .C2(n_48), .Y(n_525) );
NOR2xp33_ASAP7_75t_SL g526 ( .A(n_505), .B(n_200), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_503), .B(n_31), .Y(n_527) );
OAI211xp5_ASAP7_75t_L g528 ( .A1(n_509), .A2(n_34), .B(n_57), .C(n_60), .Y(n_528) );
NAND3xp33_ASAP7_75t_SL g529 ( .A(n_517), .B(n_61), .C(n_62), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_528), .B(n_519), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_521), .B(n_515), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_522), .A2(n_511), .B1(n_507), .B2(n_518), .C(n_67), .Y(n_532) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_525), .B(n_63), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_527), .Y(n_534) );
NOR3xp33_ASAP7_75t_L g535 ( .A(n_531), .B(n_529), .C(n_523), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_534), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_530), .Y(n_537) );
AOI22x1_ASAP7_75t_L g538 ( .A1(n_537), .A2(n_520), .B1(n_524), .B2(n_533), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_536), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_539), .Y(n_540) );
XOR2xp5_ASAP7_75t_L g541 ( .A(n_538), .B(n_535), .Y(n_541) );
OA22x2_ASAP7_75t_L g542 ( .A1(n_541), .A2(n_532), .B1(n_526), .B2(n_68), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_542), .A2(n_540), .B1(n_65), .B2(n_71), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_543), .Y(n_544) );
OAI321xp33_ASAP7_75t_L g545 ( .A1(n_544), .A2(n_64), .A3(n_72), .B1(n_73), .B2(n_76), .C(n_77), .Y(n_545) );
endmodule