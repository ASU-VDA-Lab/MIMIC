module fake_jpeg_16457_n_306 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_47),
.Y(n_93)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_2),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_21),
.C(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_60),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_2),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_66),
.Y(n_81)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_69),
.Y(n_84)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_3),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_20),
.B1(n_29),
.B2(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_88),
.B1(n_103),
.B2(n_109),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_112),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_40),
.A2(n_39),
.B1(n_20),
.B2(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_89),
.B(n_115),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_41),
.B(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_43),
.A2(n_15),
.B1(n_35),
.B2(n_34),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_28),
.C(n_26),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_76),
.C(n_95),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_49),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_38),
.B1(n_28),
.B2(n_26),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_51),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_111),
.B1(n_116),
.B2(n_90),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_48),
.A2(n_25),
.B1(n_24),
.B2(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_46),
.B(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_68),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_45),
.B(n_10),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_10),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_84),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_122),
.B(n_130),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_58),
.B1(n_62),
.B2(n_64),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_149),
.B1(n_105),
.B2(n_145),
.Y(n_166)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_145),
.B(n_150),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_76),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_13),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_132),
.B(n_143),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_134),
.B(n_142),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_82),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_146),
.C(n_140),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_144),
.Y(n_170)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_78),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_102),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_92),
.B1(n_98),
.B2(n_90),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_157),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_102),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_92),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_159),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_74),
.B(n_75),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_123),
.Y(n_167)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g181 ( 
.A(n_163),
.Y(n_181)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_133),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_167),
.B(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_144),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_182),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_141),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_124),
.Y(n_183)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_127),
.A2(n_150),
.B1(n_123),
.B2(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_184),
.B1(n_166),
.B2(n_183),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_129),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_211),
.C(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_138),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_200),
.B(n_207),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_161),
.B1(n_152),
.B2(n_163),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_133),
.B(n_152),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_220),
.B(n_226),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_SL g242 ( 
.A1(n_206),
.A2(n_181),
.B(n_185),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_198),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_178),
.B1(n_180),
.B2(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_169),
.C(n_176),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_215),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_192),
.B(n_173),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_216),
.B(n_218),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_196),
.A2(n_191),
.B1(n_192),
.B2(n_175),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_182),
.B(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_225),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_187),
.B(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_175),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_190),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_197),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_179),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_186),
.C(n_181),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_237),
.B1(n_228),
.B2(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_202),
.B1(n_208),
.B2(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_180),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_185),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_241),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_204),
.B(n_226),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_190),
.B(n_186),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_181),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.C(n_247),
.Y(n_251)
);

AO22x2_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_204),
.B1(n_206),
.B2(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_231),
.B1(n_234),
.B2(n_245),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_211),
.C(n_221),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_257),
.C(n_251),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_229),
.B(n_233),
.Y(n_271)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_209),
.C(n_215),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_236),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_265),
.B1(n_239),
.B2(n_201),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_209),
.B1(n_201),
.B2(n_210),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_278),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_251),
.C(n_254),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_244),
.B(n_235),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_271),
.B(n_272),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_249),
.B(n_260),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_275),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_261),
.B1(n_252),
.B2(n_263),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_234),
.B(n_237),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_230),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.C(n_282),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_267),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_259),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_284),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_286),
.A2(n_276),
.B1(n_269),
.B2(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_241),
.C(n_252),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_230),
.C(n_256),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_276),
.B(n_255),
.C(n_271),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_262),
.B(n_270),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_291),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_287),
.C(n_282),
.Y(n_299)
);

OAI221xp5_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_294),
.B1(n_285),
.B2(n_292),
.C(n_219),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_292),
.C(n_279),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_281),
.C(n_295),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_296),
.B(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_203),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);


endmodule