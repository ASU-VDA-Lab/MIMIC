module fake_jpeg_13373_n_426 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_56),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_31),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_64),
.B(n_66),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_72),
.Y(n_169)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_75),
.Y(n_171)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_12),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_20),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_89),
.B(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_95),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_96),
.B(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_103),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_R g142 ( 
.A(n_99),
.Y(n_142)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_13),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_102),
.B(n_109),
.Y(n_170)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_14),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_106),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_14),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_33),
.B1(n_55),
.B2(n_48),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_176),
.B1(n_32),
.B2(n_65),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_55),
.B1(n_25),
.B2(n_48),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_148),
.B1(n_32),
.B2(n_54),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_33),
.B1(n_48),
.B2(n_25),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_129),
.A2(n_6),
.B1(n_166),
.B2(n_122),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_64),
.B(n_47),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_37),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_140),
.B(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_37),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_50),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_68),
.A2(n_25),
.B1(n_49),
.B2(n_39),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_110),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_50),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_89),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_155),
.B(n_160),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_47),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_59),
.B(n_26),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_163),
.B(n_164),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_26),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_36),
.B1(n_54),
.B2(n_41),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_6),
.B1(n_129),
.B2(n_171),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_99),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_172),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_81),
.B(n_41),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_82),
.B(n_46),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_46),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_101),
.A2(n_107),
.B1(n_106),
.B2(n_36),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_196),
.Y(n_235)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_125),
.A2(n_148),
.B1(n_176),
.B2(n_113),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_179),
.A2(n_187),
.B1(n_200),
.B2(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_193),
.Y(n_233)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_124),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_217),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_3),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_201),
.B(n_232),
.C(n_126),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_208),
.Y(n_257)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_206),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_116),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_116),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_218),
.Y(n_262)
);

BUFx2_ASAP7_75t_SL g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_210),
.Y(n_246)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_211),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_137),
.B(n_16),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_212),
.B(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_170),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_150),
.B(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_117),
.Y(n_216)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_156),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_119),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_133),
.B1(n_151),
.B2(n_121),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_6),
.B1(n_113),
.B2(n_156),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_225),
.A2(n_227),
.B1(n_229),
.B2(n_132),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_169),
.A2(n_171),
.B1(n_145),
.B2(n_123),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_145),
.A2(n_123),
.B1(n_115),
.B2(n_167),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_147),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_234),
.B(n_195),
.Y(n_291)
);

AO22x2_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_131),
.B1(n_138),
.B2(n_121),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_245),
.B1(n_261),
.B2(n_270),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_183),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_242),
.A2(n_252),
.B1(n_265),
.B2(n_237),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_182),
.B(n_167),
.C(n_165),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_258),
.C(n_219),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_187),
.A2(n_188),
.B1(n_207),
.B2(n_197),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_146),
.B1(n_158),
.B2(n_135),
.Y(n_252)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_198),
.A2(n_131),
.A3(n_165),
.B1(n_146),
.B2(n_133),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_267),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_126),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_207),
.A2(n_158),
.B1(n_118),
.B2(n_132),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_197),
.A2(n_118),
.B1(n_132),
.B2(n_153),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_215),
.A2(n_153),
.B1(n_220),
.B2(n_213),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_274),
.B1(n_194),
.B2(n_217),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_213),
.A2(n_220),
.B1(n_228),
.B2(n_212),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_279),
.B(n_285),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_280),
.A2(n_284),
.B(n_304),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_281),
.A2(n_310),
.B1(n_270),
.B2(n_261),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_289),
.B1(n_300),
.B2(n_246),
.Y(n_331)
);

A2O1A1O1Ixp25_ASAP7_75t_L g284 ( 
.A1(n_233),
.A2(n_226),
.B(n_230),
.C(n_181),
.D(n_185),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_192),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_199),
.B1(n_191),
.B2(n_216),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_301),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_218),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_299),
.Y(n_318)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_245),
.A2(n_206),
.B1(n_211),
.B2(n_186),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_221),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_308),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_231),
.C(n_178),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_305),
.C(n_248),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_239),
.A2(n_190),
.B(n_203),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_184),
.C(n_204),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_309),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_205),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_252),
.B1(n_237),
.B2(n_242),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_319),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_282),
.A2(n_241),
.B1(n_251),
.B2(n_266),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_312),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_266),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_241),
.C(n_243),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_235),
.C(n_251),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_330),
.A2(n_332),
.B(n_307),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_331),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_281),
.A2(n_254),
.B(n_276),
.C(n_272),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_277),
.A2(n_244),
.B1(n_271),
.B2(n_276),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_308),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_356),
.C(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_330),
.A2(n_277),
.B1(n_289),
.B2(n_278),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_341),
.B1(n_327),
.B2(n_306),
.Y(n_371)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_332),
.A2(n_300),
.B1(n_283),
.B2(n_280),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_344),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_329),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_SL g346 ( 
.A(n_325),
.B(n_307),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_346),
.A2(n_351),
.B(n_320),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_347),
.A2(n_353),
.B1(n_316),
.B2(n_332),
.Y(n_363)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_350),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_319),
.A2(n_304),
.B(n_334),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_355),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_301),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_268),
.C(n_260),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_336),
.B(n_312),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_338),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_324),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_363),
.A2(n_373),
.B1(n_351),
.B2(n_345),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_366),
.C(n_370),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_314),
.C(n_332),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_311),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_356),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_345),
.A2(n_332),
.B1(n_328),
.B2(n_326),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_371),
.B1(n_343),
.B2(n_348),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_327),
.C(n_329),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_333),
.B1(n_317),
.B2(n_287),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_365),
.C(n_366),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_346),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_381),
.Y(n_390)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_361),
.Y(n_378)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_SL g380 ( 
.A1(n_372),
.A2(n_353),
.B(n_344),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_382),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_346),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_363),
.A2(n_347),
.B(n_343),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_385),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_387),
.Y(n_393)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_354),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_370),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_367),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_391),
.B(n_396),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_374),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_381),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_362),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_395),
.A2(n_368),
.B1(n_384),
.B2(n_382),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_393),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_397),
.A2(n_371),
.B1(n_373),
.B2(n_357),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_400),
.A2(n_404),
.B1(n_392),
.B2(n_393),
.Y(n_408)
);

AO221x1_ASAP7_75t_L g401 ( 
.A1(n_389),
.A2(n_337),
.B1(n_339),
.B2(n_355),
.C(n_340),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_402),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_398),
.A2(n_375),
.B1(n_374),
.B2(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_400),
.Y(n_411)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g414 ( 
.A1(n_407),
.A2(n_404),
.A3(n_399),
.B1(n_333),
.B2(n_317),
.C1(n_402),
.C2(n_264),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_409),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_411),
.A2(n_412),
.B(n_390),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_403),
.B(n_394),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_415),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_390),
.B(n_299),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_416),
.B(n_417),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_296),
.B(n_286),
.Y(n_417)
);

BUFx24_ASAP7_75t_SL g418 ( 
.A(n_413),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_418),
.A2(n_409),
.B(n_407),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_421),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_263),
.C(n_284),
.Y(n_422)
);

AOI322xp5_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_422),
.A3(n_419),
.B1(n_236),
.B2(n_256),
.C1(n_272),
.C2(n_255),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_424),
.A2(n_236),
.B(n_256),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_153),
.Y(n_426)
);


endmodule