module fake_jpeg_1916_n_234 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_234);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g62 ( 
.A(n_30),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_82),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_76),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_60),
.B1(n_71),
.B2(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_60),
.B1(n_61),
.B2(n_71),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_76),
.B1(n_74),
.B2(n_78),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_SL g98 ( 
.A(n_83),
.Y(n_98)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_97),
.B1(n_74),
.B2(n_89),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_70),
.C(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_116),
.B1(n_119),
.B2(n_62),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_99),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_107),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_56),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_68),
.B1(n_74),
.B2(n_66),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_63),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_66),
.B1(n_53),
.B2(n_69),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_112),
.B1(n_72),
.B2(n_73),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_129),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_87),
.A3(n_69),
.B1(n_77),
.B2(n_54),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_53),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_54),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_136),
.B(n_0),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_58),
.Y(n_136)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_97),
.B(n_87),
.C(n_90),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_23),
.B(n_5),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_139),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_87),
.B1(n_90),
.B2(n_58),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_107),
.B1(n_111),
.B2(n_104),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_72),
.B(n_62),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_151),
.B(n_163),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_159),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_112),
.B1(n_73),
.B2(n_50),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_162),
.B1(n_130),
.B2(n_6),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_6),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_128),
.B1(n_121),
.B2(n_141),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_49),
.B1(n_46),
.B2(n_43),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_36),
.C(n_35),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_4),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_133),
.CI(n_130),
.CON(n_163),
.SN(n_163)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_163),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_24),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_22),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_5),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_185),
.C(n_8),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_157),
.B1(n_152),
.B2(n_160),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_7),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_176),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_7),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_183),
.B(n_187),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_184),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_8),
.B(n_9),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_201),
.C(n_185),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_162),
.B(n_159),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_184),
.B(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_177),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_12),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_170),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_10),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_208),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_206),
.Y(n_218)
);

AO22x2_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_186),
.B1(n_177),
.B2(n_167),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_168),
.B(n_12),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_11),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_189),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_196),
.B1(n_194),
.B2(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_200),
.C(n_201),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_13),
.C(n_14),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_202),
.B1(n_200),
.B2(n_206),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_222),
.B1(n_219),
.B2(n_217),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_13),
.B(n_14),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_215),
.C(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_223),
.B(n_220),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_214),
.B(n_16),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_15),
.B(n_17),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_17),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_232),
.A2(n_20),
.B(n_21),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_20),
.Y(n_234)
);


endmodule