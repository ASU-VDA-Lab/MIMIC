module fake_jpeg_2031_n_169 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_27),
.Y(n_28)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_10),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_44),
.Y(n_86)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_48),
.Y(n_59)
);

NOR2xp67_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_2),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_2),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_53),
.Y(n_84)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_29),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_4),
.B(n_55),
.Y(n_78)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_32),
.A2(n_18),
.B1(n_19),
.B2(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_73),
.B1(n_81),
.B2(n_62),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_31),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_28),
.A2(n_4),
.B1(n_50),
.B2(n_57),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_42),
.B1(n_52),
.B2(n_70),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_30),
.A2(n_40),
.B1(n_53),
.B2(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_39),
.B(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_29),
.B(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_34),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_66),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_95),
.B1(n_100),
.B2(n_102),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_63),
.B1(n_65),
.B2(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_62),
.B1(n_79),
.B2(n_60),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_74),
.B(n_68),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_89),
.B(n_108),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_122),
.B(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_110),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_104),
.B1(n_89),
.B2(n_100),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_104),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_128),
.B(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_89),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_114),
.C(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_98),
.B1(n_76),
.B2(n_80),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_124),
.A3(n_134),
.B1(n_128),
.B2(n_121),
.C1(n_120),
.C2(n_135),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_113),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_133),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_128),
.C(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_125),
.B1(n_127),
.B2(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_120),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_139),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_151),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_145),
.B1(n_141),
.B2(n_138),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_147),
.B1(n_141),
.B2(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_153),
.C(n_75),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_120),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_146),
.B1(n_150),
.B2(n_143),
.Y(n_159)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_142),
.B(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_162),
.B(n_159),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_112),
.C(n_103),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_112),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_160),
.A3(n_165),
.B1(n_103),
.B2(n_76),
.C(n_94),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_94),
.Y(n_169)
);


endmodule