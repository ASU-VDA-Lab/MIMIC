module fake_jpeg_32163_n_476 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g152 ( 
.A(n_51),
.Y(n_152)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_19),
.Y(n_109)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_61),
.B(n_80),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_76),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_32),
.B(n_8),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_38),
.B(n_7),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_38),
.B(n_9),
.C(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_92),
.Y(n_151)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_9),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_96),
.Y(n_146)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_19),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_28),
.Y(n_147)
);

NOR4xp25_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_39),
.C(n_46),
.D(n_47),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_25),
.C(n_20),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_90),
.B1(n_50),
.B2(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_105),
.A2(n_150),
.B1(n_25),
.B2(n_30),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_46),
.B1(n_42),
.B2(n_33),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_108),
.A2(n_112),
.B1(n_114),
.B2(n_130),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_21),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_128),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_48),
.B1(n_42),
.B2(n_33),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_51),
.A2(n_42),
.B1(n_48),
.B2(n_36),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_113),
.A2(n_62),
.B1(n_57),
.B2(n_52),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_42),
.B1(n_48),
.B2(n_36),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_20),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_75),
.A2(n_48),
.B1(n_36),
.B2(n_28),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_85),
.B1(n_82),
.B2(n_79),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_134),
.A2(n_55),
.B1(n_25),
.B2(n_31),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_28),
.B1(n_36),
.B2(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_19),
.B1(n_17),
.B2(n_34),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_54),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_92),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_70),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_28),
.B1(n_41),
.B2(n_40),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_109),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_106),
.B(n_30),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_163),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_30),
.B(n_43),
.C(n_41),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_17),
.B(n_34),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_111),
.Y(n_163)
);

OR2x2_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_66),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_164),
.B(n_189),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_172),
.A2(n_135),
.B1(n_34),
.B2(n_127),
.Y(n_228)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_175),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_29),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_29),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_181),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_185),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_140),
.B(n_29),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_179),
.B(n_195),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_187),
.B1(n_193),
.B2(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_21),
.Y(n_181)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_21),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_192),
.Y(n_209)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_70),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_190),
.Y(n_231)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_67),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_102),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_146),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_199),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_120),
.B1(n_137),
.B2(n_117),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_31),
.C(n_17),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_131),
.B(n_31),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_177),
.B(n_183),
.Y(n_244)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_220),
.B(n_205),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_154),
.C(n_99),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_224),
.C(n_164),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_222),
.B1(n_226),
.B2(n_233),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_141),
.B1(n_102),
.B2(n_133),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_163),
.A2(n_118),
.B1(n_121),
.B2(n_129),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_154),
.C(n_99),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_159),
.A2(n_118),
.B1(n_117),
.B2(n_123),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_170),
.B1(n_201),
.B2(n_189),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_SL g236 ( 
.A1(n_174),
.A2(n_95),
.B(n_141),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_158),
.C(n_191),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_176),
.A2(n_132),
.B1(n_137),
.B2(n_123),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_132),
.B1(n_196),
.B2(n_144),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_174),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_239),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_179),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_174),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_216),
.C(n_237),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_249),
.Y(n_288)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_259),
.B(n_225),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_181),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_247),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_209),
.B(n_160),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_225),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_178),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_225),
.B(n_231),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_168),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_258),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_162),
.B(n_133),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_251),
.A2(n_256),
.B1(n_268),
.B2(n_269),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

AO21x1_ASAP7_75t_SL g253 ( 
.A1(n_212),
.A2(n_172),
.B(n_171),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_255),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_199),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_194),
.C(n_158),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_260),
.A2(n_266),
.B1(n_228),
.B2(n_234),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_158),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_232),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_144),
.B1(n_127),
.B2(n_120),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_231),
.B(n_182),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_267),
.B(n_232),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_227),
.A2(n_188),
.B1(n_165),
.B2(n_166),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_227),
.A2(n_166),
.B1(n_165),
.B2(n_148),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_R g329 ( 
.A(n_270),
.B(n_280),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_249),
.A2(n_221),
.B1(n_217),
.B2(n_215),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_253),
.B1(n_266),
.B2(n_227),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_273),
.A2(n_297),
.B1(n_269),
.B2(n_222),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_209),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_287),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_277),
.B(n_282),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_241),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_265),
.B(n_244),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_259),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_267),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_248),
.A2(n_211),
.B1(n_217),
.B2(n_215),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_300),
.B1(n_252),
.B2(n_210),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_224),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_298),
.C(n_246),
.Y(n_314)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_299),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_234),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_248),
.A2(n_204),
.B1(n_230),
.B2(n_219),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_243),
.Y(n_302)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_304),
.B(n_309),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_298),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_242),
.C(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_258),
.Y(n_312)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_245),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_313),
.B(n_323),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_322),
.C(n_327),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_238),
.Y(n_315)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_282),
.A2(n_240),
.B1(n_263),
.B2(n_256),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_275),
.B1(n_297),
.B2(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_325),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_320),
.A2(n_321),
.B1(n_328),
.B2(n_272),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_273),
.A2(n_262),
.B1(n_261),
.B2(n_254),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_255),
.C(n_223),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_289),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_234),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_326),
.A2(n_329),
.B1(n_295),
.B2(n_208),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_226),
.C(n_229),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_275),
.A2(n_233),
.B1(n_260),
.B2(n_208),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_279),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_303),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_333),
.B(n_350),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_338),
.B1(n_355),
.B2(n_357),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_274),
.C(n_270),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_343),
.C(n_346),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_277),
.B1(n_291),
.B2(n_300),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_307),
.A2(n_284),
.B1(n_281),
.B2(n_283),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_339),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_281),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_344),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_284),
.B1(n_294),
.B2(n_276),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_278),
.C(n_294),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_276),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_229),
.C(n_230),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_328),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_206),
.B1(n_295),
.B2(n_290),
.Y(n_348)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx3_ASAP7_75t_SL g349 ( 
.A(n_324),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_349),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_206),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_84),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_219),
.C(n_272),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_325),
.C(n_301),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_290),
.B1(n_210),
.B2(n_204),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_318),
.A2(n_290),
.B1(n_210),
.B2(n_204),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_358),
.A2(n_305),
.B1(n_301),
.B2(n_319),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_310),
.Y(n_362)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_337),
.A2(n_321),
.B(n_306),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_363),
.A2(n_374),
.B(n_377),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_375),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_371),
.B1(n_383),
.B2(n_385),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_369),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_376),
.C(n_378),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_338),
.A2(n_315),
.B1(n_312),
.B2(n_324),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_334),
.A2(n_316),
.B1(n_311),
.B2(n_305),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_148),
.C(n_173),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_354),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_349),
.A2(n_184),
.B(n_161),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_122),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_125),
.C(n_145),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_355),
.A2(n_169),
.B(n_167),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_153),
.C(n_145),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_382),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_153),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_332),
.B(n_12),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_335),
.A2(n_155),
.B1(n_55),
.B2(n_125),
.Y(n_385)
);

BUFx12_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_395),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_391),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_350),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_331),
.C(n_335),
.Y(n_393)
);

MAJx2_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_380),
.C(n_385),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_340),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_346),
.C(n_344),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_401),
.C(n_405),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_351),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_398),
.B(n_404),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_379),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_379),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_347),
.C(n_341),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_357),
.B1(n_358),
.B2(n_345),
.Y(n_403)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_356),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_361),
.B(n_341),
.C(n_345),
.Y(n_405)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_391),
.B(n_384),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_420),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_382),
.C(n_376),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_414),
.C(n_416),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_378),
.C(n_372),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_394),
.A2(n_363),
.B(n_384),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_418),
.B(n_421),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_372),
.C(n_371),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_377),
.B(n_370),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_370),
.C(n_360),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_398),
.C(n_89),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_394),
.A2(n_365),
.B(n_360),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_366),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_423),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_390),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_427),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_408),
.B(n_405),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_417),
.A2(n_388),
.B1(n_386),
.B2(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_428),
.Y(n_440)
);

AOI211xp5_ASAP7_75t_L g429 ( 
.A1(n_409),
.A2(n_383),
.B(n_387),
.C(n_400),
.Y(n_429)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_422),
.A2(n_386),
.B1(n_402),
.B2(n_387),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_431),
.B(n_434),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_395),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_436),
.C(n_438),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_69),
.C(n_72),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_14),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_14),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_0),
.C(n_1),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_421),
.B(n_407),
.Y(n_439)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_430),
.A2(n_423),
.B(n_416),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_439),
.B(n_451),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_414),
.B(n_413),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_442),
.A2(n_448),
.B(n_449),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_425),
.B(n_411),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_445),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_0),
.C(n_1),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_436),
.A2(n_14),
.B(n_13),
.Y(n_449)
);

AOI221xp5_ASAP7_75t_L g450 ( 
.A1(n_426),
.A2(n_11),
.B1(n_10),
.B2(n_12),
.C(n_3),
.Y(n_450)
);

OAI321xp33_ASAP7_75t_L g461 ( 
.A1(n_450),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.C(n_5),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_432),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_452),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_432),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_0),
.Y(n_465)
);

NAND3xp33_ASAP7_75t_SL g464 ( 
.A(n_457),
.B(n_458),
.C(n_0),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_447),
.A2(n_435),
.B(n_438),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_428),
.B(n_10),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_459),
.A2(n_456),
.B(n_453),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_5),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_461),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_455),
.A2(n_440),
.B1(n_444),
.B2(n_448),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_466),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_464),
.B(n_465),
.Y(n_468)
);

AOI211x1_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_454),
.B(n_452),
.C(n_460),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_469),
.A2(n_471),
.B(n_2),
.Y(n_473)
);

AOI321xp33_ASAP7_75t_L g471 ( 
.A1(n_467),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C(n_457),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_470),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_472),
.B(n_473),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_474),
.A2(n_468),
.B(n_2),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_2),
.C(n_5),
.Y(n_476)
);


endmodule