module fake_jpeg_14515_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_54),
.B(n_56),
.Y(n_144)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_59),
.Y(n_143)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_29),
.B(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_69),
.Y(n_135)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_95),
.Y(n_142)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_74),
.Y(n_149)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_53),
.Y(n_127)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_45),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_46),
.Y(n_153)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_9),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_31),
.B(n_9),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_38),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_51),
.B1(n_40),
.B2(n_44),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_105),
.A2(n_37),
.B1(n_32),
.B2(n_34),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_129),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_51),
.B1(n_40),
.B2(n_31),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_116),
.A2(n_133),
.B1(n_147),
.B2(n_156),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_60),
.A2(n_39),
.B1(n_46),
.B2(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_131),
.A2(n_64),
.B1(n_99),
.B2(n_97),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_51),
.B1(n_40),
.B2(n_46),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_35),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_152),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_57),
.A2(n_39),
.B1(n_46),
.B2(n_44),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_53),
.B(n_35),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_153),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_39),
.B1(n_44),
.B2(n_50),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_59),
.B(n_36),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_144),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_165),
.B(n_207),
.Y(n_236)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_72),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_167),
.B(n_215),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_169),
.Y(n_264)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_171),
.Y(n_263)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_174),
.B(n_179),
.Y(n_267)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_48),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_180),
.B(n_181),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_47),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_37),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_182),
.B(n_195),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_183),
.B(n_199),
.Y(n_271)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_185),
.A2(n_189),
.B1(n_193),
.B2(n_202),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_113),
.B(n_37),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_221),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_143),
.A2(n_100),
.B1(n_25),
.B2(n_42),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_192),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_131),
.A2(n_76),
.B1(n_66),
.B2(n_77),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_115),
.B(n_42),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_83),
.B1(n_87),
.B2(n_90),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_197),
.A2(n_211),
.B1(n_146),
.B2(n_126),
.Y(n_238)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_131),
.A2(n_74),
.B1(n_92),
.B2(n_101),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_136),
.B(n_43),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_133),
.A2(n_42),
.B1(n_25),
.B2(n_32),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_32),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_213),
.B(n_214),
.Y(n_240)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_106),
.B(n_104),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_107),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_219),
.Y(n_269)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_222),
.B1(n_149),
.B2(n_146),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_43),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_34),
.B(n_25),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_169),
.B(n_175),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_229),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_149),
.C(n_125),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_209),
.C(n_219),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_250),
.B1(n_187),
.B2(n_220),
.Y(n_277)
);

AOI22x1_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_110),
.B1(n_108),
.B2(n_86),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_245),
.Y(n_276)
);

AO22x2_ASAP7_75t_SL g250 ( 
.A1(n_208),
.A2(n_161),
.B1(n_119),
.B2(n_157),
.Y(n_250)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_119),
.B1(n_139),
.B2(n_34),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_181),
.B(n_222),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_186),
.B(n_139),
.CI(n_125),
.CON(n_255),
.SN(n_255)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_255),
.B(n_208),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_43),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_265),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_177),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_178),
.B(n_157),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_110),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_187),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_218),
.A2(n_21),
.B1(n_102),
.B2(n_128),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_21),
.B1(n_191),
.B2(n_0),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_293),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_277),
.A2(n_245),
.B1(n_272),
.B2(n_269),
.Y(n_336)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_198),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_284),
.B(n_305),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_285),
.A2(n_309),
.B(n_251),
.Y(n_332)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_168),
.B(n_176),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_315),
.B(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_205),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_292),
.B(n_297),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_212),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_216),
.B1(n_204),
.B2(n_170),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_310),
.B1(n_312),
.B2(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_166),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_171),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_301),
.Y(n_354)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_300),
.A2(n_318),
.B1(n_5),
.B2(n_6),
.Y(n_360)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_302),
.B(n_304),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_214),
.C(n_201),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_320),
.C(n_224),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_229),
.B(n_184),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_250),
.A2(n_164),
.B1(n_172),
.B2(n_102),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_306),
.A2(n_256),
.B1(n_253),
.B2(n_245),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_0),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_311),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_271),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_233),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_259),
.A2(n_191),
.B1(n_21),
.B2(n_0),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_255),
.B(n_0),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_313),
.B(n_319),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_250),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_1),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_317),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_247),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_16),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_234),
.B(n_1),
.C(n_2),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_223),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_335),
.C(n_339),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_330),
.B(n_335),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_332),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_344),
.B1(n_352),
.B2(n_360),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_243),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_336),
.A2(n_342),
.B1(n_343),
.B2(n_351),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g373 ( 
.A(n_338),
.B(n_290),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_274),
.B(n_248),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_230),
.C(n_253),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_346),
.C(n_347),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_284),
.A2(n_254),
.B1(n_270),
.B2(n_258),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_276),
.A2(n_258),
.B1(n_241),
.B2(n_228),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_241),
.B1(n_244),
.B2(n_226),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_232),
.C(n_244),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_274),
.B(n_231),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_231),
.C(n_242),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_356),
.C(n_359),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_313),
.A2(n_231),
.B(n_264),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_285),
.B(n_332),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_276),
.A2(n_226),
.B1(n_261),
.B2(n_239),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_295),
.A2(n_261),
.B1(n_239),
.B2(n_242),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_1),
.C(n_3),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_3),
.C(n_5),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_354),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_363),
.B(n_390),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_364),
.A2(n_373),
.B(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_326),
.Y(n_366)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_327),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_368),
.B(n_386),
.C(n_288),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_323),
.A2(n_355),
.B1(n_353),
.B2(n_334),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_369),
.A2(n_372),
.B1(n_325),
.B2(n_330),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_323),
.A2(n_319),
.B1(n_299),
.B2(n_293),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_308),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_374),
.B(n_379),
.C(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_275),
.Y(n_375)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_378),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_353),
.A2(n_286),
.B(n_320),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_338),
.A2(n_333),
.B(n_350),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_283),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_309),
.C(n_279),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_385),
.C(n_387),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_297),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_331),
.B(n_296),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_292),
.C(n_278),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_314),
.B1(n_310),
.B2(n_318),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_388),
.A2(n_345),
.B1(n_356),
.B2(n_300),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_324),
.B(n_315),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_398),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_357),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

XOR2x1_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_281),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_396),
.Y(n_410)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_305),
.C(n_302),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_294),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_324),
.B(n_301),
.Y(n_398)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_382),
.A2(n_354),
.B1(n_357),
.B2(n_348),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_405),
.B1(n_415),
.B2(n_423),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_403),
.A2(n_408),
.B1(n_424),
.B2(n_6),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_362),
.Y(n_404)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

OAI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_365),
.A2(n_344),
.B1(n_341),
.B2(n_343),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_369),
.A2(n_351),
.B1(n_346),
.B2(n_358),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_393),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_409),
.B(n_380),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_358),
.Y(n_413)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_364),
.A2(n_361),
.B1(n_300),
.B2(n_359),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_298),
.B1(n_291),
.B2(n_289),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_425),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_5),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_427),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_6),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_428),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_383),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_439),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_370),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_445),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_387),
.C(n_376),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_434),
.C(n_443),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_376),
.C(n_370),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_385),
.Y(n_435)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_414),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_419),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_374),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_410),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_427),
.Y(n_469)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_384),
.C(n_377),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_365),
.Y(n_444)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_403),
.B(n_392),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_411),
.A2(n_373),
.B(n_367),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_448),
.A2(n_408),
.B(n_407),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_377),
.C(n_389),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_429),
.C(n_428),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_417),
.B(n_388),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_413),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_453),
.A2(n_400),
.B1(n_417),
.B2(n_423),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_402),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_455),
.A2(n_420),
.B1(n_426),
.B2(n_400),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_458),
.A2(n_440),
.B(n_431),
.Y(n_490)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_461),
.B(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_464),
.B(n_466),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g467 ( 
.A(n_449),
.B(n_445),
.CI(n_435),
.CON(n_467),
.SN(n_467)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_467),
.Y(n_493)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_468),
.B(n_470),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_477),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_419),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_424),
.C(n_406),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_475),
.C(n_476),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_399),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_474),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_426),
.C(n_420),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_401),
.C(n_422),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_460),
.A2(n_447),
.B1(n_450),
.B2(n_436),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_479),
.A2(n_451),
.B1(n_476),
.B2(n_466),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_441),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_481),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_432),
.Y(n_481)
);

AOI21xp33_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_454),
.B(n_436),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_482),
.A2(n_483),
.B(n_458),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_465),
.A2(n_448),
.B(n_447),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_430),
.C(n_453),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_475),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_467),
.B(n_422),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_440),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_494),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_431),
.Y(n_494)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_465),
.C(n_457),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_496),
.B(n_499),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_488),
.A2(n_463),
.B1(n_450),
.B2(n_456),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_500),
.A2(n_480),
.B1(n_481),
.B2(n_13),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_492),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_501),
.B(n_503),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_502),
.A2(n_504),
.B1(n_491),
.B2(n_478),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_457),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_485),
.A2(n_467),
.B(n_455),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_506),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_401),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_502),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_8),
.C(n_9),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_509),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_11),
.C(n_12),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_500),
.A2(n_479),
.B1(n_493),
.B2(n_490),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_511),
.Y(n_524)
);

AOI21xp33_ASAP7_75t_L g512 ( 
.A1(n_498),
.A2(n_484),
.B(n_478),
.Y(n_512)
);

OA21x2_ASAP7_75t_SL g521 ( 
.A1(n_512),
.A2(n_496),
.B(n_497),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_518),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_11),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_515),
.Y(n_523)
);

AOI31xp33_ASAP7_75t_L g530 ( 
.A1(n_521),
.A2(n_526),
.A3(n_516),
.B(n_517),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_523),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_497),
.C(n_509),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_527),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_508),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_12),
.C(n_13),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_514),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_528),
.B(n_524),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_SL g533 ( 
.A1(n_530),
.A2(n_522),
.B(n_510),
.C(n_518),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_SL g534 ( 
.A1(n_532),
.A2(n_533),
.B(n_529),
.C(n_531),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_535),
.B(n_13),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_532),
.A2(n_520),
.B(n_527),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_536),
.B(n_13),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_14),
.B(n_15),
.Y(n_538)
);

OAI21xp33_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_14),
.B(n_15),
.Y(n_539)
);


endmodule