module real_jpeg_26351_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_2),
.B(n_76),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_2),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_2),
.B(n_51),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_2),
.B(n_32),
.C(n_64),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_67),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_210),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_2),
.B(n_25),
.C(n_27),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_2),
.A2(n_99),
.B(n_271),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g49 ( 
.A(n_4),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_5),
.A2(n_41),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_5),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_5),
.A2(n_52),
.B1(n_54),
.B2(n_142),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_142),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_142),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_39),
.B1(n_42),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_25),
.B1(n_28),
.B2(n_56),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_39),
.B1(n_77),
.B2(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_114),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_114),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_114),
.Y(n_241)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_60),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_60),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_60),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_11),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_43),
.B1(n_52),
.B2(n_54),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_43),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_52),
.B1(n_54),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_25),
.B1(n_28),
.B2(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_14),
.A2(n_77),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_14),
.A2(n_52),
.B1(n_54),
.B2(n_159),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_159),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_159),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_15),
.A2(n_36),
.B1(n_52),
.B2(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_25),
.B1(n_28),
.B2(n_36),
.Y(n_104)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_16),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_115),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_84),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_20),
.B(n_84),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.C(n_57),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_22),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_22),
.A2(n_57),
.B1(n_82),
.B2(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_23),
.A2(n_29),
.B1(n_96),
.B2(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_23),
.A2(n_29),
.B1(n_108),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_23),
.A2(n_29),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_23),
.B(n_207),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_24),
.A2(n_35),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_24),
.A2(n_94),
.B1(n_136),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_24),
.A2(n_170),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_24),
.A2(n_206),
.B(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_24),
.B(n_210),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_100),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_28),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_29),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_31),
.A2(n_32),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_32),
.B(n_278),
.Y(n_277)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_37),
.A2(n_72),
.B1(n_73),
.B2(n_83),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_37),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_50),
.B2(n_55),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_38),
.A2(n_50),
.B(n_111),
.Y(n_110)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_40),
.A2(n_48),
.A3(n_54),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_41),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_50),
.B1(n_55),
.B2(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_44),
.A2(n_140),
.B(n_144),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_45),
.A2(n_51),
.B1(n_141),
.B2(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_45),
.A2(n_145),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_47),
.B(n_52),
.Y(n_187)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_113),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_50),
.A2(n_111),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_52),
.B(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_61),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_61),
.A2(n_67),
.B1(n_178),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_63),
.B1(n_69),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_62),
.A2(n_63),
.B1(n_92),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_62),
.A2(n_177),
.B(n_179),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_62),
.A2(n_179),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_63),
.A2(n_138),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_63),
.A2(n_163),
.B(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_67),
.B(n_164),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_77),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_97),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_94),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_94),
.A2(n_259),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_147),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_105),
.B(n_109),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_109),
.B1(n_110),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_98),
.A2(n_106),
.B1(n_107),
.B2(n_122),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B(n_104),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_104),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_99),
.A2(n_101),
.B1(n_130),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_99),
.A2(n_100),
.B1(n_184),
.B2(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_99),
.B(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_99),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_100),
.Y(n_284)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_102),
.B(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_103),
.B(n_210),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_149),
.B(n_327),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_146),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_119),
.B(n_146),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_120),
.Y(n_323)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_125),
.A2(n_126),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.C(n_139),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_127),
.A2(n_128),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_168),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_137),
.B(n_139),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_320),
.B(n_326),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_195),
.B(n_319),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_188),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_152),
.B(n_188),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_171),
.C(n_173),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_153),
.A2(n_154),
.B1(n_171),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_161),
.C(n_165),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_169),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_171),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_173),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_176),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_180),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_182),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_190),
.B(n_191),
.C(n_194),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_226),
.B(n_313),
.C(n_318),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_220),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_220),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_212),
.C(n_213),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_198),
.A2(n_199),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_204),
.C(n_208),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_212),
.B(n_213),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_307),
.B(n_312),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_260),
.B(n_306),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_249),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_249),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_242),
.C(n_246),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_232),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B(n_240),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_283),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_242),
.A2(n_246),
.B1(n_247),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_254),
.B2(n_255),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_256),
.C(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_300),
.B(n_305),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_279),
.B(n_299),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_273),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_273),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_277),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_288),
.B(n_298),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_286),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_293),
.B(n_297),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_304),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_311),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_311),
.Y(n_312)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule