module fake_jpeg_13063_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_52),
.B1(n_34),
.B2(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_33),
.B1(n_26),
.B2(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_64),
.Y(n_102)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx11_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_72),
.Y(n_88)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_85),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_29),
.C(n_32),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_34),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_57),
.B1(n_65),
.B2(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_91),
.B1(n_103),
.B2(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_94),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_18),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_42),
.B1(n_43),
.B2(n_37),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_98),
.B1(n_39),
.B2(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_37),
.B1(n_43),
.B2(n_42),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_18),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_21),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_30),
.B1(n_35),
.B2(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_104),
.B(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_89),
.B1(n_77),
.B2(n_27),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_108),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_96),
.A3(n_86),
.B1(n_84),
.B2(n_101),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_118),
.Y(n_133)
);

INVxp67_ASAP7_75t_SL g134 ( 
.A(n_112),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_130),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_129),
.B(n_1),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_71),
.B1(n_69),
.B2(n_59),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_125),
.B1(n_98),
.B2(n_100),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_46),
.A3(n_23),
.B1(n_62),
.B2(n_61),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_61),
.B(n_30),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_31),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_18),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_83),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_71),
.B1(n_27),
.B2(n_20),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_46),
.B1(n_24),
.B2(n_62),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_61),
.B1(n_62),
.B2(n_27),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_76),
.B(n_23),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_23),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_73),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_155),
.B(n_156),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_76),
.B(n_94),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_142),
.B1(n_116),
.B2(n_123),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_92),
.B1(n_89),
.B2(n_74),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_147),
.B1(n_150),
.B2(n_115),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_119),
.B1(n_113),
.B2(n_109),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_77),
.C(n_74),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_153),
.C(n_131),
.Y(n_184)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_81),
.B(n_35),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_4),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_111),
.B1(n_108),
.B2(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_23),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_158),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_83),
.C(n_62),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_24),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_23),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_161),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_1),
.B(n_3),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_0),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_61),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_160),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_176),
.B1(n_192),
.B2(n_155),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_118),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_184),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_170),
.B(n_172),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_122),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_120),
.B1(n_125),
.B2(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_138),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_131),
.B1(n_117),
.B2(n_112),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_148),
.B1(n_147),
.B2(n_6),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_140),
.B(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_117),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_4),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_22),
.B1(n_10),
.B2(n_11),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_161),
.B(n_156),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_10),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_164),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_22),
.B1(n_11),
.B2(n_12),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_9),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_196),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_133),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_8),
.C(n_13),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_134),
.B(n_133),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_223),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_145),
.B(n_139),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NAND2x1_ASAP7_75t_SL g210 ( 
.A(n_168),
.B(n_164),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_211),
.B(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_185),
.A2(n_155),
.B1(n_137),
.B2(n_157),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_173),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_171),
.B(n_154),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_176),
.B1(n_192),
.B2(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_222),
.A2(n_173),
.B1(n_191),
.B2(n_166),
.Y(n_243)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_225),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_184),
.C(n_169),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_236),
.C(n_216),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_215),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_234),
.A2(n_243),
.B1(n_244),
.B2(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_193),
.C(n_197),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_196),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_208),
.B(n_167),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_242),
.B(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_181),
.B1(n_180),
.B2(n_174),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_201),
.B(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_263),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_209),
.B1(n_221),
.B2(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_234),
.B1(n_244),
.B2(n_239),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_270),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_216),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_251),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_206),
.C(n_211),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_200),
.C(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_203),
.C(n_220),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_220),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_272),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_213),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_268),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_219),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_250),
.B(n_210),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_251),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_203),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_238),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_251),
.C(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_287),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_243),
.B(n_246),
.Y(n_282)
);

OAI21x1_ASAP7_75t_SL g294 ( 
.A1(n_282),
.A2(n_271),
.B(n_267),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_239),
.C(n_222),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_278),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_207),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_245),
.C(n_212),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_245),
.C(n_253),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_265),
.C(n_273),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_240),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_265),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_300),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_301),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_259),
.B(n_264),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_275),
.B(n_287),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_269),
.B1(n_209),
.B2(n_270),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_283),
.B1(n_284),
.B2(n_222),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_202),
.C(n_238),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_240),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_235),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_288),
.Y(n_310)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_235),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_316),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_317),
.B(n_318),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.Y(n_320)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_314),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_298),
.A2(n_283),
.B1(n_202),
.B2(n_223),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_303),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_223),
.B1(n_9),
.B2(n_7),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_7),
.C(n_12),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_293),
.C(n_292),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_297),
.C(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_5),
.B(n_6),
.Y(n_333)
);

AOI221xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_299),
.B1(n_302),
.B2(n_12),
.C(n_7),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_317),
.B1(n_13),
.B2(n_16),
.Y(n_331)
);

OA21x2_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_311),
.B(n_310),
.Y(n_330)
);

OAI311xp33_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_329),
.A3(n_327),
.B1(n_320),
.C1(n_328),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_4),
.C(n_5),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_326),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_335),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_330),
.C(n_334),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_320),
.B1(n_5),
.B2(n_6),
.Y(n_340)
);


endmodule