module fake_jpeg_1669_n_455 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_455);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_48),
.Y(n_108)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_20),
.A2(n_8),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_6),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_24),
.Y(n_100)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_114),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_0),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_40),
.B1(n_29),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_125),
.B1(n_31),
.B2(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_45),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_45),
.B1(n_44),
.B2(n_26),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_87),
.B1(n_83),
.B2(n_74),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_41),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_129),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_48),
.A2(n_40),
.B1(n_39),
.B2(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_49),
.B(n_44),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_30),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_145),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_39),
.C(n_33),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_31),
.C(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_69),
.B(n_34),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_9),
.Y(n_189)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_106),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_156),
.B(n_165),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_158),
.A2(n_168),
.B1(n_170),
.B2(n_179),
.Y(n_225)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_160),
.B(n_162),
.Y(n_236)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_67),
.A3(n_21),
.B1(n_38),
.B2(n_43),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_40),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_38),
.B1(n_68),
.B2(n_64),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_112),
.A2(n_50),
.B1(n_63),
.B2(n_60),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_176),
.B(n_189),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_97),
.A2(n_125),
.B1(n_53),
.B2(n_57),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

AND2x4_ASAP7_75t_SL g172 ( 
.A(n_96),
.B(n_71),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_172),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_109),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_109),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_35),
.B1(n_23),
.B2(n_17),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_101),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_193),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_117),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_128),
.B1(n_121),
.B2(n_148),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_119),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_126),
.B(n_6),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_147),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_197),
.Y(n_235)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_131),
.A2(n_5),
.A3(n_13),
.B1(n_11),
.B2(n_3),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_11),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_199),
.Y(n_228)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx6p67_ASAP7_75t_R g200 ( 
.A(n_137),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_147),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_160),
.C(n_188),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_205),
.C(n_200),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_110),
.B1(n_127),
.B2(n_120),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_204),
.A2(n_227),
.B1(n_174),
.B2(n_141),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_150),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_222),
.B1(n_128),
.B2(n_185),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_220),
.A2(n_153),
.B1(n_184),
.B2(n_157),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_148),
.B1(n_113),
.B2(n_124),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_169),
.A2(n_172),
.B1(n_127),
.B2(n_196),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_180),
.B(n_142),
.CI(n_115),
.CON(n_231),
.SN(n_231)
);

AOI32xp33_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_141),
.A3(n_138),
.B1(n_4),
.B2(n_3),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_172),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_199),
.B1(n_175),
.B2(n_113),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_242),
.A2(n_254),
.B1(n_220),
.B2(n_202),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_244),
.B(n_260),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_155),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_250),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_178),
.B(n_152),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_247),
.A2(n_267),
.B(n_240),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_151),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_159),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_236),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_273),
.B1(n_249),
.B2(n_220),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_124),
.B1(n_164),
.B2(n_177),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_144),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_258),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_261),
.C(n_260),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_203),
.B(n_167),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_182),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_200),
.C(n_171),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_194),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_265),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_264),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_200),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_266),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_187),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_272),
.Y(n_285)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_211),
.A2(n_9),
.B(n_14),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_220),
.B(n_210),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_225),
.B(n_138),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_225),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_275),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_204),
.A2(n_3),
.B1(n_4),
.B2(n_10),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_237),
.B1(n_233),
.B2(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_278),
.A2(n_288),
.B1(n_307),
.B2(n_273),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_250),
.A2(n_211),
.B1(n_240),
.B2(n_231),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_295),
.A2(n_266),
.B(n_207),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_268),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_243),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_298),
.A2(n_256),
.B1(n_275),
.B2(n_269),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_234),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_305),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_235),
.B1(n_231),
.B2(n_209),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_244),
.B1(n_247),
.B2(n_253),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_207),
.C(n_201),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_255),
.C(n_246),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_263),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_312),
.B(n_318),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_313),
.A2(n_328),
.B1(n_334),
.B2(n_337),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_270),
.B(n_271),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_314),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_276),
.B(n_261),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_321),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_280),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_323),
.Y(n_351)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_282),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_327),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_237),
.B1(n_229),
.B2(n_277),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_307),
.B1(n_289),
.B2(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_274),
.B1(n_262),
.B2(n_264),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_264),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_329),
.Y(n_356)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_331),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_297),
.B(n_245),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_293),
.B(n_245),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_338),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_333),
.A2(n_339),
.B1(n_287),
.B2(n_290),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_294),
.A2(n_229),
.B1(n_217),
.B2(n_216),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_233),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_335),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_294),
.A2(n_217),
.B1(n_201),
.B2(n_230),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_213),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_283),
.B1(n_308),
.B2(n_300),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_306),
.C(n_305),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_353),
.C(n_365),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_308),
.B1(n_300),
.B2(n_288),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_297),
.B1(n_285),
.B2(n_299),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_320),
.C(n_309),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_352),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_285),
.B1(n_291),
.B2(n_279),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_350),
.A2(n_358),
.B1(n_364),
.B2(n_332),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_303),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_357),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_301),
.C(n_289),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_301),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_314),
.A2(n_318),
.B1(n_319),
.B2(n_322),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_359),
.A2(n_364),
.B1(n_351),
.B2(n_356),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_312),
.A2(n_287),
.B1(n_290),
.B2(n_302),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_329),
.C(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g368 ( 
.A1(n_341),
.A2(n_319),
.B(n_315),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_321),
.C(n_335),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_370),
.C(n_381),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_333),
.C(n_325),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_371),
.A2(n_377),
.B1(n_380),
.B2(n_382),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_385),
.Y(n_398)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_375),
.Y(n_401)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_311),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_378),
.B(n_383),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_343),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_379),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_SL g380 ( 
.A(n_341),
.B(n_331),
.C(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_330),
.C(n_327),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_355),
.A2(n_328),
.B1(n_326),
.B2(n_334),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_361),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_323),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_302),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_363),
.B(n_342),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_376),
.B(n_345),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_389),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_350),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_357),
.C(n_360),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_392),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_360),
.C(n_359),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_396),
.Y(n_417)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_358),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_402),
.C(n_371),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_340),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_347),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_366),
.C(n_381),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_405),
.B(n_411),
.Y(n_428)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_388),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_362),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_401),
.Y(n_407)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

AO21x1_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_377),
.B(n_375),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_416),
.Y(n_426)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_412),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_400),
.A2(n_379),
.B1(n_385),
.B2(n_382),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_389),
.C(n_391),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_373),
.C(n_372),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_416),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_374),
.C(n_368),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_392),
.C(n_402),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_422),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_387),
.C(n_398),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_404),
.A2(n_347),
.B1(n_403),
.B2(n_368),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_423),
.A2(n_429),
.B(n_292),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_414),
.A2(n_395),
.B(n_393),
.Y(n_424)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_426),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_427),
.B(n_415),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_337),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_418),
.B(n_417),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_431),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_408),
.C(n_290),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_433),
.B(n_434),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_292),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_292),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_436),
.B(n_419),
.Y(n_443)
);

AO21x1_ASAP7_75t_L g439 ( 
.A1(n_437),
.A2(n_426),
.B(n_423),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_443),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_420),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_441),
.A2(n_444),
.B(n_434),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_428),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_435),
.B(n_432),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_445),
.A2(n_446),
.B(n_436),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_442),
.A2(n_437),
.B(n_429),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_213),
.Y(n_450)
);

OAI31xp33_ASAP7_75t_SL g451 ( 
.A1(n_449),
.A2(n_450),
.A3(n_447),
.B(n_230),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_4),
.C(n_14),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_0),
.B(n_1),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_0),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_1),
.B1(n_388),
.B2(n_419),
.Y(n_455)
);


endmodule