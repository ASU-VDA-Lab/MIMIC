module real_jpeg_20634_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_5),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_2),
.A2(n_5),
.B1(n_26),
.B2(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_2),
.A2(n_3),
.B1(n_41),
.B2(n_60),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_2),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_64),
.B(n_70),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_2),
.B(n_75),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_2),
.A2(n_35),
.B(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_61),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_3),
.A2(n_8),
.B1(n_39),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_41),
.B(n_65),
.C(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_5),
.B(n_24),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_5),
.A2(n_7),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_5),
.A2(n_10),
.B1(n_26),
.B2(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_5),
.A2(n_8),
.B1(n_26),
.B2(n_39),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_60),
.B(n_62),
.C(n_69),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_110),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_109),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_97),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_16),
.B(n_97),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_96),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_43),
.B2(n_44),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_31),
.B2(n_42),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_23),
.A2(n_24),
.B1(n_49),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_23),
.B(n_28),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_28),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_26),
.B(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_28),
.B(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_31),
.A2(n_42),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_31),
.B(n_90),
.C(n_140),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_31),
.A2(n_42),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_31),
.B(n_160),
.C(n_169),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_32),
.B(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_34),
.A2(n_35),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_35),
.A2(n_36),
.B(n_41),
.C(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_37),
.B(n_41),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_41),
.A2(n_64),
.B(n_78),
.C(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_56),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_46),
.A2(n_51),
.B1(n_52),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_46),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_47),
.A2(n_91),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_48),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_51),
.A2(n_52),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_51),
.A2(n_52),
.B1(n_104),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_52),
.B(n_125),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_52),
.B(n_104),
.C(n_147),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_57),
.A2(n_58),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_104),
.C(n_106),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_66),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_61),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_76),
.B(n_77),
.C(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_77),
.Y(n_81)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_76),
.B1(n_80),
.B2(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_95),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.C(n_92),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_132),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_92),
.A2(n_93),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_93),
.B(n_120),
.C(n_163),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.C(n_103),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_98),
.B(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_101),
.B(n_103),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_104),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_104),
.A2(n_106),
.B1(n_155),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_186),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_182),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_171),
.B(n_181),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_157),
.B(n_170),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_144),
.B(n_156),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_135),
.B(n_143),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_127),
.B(n_134),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_120),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_131),
.B(n_133),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_153),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_168),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_173),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);


endmodule