module fake_jpeg_9155_n_60 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_16),
.C(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_17),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_11),
.B(n_12),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_10),
.B(n_16),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_23),
.B(n_20),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.C(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_20),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_9),
.B1(n_14),
.B2(n_21),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_21),
.B1(n_7),
.B2(n_8),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_35),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_35),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_44),
.B(n_45),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_21),
.B1(n_17),
.B2(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_7),
.C(n_4),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_40),
.C(n_5),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_51),
.Y(n_55)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_43),
.B1(n_47),
.B2(n_45),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_54),
.B(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.C(n_54),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_49),
.C(n_3),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_53),
.C(n_6),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_6),
.Y(n_60)
);


endmodule