module fake_jpeg_21663_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_11),
.B1(n_17),
.B2(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_38),
.B1(n_20),
.B2(n_29),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_20),
.B1(n_11),
.B2(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_9),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_37),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_26),
.B1(n_21),
.B2(n_10),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_26),
.B1(n_17),
.B2(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_41),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_47),
.B1(n_42),
.B2(n_10),
.C(n_16),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_69),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_57),
.B1(n_42),
.B2(n_53),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_21),
.B1(n_17),
.B2(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_55),
.B(n_58),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_81),
.B(n_5),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_14),
.B1(n_12),
.B2(n_22),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_14),
.C(n_7),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_14),
.C(n_8),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_7),
.B(n_8),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI321xp33_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_69),
.A3(n_70),
.B1(n_67),
.B2(n_22),
.C(n_4),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_77),
.B(n_6),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_22),
.C(n_12),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_78),
.B1(n_76),
.B2(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_93),
.B1(n_5),
.B2(n_9),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_78),
.C(n_22),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_88),
.C(n_15),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_4),
.B(n_6),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_99),
.B(n_0),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_12),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_5),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_9),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_95),
.C(n_92),
.Y(n_104)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_104),
.C(n_97),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_1),
.B(n_2),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_92),
.C(n_2),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.B(n_2),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_3),
.B(n_109),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_110),
.Y(n_111)
);


endmodule