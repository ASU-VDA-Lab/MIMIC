module fake_jpeg_11166_n_307 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_29),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_24),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_34),
.B1(n_22),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_26),
.B1(n_22),
.B2(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_17),
.B1(n_29),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_26),
.B1(n_39),
.B2(n_45),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_26),
.B(n_30),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_64),
.B(n_36),
.C(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_46),
.B1(n_62),
.B2(n_24),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_17),
.B1(n_20),
.B2(n_32),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_26),
.B(n_30),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_95),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_73),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_77),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_84),
.B1(n_94),
.B2(n_33),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_45),
.B1(n_44),
.B2(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_53),
.B1(n_55),
.B2(n_60),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_37),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_36),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_32),
.B1(n_20),
.B2(n_21),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_102),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_44),
.B1(n_37),
.B2(n_36),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_104),
.B(n_87),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_49),
.B1(n_66),
.B2(n_88),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_89),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_63),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_61),
.C(n_68),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_102),
.B1(n_79),
.B2(n_101),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_118),
.C(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_68),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_73),
.C(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_89),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_140),
.B1(n_146),
.B2(n_156),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_150),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_120),
.C(n_115),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_18),
.Y(n_187)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_139),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_84),
.B1(n_61),
.B2(n_66),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_148),
.Y(n_169)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_66),
.B1(n_49),
.B2(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_95),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_151),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_92),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_75),
.A3(n_57),
.B1(n_21),
.B2(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_158),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_155),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_49),
.B1(n_21),
.B2(n_28),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_161),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_33),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_110),
.A2(n_28),
.B1(n_83),
.B2(n_71),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_112),
.B1(n_109),
.B2(n_117),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_105),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_123),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_188),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_180),
.B1(n_144),
.B2(n_147),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_176),
.B1(n_6),
.B2(n_14),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_130),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_183),
.C(n_190),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_152),
.B1(n_145),
.B2(n_133),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_109),
.B(n_126),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_189),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_109),
.B1(n_128),
.B2(n_126),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_158),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_57),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_24),
.B(n_18),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_187),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_80),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_18),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_7),
.C(n_15),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_0),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_134),
.B(n_7),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_9),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_156),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_183),
.C(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_150),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_197),
.B(n_205),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_146),
.B(n_139),
.C(n_153),
.D(n_140),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_204),
.B(n_219),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_158),
.B1(n_138),
.B2(n_143),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_7),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_9),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_165),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_185),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_9),
.B1(n_15),
.B2(n_2),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_12),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_164),
.B1(n_163),
.B2(n_187),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_6),
.B(n_13),
.C(n_3),
.D(n_4),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_217),
.B1(n_213),
.B2(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_178),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_238),
.C(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_164),
.B1(n_170),
.B2(n_180),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_236),
.B1(n_241),
.B2(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_171),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_182),
.C(n_173),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_187),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_199),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_253),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_194),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_201),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_202),
.C(n_203),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_231),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_206),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_258),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_206),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_234),
.B1(n_220),
.B2(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_267),
.B1(n_226),
.B2(n_239),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_228),
.B(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_271),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_240),
.B1(n_223),
.B2(n_235),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_230),
.B(n_237),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

OAI211xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_272),
.B(n_268),
.C(n_262),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_248),
.B(n_221),
.CI(n_218),
.CON(n_272),
.SN(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_243),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_282),
.Y(n_284)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_277),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_242),
.C(n_258),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_280),
.B(n_259),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_255),
.C(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_249),
.B(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_225),
.B1(n_223),
.B2(n_235),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_181),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_283),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_219),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_286),
.B(n_287),
.Y(n_292)
);

OA21x2_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_272),
.B(n_270),
.Y(n_291)
);

OAI221xp5_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_222),
.B1(n_6),
.B2(n_3),
.C(n_4),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_294),
.B(n_5),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_283),
.A3(n_230),
.B1(n_261),
.B2(n_175),
.C1(n_270),
.C2(n_172),
.Y(n_293)
);

AOI31xp67_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_296),
.A3(n_297),
.B(n_10),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_186),
.B(n_175),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_284),
.Y(n_299)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_300),
.B(n_301),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_284),
.B(n_4),
.C(n_5),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_12),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_303),
.B(n_16),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_0),
.C(n_1),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_1),
.Y(n_307)
);


endmodule