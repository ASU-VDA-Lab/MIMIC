module fake_jpeg_2990_n_614 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_614);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_614;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_105),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_62),
.Y(n_169)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_75),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_96),
.Y(n_131)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_81),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_82),
.Y(n_216)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g135 ( 
.A(n_84),
.Y(n_135)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_0),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_92),
.A2(n_118),
.B(n_39),
.C(n_43),
.Y(n_185)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_94),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_95),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_97),
.Y(n_193)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_52),
.Y(n_140)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_102),
.Y(n_218)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_18),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx2_ASAP7_75t_SL g202 ( 
.A(n_111),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_1),
.C(n_2),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_49),
.C(n_41),
.Y(n_190)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_34),
.B(n_1),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_23),
.Y(n_124)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_129),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_53),
.B1(n_34),
.B2(n_43),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_137),
.A2(n_139),
.B1(n_213),
.B2(n_32),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_90),
.B1(n_85),
.B2(n_75),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_140),
.B(n_145),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_66),
.A2(n_52),
.B1(n_51),
.B2(n_55),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_111),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_155),
.A2(n_161),
.B1(n_174),
.B2(n_200),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_69),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_77),
.B(n_39),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_163),
.B(n_184),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_72),
.A2(n_58),
.B1(n_56),
.B2(n_54),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_70),
.B(n_52),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_196),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_65),
.B(n_54),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_189),
.B(n_192),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_190),
.B(n_220),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_83),
.B(n_87),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_88),
.B(n_49),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_195),
.B(n_207),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_68),
.B(n_41),
.Y(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_198),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_71),
.A2(n_47),
.B1(n_51),
.B2(n_40),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_205),
.Y(n_253)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_81),
.B(n_40),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_82),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_122),
.Y(n_249)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_95),
.A2(n_47),
.B1(n_32),
.B2(n_37),
.Y(n_213)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_127),
.B(n_32),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g222 ( 
.A(n_202),
.Y(n_222)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_222),
.Y(n_340)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_223),
.A2(n_158),
.B1(n_141),
.B2(n_172),
.Y(n_337)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_171),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_162),
.A2(n_44),
.B(n_3),
.C(n_4),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_231),
.B(n_6),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_244),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_234),
.Y(n_333)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g356 ( 
.A(n_235),
.Y(n_356)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_237),
.B(n_238),
.Y(n_309)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_239),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_154),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_240),
.Y(n_353)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_131),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_140),
.A2(n_44),
.B(n_4),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_247),
.A2(n_265),
.B(n_155),
.Y(n_303)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_259),
.Y(n_318)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_250),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_2),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_251),
.B(n_256),
.Y(n_310)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_135),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_2),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_159),
.Y(n_258)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_258),
.Y(n_352)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_178),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_261),
.Y(n_315)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_263),
.Y(n_317)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_143),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_189),
.A2(n_44),
.B(n_114),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_268),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_147),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_267),
.Y(n_312)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_269),
.B(n_271),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_149),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_270),
.Y(n_344)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_182),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_163),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_272),
.B(n_273),
.Y(n_341)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_130),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_160),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_274),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_184),
.A2(n_119),
.B1(n_110),
.B2(n_108),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_167),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_145),
.A2(n_104),
.B1(n_5),
.B2(n_6),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_194),
.B1(n_199),
.B2(n_193),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_166),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_347)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_183),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_134),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_196),
.A2(n_194),
.B1(n_201),
.B2(n_209),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_168),
.B1(n_221),
.B2(n_164),
.Y(n_314)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_142),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_286),
.B(n_289),
.Y(n_328)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_187),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_288),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_179),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_146),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_152),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_290),
.B(n_294),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_179),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_293),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_165),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_136),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_148),
.B(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_296),
.B(n_298),
.Y(n_348)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_165),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_303),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_306),
.A2(n_325),
.B1(n_327),
.B2(n_332),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_227),
.A2(n_221),
.B1(n_164),
.B2(n_186),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_313),
.A2(n_330),
.B1(n_349),
.B2(n_283),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_314),
.A2(n_327),
.B1(n_332),
.B2(n_324),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g316 ( 
.A(n_297),
.B(n_150),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_316),
.Y(n_386)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_229),
.A2(n_200),
.A3(n_169),
.B1(n_186),
.B2(n_181),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_342),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_227),
.A2(n_223),
.B1(n_285),
.B2(n_297),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_265),
.A2(n_216),
.B1(n_191),
.B2(n_214),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_279),
.A2(n_247),
.B1(n_291),
.B2(n_231),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_264),
.B(n_246),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_331),
.B(n_343),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_275),
.A2(n_216),
.B1(n_214),
.B2(n_181),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_284),
.B(n_215),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_338),
.C(n_354),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_337),
.A2(n_314),
.B1(n_305),
.B2(n_340),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_224),
.B(n_172),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_228),
.B(n_6),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_225),
.B(n_18),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_284),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_284),
.A2(n_8),
.B(n_9),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_350),
.A2(n_347),
.B(n_351),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_239),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_351),
.A2(n_240),
.B1(n_293),
.B2(n_292),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_236),
.B(n_226),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_268),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_358),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_333),
.B(n_263),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_350),
.A2(n_303),
.B1(n_330),
.B2(n_336),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_360),
.A2(n_361),
.B1(n_363),
.B2(n_373),
.Y(n_412)
);

A2O1A1O1Ixp25_ASAP7_75t_L g365 ( 
.A1(n_331),
.A2(n_255),
.B(n_253),
.C(n_233),
.D(n_230),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_365),
.A2(n_385),
.B(n_396),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_233),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_369),
.Y(n_415)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_310),
.B(n_243),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_253),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_371),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_245),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_248),
.B1(n_288),
.B2(n_242),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_341),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_380),
.Y(n_425)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_325),
.A2(n_235),
.B1(n_287),
.B2(n_241),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_377),
.A2(n_356),
.B1(n_302),
.B2(n_301),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_313),
.A2(n_295),
.B1(n_261),
.B2(n_14),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_381),
.B1(n_382),
.B2(n_391),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_11),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_384),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_309),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_306),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_323),
.A2(n_13),
.B1(n_15),
.B2(n_316),
.Y(n_382)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_318),
.B(n_13),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_328),
.B(n_317),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_310),
.B(n_338),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_395),
.Y(n_409)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_316),
.A2(n_337),
.B1(n_300),
.B2(n_322),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_321),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_309),
.B(n_346),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_354),
.B(n_342),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_397),
.Y(n_435)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_398),
.Y(n_437)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_SL g400 ( 
.A(n_316),
.B(n_329),
.C(n_337),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_364),
.C(n_386),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_344),
.A2(n_305),
.B(n_346),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_401),
.A2(n_299),
.B(n_311),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_337),
.B1(n_343),
.B2(n_344),
.Y(n_403)
);

OAI22x1_ASAP7_75t_L g454 ( 
.A1(n_403),
.A2(n_385),
.B1(n_370),
.B2(n_366),
.Y(n_454)
);

AND2x2_ASAP7_75t_SL g404 ( 
.A(n_364),
.B(n_335),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_404),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_360),
.A2(n_315),
.B(n_301),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_365),
.B(n_368),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_406),
.A2(n_373),
.B1(n_389),
.B2(n_394),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_357),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_339),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_410),
.B(n_387),
.Y(n_456)
);

OAI31xp33_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_428),
.A3(n_400),
.B(n_386),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_326),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_390),
.C(n_376),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_362),
.A2(n_324),
.B1(n_302),
.B2(n_355),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_420),
.A2(n_422),
.B1(n_431),
.B2(n_432),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_393),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_424),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_362),
.A2(n_355),
.B1(n_320),
.B2(n_299),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_401),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_319),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_359),
.A2(n_383),
.B1(n_368),
.B2(n_367),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_359),
.A2(n_320),
.B1(n_353),
.B2(n_326),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_361),
.A2(n_356),
.B1(n_312),
.B2(n_335),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_436),
.A2(n_358),
.B1(n_371),
.B2(n_379),
.Y(n_461)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_438),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_423),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_447),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_459),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_445),
.A2(n_460),
.B(n_462),
.Y(n_476)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_425),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_SL g500 ( 
.A(n_446),
.B(n_454),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_433),
.A2(n_382),
.B(n_369),
.C(n_368),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_380),
.Y(n_448)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_450),
.A2(n_428),
.B(n_415),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_416),
.A2(n_365),
.B1(n_434),
.B2(n_411),
.Y(n_451)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_416),
.A2(n_403),
.B1(n_412),
.B2(n_413),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_461),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_431),
.A2(n_396),
.B1(n_377),
.B2(n_395),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_385),
.B1(n_363),
.B2(n_374),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_471),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_430),
.B(n_375),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_457),
.B(n_407),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_466),
.C(n_470),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_409),
.B(n_392),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_433),
.A2(n_405),
.B(n_417),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_408),
.A2(n_378),
.B(n_394),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_418),
.B(n_374),
.Y(n_463)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_413),
.A2(n_384),
.B1(n_381),
.B2(n_353),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_464),
.A2(n_465),
.B1(n_472),
.B2(n_406),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_422),
.A2(n_397),
.B1(n_312),
.B2(n_352),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_352),
.C(n_334),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_397),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_414),
.B(n_334),
.Y(n_469)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_404),
.B(n_399),
.C(n_419),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_399),
.C(n_409),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_414),
.B1(n_427),
.B2(n_420),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_415),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_475),
.B(n_482),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_478),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_467),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_480),
.B(n_484),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_471),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_459),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_491),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_448),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_492),
.B(n_495),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_450),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g528 ( 
.A(n_493),
.B(n_494),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_444),
.B(n_418),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_440),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_496),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_463),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_499),
.B1(n_502),
.B2(n_503),
.Y(n_510)
);

OA22x2_ASAP7_75t_L g498 ( 
.A1(n_449),
.A2(n_428),
.B1(n_427),
.B2(n_432),
.Y(n_498)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_498),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_472),
.Y(n_501)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_402),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_482),
.C(n_473),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_485),
.C(n_494),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_486),
.A2(n_454),
.B1(n_455),
.B2(n_449),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_505),
.A2(n_513),
.B1(n_521),
.B2(n_523),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_474),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_511),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_470),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_445),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_519),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_486),
.A2(n_453),
.B1(n_441),
.B2(n_462),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_481),
.A2(n_428),
.B1(n_461),
.B2(n_447),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_515),
.B(n_493),
.Y(n_547)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_516),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_475),
.B(n_428),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_520),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_497),
.A2(n_465),
.B1(n_464),
.B2(n_402),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_481),
.A2(n_468),
.B1(n_439),
.B2(n_438),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_485),
.A2(n_439),
.B1(n_437),
.B2(n_423),
.Y(n_525)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_525),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_499),
.A2(n_429),
.B1(n_435),
.B2(n_426),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_498),
.Y(n_538)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_527),
.Y(n_543)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_529),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_476),
.B(n_407),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_530),
.B(n_476),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_536),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_507),
.B(n_512),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_537),
.B(n_546),
.Y(n_567)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_538),
.Y(n_558)
);

XNOR2x1_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_493),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_539),
.B(n_545),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_507),
.B(n_489),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_547),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_496),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_504),
.B(n_493),
.C(n_487),
.Y(n_546)
);

BUFx24_ASAP7_75t_SL g548 ( 
.A(n_517),
.Y(n_548)
);

BUFx24_ASAP7_75t_SL g559 ( 
.A(n_548),
.Y(n_559)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_549),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_518),
.B(n_484),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_550),
.A2(n_522),
.B(n_489),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_540),
.A2(n_510),
.B1(n_521),
.B2(n_513),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_551),
.A2(n_557),
.B1(n_563),
.B2(n_480),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_509),
.C(n_511),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_552),
.B(n_553),
.C(n_554),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_519),
.C(n_514),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_514),
.C(n_508),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_541),
.A2(n_505),
.B1(n_515),
.B2(n_516),
.Y(n_557)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_560),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_531),
.B(n_528),
.C(n_477),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_561),
.B(n_562),
.C(n_542),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_536),
.B(n_528),
.C(n_477),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_534),
.A2(n_520),
.B1(n_506),
.B2(n_522),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_547),
.A2(n_500),
.B(n_506),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_564),
.A2(n_535),
.B(n_487),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_568),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_571),
.B(n_579),
.Y(n_592)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_563),
.Y(n_572)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_572),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_533),
.Y(n_573)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_573),
.Y(n_588)
);

INVxp33_ASAP7_75t_SL g574 ( 
.A(n_558),
.Y(n_574)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_532),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_575),
.B(n_576),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_523),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_566),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_581),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_567),
.B(n_532),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_578),
.B(n_579),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_552),
.B(n_539),
.C(n_526),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_580),
.A2(n_556),
.B(n_561),
.Y(n_591)
);

CKINVDCx14_ASAP7_75t_R g581 ( 
.A(n_565),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_575),
.C(n_578),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_590),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_570),
.B(n_557),
.C(n_555),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_591),
.A2(n_573),
.B(n_569),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_592),
.B(n_584),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_593),
.A2(n_595),
.B(n_599),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_588),
.B(n_555),
.Y(n_594)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_594),
.Y(n_604)
);

INVx11_ASAP7_75t_L g595 ( 
.A(n_591),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_596),
.B(n_598),
.Y(n_603)
);

OA21x2_ASAP7_75t_SL g598 ( 
.A1(n_586),
.A2(n_574),
.B(n_490),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_587),
.B(n_559),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_592),
.B(n_571),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_600),
.A2(n_585),
.B(n_582),
.Y(n_601)
);

AO21x1_ASAP7_75t_L g606 ( 
.A1(n_601),
.A2(n_595),
.B(n_600),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_597),
.A2(n_589),
.B(n_583),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_605),
.A2(n_543),
.B(n_544),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_606),
.A2(n_608),
.B(n_603),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_602),
.B(n_590),
.C(n_594),
.Y(n_607)
);

A2O1A1O1Ixp25_ASAP7_75t_L g610 ( 
.A1(n_607),
.A2(n_604),
.B(n_562),
.C(n_490),
.D(n_528),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_609),
.B(n_610),
.C(n_529),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_435),
.C(n_498),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_612),
.A2(n_429),
.B(n_498),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_613),
.B(n_426),
.Y(n_614)
);


endmodule