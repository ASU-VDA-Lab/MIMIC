module fake_ariane_2001_n_108 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_108);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_108;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_1),
.C(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_24),
.B1(n_33),
.B2(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_53)
);

OR2x6_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_34),
.Y(n_54)
);

OAI221xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_34),
.B1(n_23),
.B2(n_8),
.C(n_9),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_34),
.B1(n_6),
.B2(n_8),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_3),
.B1(n_15),
.B2(n_16),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_44),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_56),
.B(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_52),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_53),
.B1(n_57),
.B2(n_55),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_40),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_52),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_53),
.B(n_51),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_36),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_63),
.B(n_36),
.C(n_46),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_60),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI211xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_46),
.B(n_37),
.C(n_62),
.Y(n_74)
);

AO21x2_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_68),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_64),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_72),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_70),
.B(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_67),
.Y(n_82)
);

AND3x1_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_76),
.C(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_75),
.Y(n_86)
);

AOI222xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_37),
.B1(n_76),
.B2(n_78),
.C1(n_62),
.C2(n_75),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_75),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_81),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

AND3x4_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_37),
.C(n_85),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_88),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_17),
.B(n_42),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NAND4xp25_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.C(n_100),
.D(n_101),
.Y(n_105)
);

AOI211xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_99),
.B(n_62),
.C(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_42),
.B1(n_62),
.B2(n_105),
.C(n_106),
.Y(n_108)
);


endmodule