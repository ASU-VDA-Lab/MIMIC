module real_jpeg_29730_n_18 (n_17, n_8, n_0, n_2, n_297, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_297;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_286;
wire n_215;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_293;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_70;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_0),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_1),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_29),
.B1(n_35),
.B2(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_72),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_42),
.B1(n_44),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_104),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_104),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_104),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_86),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_86),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_6),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_47),
.B(n_51),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_42),
.B1(n_44),
.B2(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_6),
.B(n_49),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_62),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_6),
.B(n_62),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_6),
.B(n_96),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_27),
.B1(n_235),
.B2(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_6),
.A2(n_50),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_42),
.B1(n_44),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_7),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_135),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_135),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_135),
.Y(n_229)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_64),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_41),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_11),
.A2(n_42),
.B1(n_44),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_11),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_11),
.A2(n_29),
.B1(n_35),
.B2(n_54),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_68),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_35),
.A3(n_62),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_17),
.A2(n_42),
.B1(n_44),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_17),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_17),
.A2(n_50),
.B1(n_51),
.B2(n_142),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_142),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_17),
.A2(n_29),
.B1(n_35),
.B2(n_142),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_22),
.B(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.C(n_91),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_23),
.B(n_75),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_56),
.B1(n_57),
.B2(n_74),
.Y(n_23)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_38),
.B(n_56),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_25),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_27),
.A2(n_31),
.B1(n_34),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_27),
.A2(n_33),
.B1(n_99),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_27),
.A2(n_33),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_27),
.A2(n_33),
.B1(n_229),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_27),
.A2(n_224),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_28),
.A2(n_128),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_28),
.A2(n_32),
.B1(n_149),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_28),
.A2(n_32),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_29),
.B(n_68),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_29),
.B(n_241),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_31),
.Y(n_150)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g263 ( 
.A(n_32),
.Y(n_263)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_33),
.B(n_146),
.Y(n_241)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_53),
.B2(n_55),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_42),
.A2(n_52),
.B(n_146),
.C(n_147),
.Y(n_145)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_45),
.A2(n_53),
.B1(n_55),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_45),
.A2(n_55),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_46),
.A2(n_49),
.B1(n_103),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_46),
.A2(n_49),
.B1(n_141),
.B2(n_179),
.Y(n_178)
);

AO22x1_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_78),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_50),
.A2(n_63),
.A3(n_82),
.B1(n_252),
.B2(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_51),
.B(n_146),
.Y(n_252)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_70),
.B2(n_73),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_63),
.B1(n_79),
.B2(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_62),
.B(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_65),
.A2(n_73),
.B1(n_131),
.B2(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_65),
.A2(n_73),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_67),
.B(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_66),
.A2(n_67),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_66),
.A2(n_67),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_66),
.A2(n_67),
.B1(n_210),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_66),
.A2(n_67),
.B1(n_177),
.B2(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_67),
.B(n_146),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_88),
.B(n_90),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_88),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_81),
.B1(n_84),
.B2(n_87),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_77),
.A2(n_81),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_77),
.A2(n_81),
.B1(n_152),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_77),
.A2(n_81),
.B1(n_185),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

FAx1_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_106),
.CI(n_118),
.CON(n_105),
.SN(n_105)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_91),
.A2(n_92),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_102),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_93),
.B(n_97),
.CI(n_102),
.CON(n_158),
.SN(n_158)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_96),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_95),
.A2(n_96),
.B1(n_173),
.B2(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_100),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_105),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_117),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_114),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_160),
.A3(n_165),
.B1(n_288),
.B2(n_293),
.C(n_297),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_122),
.A2(n_289),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_155),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_123),
.B(n_155),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.C(n_154),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_124),
.B(n_154),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_133),
.C(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_129),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_138),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.C(n_151),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_144),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_148),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.C(n_159),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_158),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_161),
.B(n_162),
.Y(n_293)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_195),
.C(n_200),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_189),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_167),
.B(n_189),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_180),
.C(n_181),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_168),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_175),
.C(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_180),
.Y(n_286)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_183),
.B(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_186),
.B(n_188),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_187),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_196),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_197),
.B(n_198),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_282),
.B(n_287),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_268),
.B(n_281),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_245),
.B(n_267),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_225),
.B(n_244),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_215),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_222),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_223),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_243),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_242),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_246),
.B(n_247),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_258),
.B1(n_265),
.B2(n_266),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_257),
.C(n_266),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_258),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_262),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_277),
.C(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);


endmodule