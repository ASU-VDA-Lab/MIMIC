module real_aes_7674_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_1), .A2(n_102), .B1(n_115), .B2(n_727), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_2), .A2(n_145), .B(n_150), .C(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_3), .A2(n_140), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g456 ( .A(n_4), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_5), .B(n_164), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_6), .A2(n_16), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_6), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g473 ( .A1(n_7), .A2(n_140), .B(n_474), .Y(n_473) );
AND2x6_ASAP7_75t_L g145 ( .A(n_8), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g174 ( .A(n_9), .Y(n_174) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_10), .B(n_44), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_11), .A2(n_252), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_12), .B(n_155), .Y(n_191) );
INVx1_ASAP7_75t_L g478 ( .A(n_13), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_14), .B(n_154), .Y(n_526) );
INVx1_ASAP7_75t_L g138 ( .A(n_15), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_16), .Y(n_716) );
INVx1_ASAP7_75t_L g538 ( .A(n_17), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_18), .A2(n_175), .B(n_200), .C(n_202), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_19), .B(n_164), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_20), .B(n_467), .Y(n_517) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_21), .A2(n_444), .B1(n_715), .B2(n_718), .C1(n_721), .C2(n_725), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_22), .B(n_140), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_23), .B(n_260), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_24), .A2(n_154), .B(n_156), .C(n_160), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_25), .B(n_164), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_26), .B(n_155), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_27), .A2(n_158), .B(n_202), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_28), .B(n_155), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_29), .Y(n_220) );
INVx1_ASAP7_75t_L g234 ( .A(n_30), .Y(n_234) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_31), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_32), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_33), .B(n_155), .Y(n_457) );
INVx1_ASAP7_75t_L g257 ( .A(n_34), .Y(n_257) );
INVx1_ASAP7_75t_L g491 ( .A(n_35), .Y(n_491) );
INVx2_ASAP7_75t_L g143 ( .A(n_36), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_37), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_38), .A2(n_154), .B(n_213), .C(n_215), .Y(n_212) );
INVxp67_ASAP7_75t_L g258 ( .A(n_39), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g211 ( .A(n_40), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_41), .A2(n_150), .B(n_233), .C(n_239), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_42), .A2(n_145), .B(n_150), .C(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_43), .A2(n_90), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_43), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_44), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g490 ( .A(n_45), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_46), .A2(n_172), .B(n_173), .C(n_176), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_47), .B(n_155), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_48), .B(n_441), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_49), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_50), .Y(n_254) );
INVx1_ASAP7_75t_L g148 ( .A(n_51), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_52), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_53), .B(n_140), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_54), .A2(n_150), .B1(n_160), .B2(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_55), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_56), .Y(n_453) );
CKINVDCx14_ASAP7_75t_R g170 ( .A(n_57), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_58), .A2(n_172), .B(n_215), .C(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_59), .Y(n_519) );
INVx1_ASAP7_75t_L g475 ( .A(n_60), .Y(n_475) );
INVx1_ASAP7_75t_L g146 ( .A(n_61), .Y(n_146) );
INVx1_ASAP7_75t_L g137 ( .A(n_62), .Y(n_137) );
INVx1_ASAP7_75t_SL g214 ( .A(n_63), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_64), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_65), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g223 ( .A(n_66), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_SL g466 ( .A1(n_67), .A2(n_215), .B(n_467), .C(n_468), .Y(n_466) );
INVxp67_ASAP7_75t_L g469 ( .A(n_68), .Y(n_469) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_70), .A2(n_140), .B(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_71), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_72), .A2(n_140), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_73), .Y(n_494) );
INVx1_ASAP7_75t_L g513 ( .A(n_74), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_75), .A2(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g198 ( .A(n_76), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_77), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_78), .A2(n_145), .B(n_150), .C(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_79), .A2(n_140), .B(n_147), .Y(n_139) );
INVx1_ASAP7_75t_L g201 ( .A(n_80), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_81), .B(n_235), .Y(n_507) );
INVx2_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
INVx1_ASAP7_75t_L g188 ( .A(n_83), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_84), .B(n_467), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_85), .A2(n_145), .B(n_150), .C(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
OR2x2_ASAP7_75t_L g436 ( .A(n_86), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g714 ( .A(n_86), .B(n_438), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_87), .A2(n_150), .B(n_222), .C(n_225), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_88), .B(n_167), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_89), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_90), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_91), .A2(n_145), .B(n_150), .C(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_92), .Y(n_530) );
INVx1_ASAP7_75t_L g465 ( .A(n_93), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_94), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_95), .B(n_235), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_96), .B(n_133), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_97), .B(n_133), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_100), .A2(n_140), .B(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g729 ( .A(n_104), .Y(n_729) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g438 ( .A(n_110), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g713 ( .A(n_111), .B(n_438), .Y(n_713) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_111), .B(n_437), .Y(n_720) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_442), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g726 ( .A(n_118), .Y(n_726) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_433), .B(n_440), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_431), .B2(n_432), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_122), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_125), .A2(n_713), .B1(n_722), .B2(n_723), .Y(n_721) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g432 ( .A(n_126), .Y(n_432) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_357), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_299), .C(n_329), .D(n_339), .Y(n_127) );
OAI211xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_204), .B(n_262), .C(n_289), .Y(n_128) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_129), .A2(n_304), .B1(n_385), .B2(n_386), .C1(n_387), .C2(n_388), .Y(n_384) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_179), .Y(n_129) );
AOI33xp33_ASAP7_75t_L g310 ( .A1(n_130), .A2(n_297), .A3(n_298), .B1(n_311), .B2(n_316), .B3(n_318), .Y(n_310) );
OAI211xp5_ASAP7_75t_SL g367 ( .A1(n_130), .A2(n_368), .B(n_370), .C(n_372), .Y(n_367) );
OR2x2_ASAP7_75t_L g383 ( .A(n_130), .B(n_369), .Y(n_383) );
INVx1_ASAP7_75t_L g416 ( .A(n_130), .Y(n_416) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
INVx2_ASAP7_75t_L g293 ( .A(n_131), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_131), .B(n_195), .Y(n_309) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_131), .Y(n_344) );
AND2x2_ASAP7_75t_L g373 ( .A(n_131), .B(n_166), .Y(n_373) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_163), .Y(n_131) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_132), .A2(n_196), .B(n_203), .Y(n_195) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_132), .A2(n_209), .B(n_217), .Y(n_208) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx4_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_133), .A2(n_463), .B(n_470), .Y(n_462) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g250 ( .A(n_134), .Y(n_250) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_135), .B(n_136), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g252 ( .A(n_140), .Y(n_252) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_141), .B(n_145), .Y(n_185) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g238 ( .A(n_142), .Y(n_238) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx1_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
INVx3_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx1_ASAP7_75t_L g467 ( .A(n_144), .Y(n_467) );
INVx4_ASAP7_75t_SL g162 ( .A(n_145), .Y(n_162) );
BUFx3_ASAP7_75t_L g239 ( .A(n_145), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g147 ( .A1(n_148), .A2(n_149), .B(n_153), .C(n_162), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_149), .A2(n_162), .B(n_170), .C(n_171), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g197 ( .A1(n_149), .A2(n_162), .B(n_198), .C(n_199), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_149), .A2(n_162), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_149), .A2(n_162), .B(n_254), .C(n_255), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_149), .A2(n_162), .B(n_465), .C(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_149), .A2(n_162), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_149), .A2(n_162), .B(n_535), .C(n_536), .Y(n_534) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx3_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_154), .B(n_214), .Y(n_213) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_158), .B(n_201), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_158), .A2(n_235), .B1(n_257), .B2(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_158), .B(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_159), .A2(n_190), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g458 ( .A(n_160), .Y(n_458) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_162), .A2(n_185), .B1(n_488), .B2(n_492), .Y(n_487) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_164), .A2(n_473), .B(n_479), .Y(n_472) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_165), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_219), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_165), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g509 ( .A(n_165), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g273 ( .A(n_166), .Y(n_273) );
BUFx3_ASAP7_75t_L g281 ( .A(n_166), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_166), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g292 ( .A(n_166), .B(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_166), .B(n_180), .Y(n_321) );
AND2x2_ASAP7_75t_L g390 ( .A(n_166), .B(n_324), .Y(n_390) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_178), .Y(n_166) );
INVx1_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
INVx2_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_167), .A2(n_185), .B(n_231), .C(n_232), .Y(n_230) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_167), .A2(n_533), .B(n_539), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
INVx5_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_175), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_175), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
INVx2_ASAP7_75t_SL g284 ( .A(n_179), .Y(n_284) );
OR2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_195), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_180), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g326 ( .A(n_180), .Y(n_326) );
AND2x2_ASAP7_75t_L g337 ( .A(n_180), .B(n_293), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_180), .B(n_322), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_180), .B(n_324), .Y(n_369) );
AND2x2_ASAP7_75t_L g428 ( .A(n_180), .B(n_373), .Y(n_428) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g298 ( .A(n_181), .B(n_195), .Y(n_298) );
AND2x2_ASAP7_75t_L g308 ( .A(n_181), .B(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g330 ( .A(n_181), .Y(n_330) );
AND3x2_ASAP7_75t_L g389 ( .A(n_181), .B(n_390), .C(n_391), .Y(n_389) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_193), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_182), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_182), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_182), .B(n_530), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_185), .A2(n_220), .B(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_185), .A2(n_453), .B(n_454), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_185), .A2(n_513), .B(n_514), .Y(n_512) );
O2A1O1Ixp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .C(n_192), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_192), .B(n_223), .C(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_192), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_192), .A2(n_516), .B(n_517), .Y(n_515) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
INVx1_ASAP7_75t_SL g324 ( .A(n_195), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_195), .B(n_273), .C(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_242), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_205), .A2(n_308), .B(n_360), .C(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_229), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_207), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g376 ( .A(n_207), .Y(n_376) );
AND2x2_ASAP7_75t_L g397 ( .A(n_207), .B(n_244), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_207), .B(n_306), .Y(n_425) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_261), .Y(n_270) );
INVx2_ASAP7_75t_L g277 ( .A(n_208), .Y(n_277) );
AND2x2_ASAP7_75t_L g297 ( .A(n_208), .B(n_244), .Y(n_297) );
AND2x2_ASAP7_75t_L g347 ( .A(n_208), .B(n_229), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_208), .Y(n_351) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_216), .Y(n_527) );
INVx2_ASAP7_75t_SL g261 ( .A(n_218), .Y(n_261) );
BUFx2_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
AND2x2_ASAP7_75t_L g414 ( .A(n_218), .B(n_229), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_228), .A2(n_522), .B(n_529), .Y(n_521) );
INVx3_ASAP7_75t_SL g244 ( .A(n_229), .Y(n_244) );
AND2x2_ASAP7_75t_L g269 ( .A(n_229), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g276 ( .A(n_229), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g306 ( .A(n_229), .B(n_266), .Y(n_306) );
OR2x2_ASAP7_75t_L g315 ( .A(n_229), .B(n_261), .Y(n_315) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_229), .Y(n_333) );
AND2x2_ASAP7_75t_L g338 ( .A(n_229), .B(n_291), .Y(n_338) );
AND2x2_ASAP7_75t_L g366 ( .A(n_229), .B(n_246), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_229), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_229), .B(n_245), .Y(n_404) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_240), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .C(n_237), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_235), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_238), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g328 ( .A(n_244), .B(n_277), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_244), .B(n_270), .Y(n_356) );
AND2x2_ASAP7_75t_L g374 ( .A(n_244), .B(n_291), .Y(n_374) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_261), .Y(n_245) );
AND2x2_ASAP7_75t_L g275 ( .A(n_246), .B(n_261), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_246), .B(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
OR2x2_ASAP7_75t_L g361 ( .A(n_246), .B(n_281), .Y(n_361) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_251), .B(n_259), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_248), .A2(n_267), .B(n_268), .Y(n_266) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_248), .A2(n_512), .B(n_518), .Y(n_511) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_SL g503 ( .A1(n_249), .A2(n_504), .B(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_250), .A2(n_452), .B(n_459), .Y(n_451) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_250), .A2(n_487), .B(n_493), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_250), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_259), .Y(n_268) );
AND2x2_ASAP7_75t_L g296 ( .A(n_261), .B(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g304 ( .A(n_261), .Y(n_304) );
AND2x2_ASAP7_75t_L g399 ( .A(n_261), .B(n_277), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_271), .B1(n_274), .B2(n_278), .C1(n_282), .C2(n_285), .Y(n_262) );
INVx1_ASAP7_75t_L g394 ( .A(n_263), .Y(n_394) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_269), .Y(n_263) );
AND2x2_ASAP7_75t_L g290 ( .A(n_264), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g301 ( .A(n_264), .B(n_270), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_264), .B(n_292), .Y(n_317) );
OAI222xp33_ASAP7_75t_L g339 ( .A1(n_264), .A2(n_340), .B1(n_345), .B2(n_346), .C1(n_354), .C2(n_356), .Y(n_339) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g327 ( .A(n_266), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_266), .B(n_347), .Y(n_387) );
AND2x2_ASAP7_75t_L g398 ( .A(n_266), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g406 ( .A(n_269), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_271), .B(n_322), .Y(n_385) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_273), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g343 ( .A(n_273), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx3_ASAP7_75t_L g288 ( .A(n_276), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_276), .A2(n_379), .B(n_382), .C(n_384), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_276), .B(n_313), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_276), .B(n_296), .Y(n_418) );
AND2x2_ASAP7_75t_L g291 ( .A(n_277), .B(n_287), .Y(n_291) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_281), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g370 ( .A(n_281), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g409 ( .A(n_281), .B(n_309), .Y(n_409) );
INVx1_ASAP7_75t_L g421 ( .A(n_281), .Y(n_421) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_284), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g402 ( .A(n_287), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .B(n_294), .C(n_298), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_290), .A2(n_320), .B1(n_335), .B2(n_338), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_291), .B(n_305), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_291), .B(n_313), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_292), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g355 ( .A(n_292), .Y(n_355) );
AND2x2_ASAP7_75t_L g362 ( .A(n_292), .B(n_342), .Y(n_362) );
INVx2_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NOR4xp25_ASAP7_75t_L g300 ( .A(n_297), .B(n_301), .C(n_302), .D(n_305), .Y(n_300) );
INVx1_ASAP7_75t_SL g371 ( .A(n_298), .Y(n_371) );
AND2x2_ASAP7_75t_L g415 ( .A(n_298), .B(n_416), .Y(n_415) );
OAI211xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_307), .B(n_310), .C(n_319), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_306), .B(n_376), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_308), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_426) );
INVx1_ASAP7_75t_SL g381 ( .A(n_309), .Y(n_381) );
AND2x2_ASAP7_75t_L g420 ( .A(n_309), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_313), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_317), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_318), .B(n_343), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_325), .B(n_327), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g395 ( .A(n_322), .Y(n_395) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g423 ( .A(n_323), .Y(n_423) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B(n_334), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_330), .Y(n_342) );
OR2x2_ASAP7_75t_L g380 ( .A(n_330), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_333), .A2(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_337), .A2(n_364), .B1(n_367), .B2(n_374), .C(n_375), .Y(n_363) );
INVx1_ASAP7_75t_SL g407 ( .A(n_338), .Y(n_407) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OR2x2_ASAP7_75t_L g354 ( .A(n_342), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_351), .B2(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_350), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_392), .C(n_405), .D(n_417), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g358 ( .A(n_359), .B(n_363), .C(n_378), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_361), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_368), .B(n_373), .Y(n_377) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g405 ( .A1(n_380), .A2(n_406), .B1(n_407), .B2(n_408), .C(n_410), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_382), .A2(n_397), .B(n_398), .C(n_400), .Y(n_396) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_383), .A2(n_401), .B1(n_403), .B2(n_404), .Y(n_400) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B(n_395), .C(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g411 ( .A(n_404), .Y(n_411) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI221xp5_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_432), .A2(n_445), .B1(n_713), .B2(n_714), .Y(n_444) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g441 ( .A(n_436), .Y(n_441) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_440), .A2(n_443), .B(n_726), .Y(n_442) );
INVx1_ASAP7_75t_L g722 ( .A(n_445), .Y(n_722) );
NAND2x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_629), .Y(n_445) );
NOR5xp2_ASAP7_75t_L g446 ( .A(n_447), .B(n_552), .C(n_584), .D(n_599), .E(n_616), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_480), .B(n_499), .C(n_540), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_461), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_449), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_449), .B(n_604), .Y(n_667) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_450), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_450), .B(n_496), .Y(n_553) );
AND2x2_ASAP7_75t_L g594 ( .A(n_450), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_450), .B(n_563), .Y(n_598) );
OR2x2_ASAP7_75t_L g635 ( .A(n_450), .B(n_486), .Y(n_635) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g485 ( .A(n_451), .B(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g543 ( .A(n_451), .Y(n_543) );
OR2x2_ASAP7_75t_L g706 ( .A(n_451), .B(n_546), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_461), .A2(n_609), .B1(n_610), .B2(n_613), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_461), .B(n_543), .Y(n_692) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_471), .Y(n_461) );
AND2x2_ASAP7_75t_L g498 ( .A(n_462), .B(n_486), .Y(n_498) );
AND2x2_ASAP7_75t_L g545 ( .A(n_462), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g550 ( .A(n_462), .Y(n_550) );
INVx3_ASAP7_75t_L g563 ( .A(n_462), .Y(n_563) );
OR2x2_ASAP7_75t_L g583 ( .A(n_462), .B(n_546), .Y(n_583) );
AND2x2_ASAP7_75t_L g602 ( .A(n_462), .B(n_472), .Y(n_602) );
BUFx2_ASAP7_75t_L g634 ( .A(n_462), .Y(n_634) );
AND2x4_ASAP7_75t_L g549 ( .A(n_471), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g484 ( .A(n_472), .Y(n_484) );
INVx2_ASAP7_75t_L g497 ( .A(n_472), .Y(n_497) );
OR2x2_ASAP7_75t_L g565 ( .A(n_472), .B(n_546), .Y(n_565) );
AND2x2_ASAP7_75t_L g595 ( .A(n_472), .B(n_486), .Y(n_595) );
AND2x2_ASAP7_75t_L g612 ( .A(n_472), .B(n_543), .Y(n_612) );
AND2x2_ASAP7_75t_L g652 ( .A(n_472), .B(n_563), .Y(n_652) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_472), .B(n_498), .Y(n_688) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp33_ASAP7_75t_SL g481 ( .A(n_482), .B(n_495), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_483), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
OAI21xp33_ASAP7_75t_L g626 ( .A1(n_484), .A2(n_498), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_484), .B(n_486), .Y(n_682) );
AND2x2_ASAP7_75t_L g618 ( .A(n_485), .B(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g546 ( .A(n_486), .Y(n_546) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_486), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_495), .B(n_543), .Y(n_711) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_496), .A2(n_654), .B1(n_655), .B2(n_660), .Y(n_653) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x2_ASAP7_75t_L g544 ( .A(n_497), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g582 ( .A(n_497), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g619 ( .A(n_497), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_498), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g673 ( .A(n_498), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_520), .Y(n_500) );
INVx4_ASAP7_75t_L g559 ( .A(n_501), .Y(n_559) );
AND2x2_ASAP7_75t_L g637 ( .A(n_501), .B(n_604), .Y(n_637) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
INVx3_ASAP7_75t_L g556 ( .A(n_502), .Y(n_556) );
AND2x2_ASAP7_75t_L g570 ( .A(n_502), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g574 ( .A(n_502), .Y(n_574) );
INVx2_ASAP7_75t_L g588 ( .A(n_502), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_502), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g645 ( .A(n_502), .B(n_640), .Y(n_645) );
AND2x2_ASAP7_75t_L g710 ( .A(n_502), .B(n_680), .Y(n_710) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
AND2x2_ASAP7_75t_L g551 ( .A(n_511), .B(n_532), .Y(n_551) );
INVx2_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
INVx1_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
AND2x2_ASAP7_75t_L g622 ( .A(n_520), .B(n_570), .Y(n_622) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
INVx2_ASAP7_75t_L g561 ( .A(n_521), .Y(n_561) );
INVx1_ASAP7_75t_L g569 ( .A(n_521), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_521), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_521), .B(n_571), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_527), .Y(n_524) );
AND2x2_ASAP7_75t_L g604 ( .A(n_531), .B(n_561), .Y(n_604) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g557 ( .A(n_532), .Y(n_557) );
AND2x2_ASAP7_75t_L g640 ( .A(n_532), .B(n_571), .Y(n_640) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_547), .B(n_551), .Y(n_540) );
INVx1_ASAP7_75t_SL g585 ( .A(n_541), .Y(n_585) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_542), .B(n_549), .Y(n_642) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g591 ( .A(n_543), .B(n_546), .Y(n_591) );
AND2x2_ASAP7_75t_L g620 ( .A(n_543), .B(n_564), .Y(n_620) );
OR2x2_ASAP7_75t_L g623 ( .A(n_543), .B(n_583), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_544), .A2(n_636), .B1(n_688), .B2(n_689), .C1(n_691), .C2(n_693), .Y(n_687) );
BUFx2_ASAP7_75t_L g601 ( .A(n_546), .Y(n_601) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g590 ( .A(n_549), .B(n_591), .Y(n_590) );
INVx3_ASAP7_75t_SL g607 ( .A(n_549), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_549), .B(n_601), .Y(n_661) );
AND2x2_ASAP7_75t_L g596 ( .A(n_551), .B(n_556), .Y(n_596) );
INVx1_ASAP7_75t_L g615 ( .A(n_551), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_554), .B1(n_558), .B2(n_562), .C(n_566), .Y(n_552) );
OR2x2_ASAP7_75t_L g624 ( .A(n_554), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g609 ( .A(n_556), .B(n_579), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_556), .B(n_569), .Y(n_649) );
AND2x2_ASAP7_75t_L g654 ( .A(n_556), .B(n_604), .Y(n_654) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_556), .Y(n_664) );
NAND2x1_ASAP7_75t_SL g675 ( .A(n_556), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g560 ( .A(n_557), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g580 ( .A(n_557), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_557), .B(n_575), .Y(n_606) );
INVx1_ASAP7_75t_L g672 ( .A(n_557), .Y(n_672) );
INVx1_ASAP7_75t_L g647 ( .A(n_558), .Y(n_647) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g659 ( .A(n_559), .Y(n_659) );
NOR2xp67_ASAP7_75t_L g671 ( .A(n_559), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g676 ( .A(n_560), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_560), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g579 ( .A(n_561), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_561), .B(n_571), .Y(n_592) );
INVx1_ASAP7_75t_L g658 ( .A(n_561), .Y(n_658) );
INVx1_ASAP7_75t_L g679 ( .A(n_562), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI21xp5_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_572), .B(n_581), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
AND2x2_ASAP7_75t_L g712 ( .A(n_568), .B(n_645), .Y(n_712) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g680 ( .A(n_569), .B(n_640), .Y(n_680) );
AOI32xp33_ASAP7_75t_L g593 ( .A1(n_570), .A2(n_576), .A3(n_594), .B1(n_596), .B2(n_597), .Y(n_593) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_570), .A2(n_602), .A3(n_685), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_700), .Y(n_695) );
INVx2_ASAP7_75t_L g575 ( .A(n_571), .Y(n_575) );
INVx1_ASAP7_75t_L g685 ( .A(n_571), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_573), .B(n_579), .Y(n_628) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_574), .B(n_640), .Y(n_690) );
INVx1_ASAP7_75t_L g577 ( .A(n_575), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_575), .B(n_604), .Y(n_694) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_583), .B(n_678), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_586), .B1(n_589), .B2(n_592), .C(n_593), .Y(n_584) );
OR2x2_ASAP7_75t_L g605 ( .A(n_586), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g614 ( .A(n_586), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g639 ( .A(n_587), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g643 ( .A(n_597), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_605), .B2(n_607), .C(n_608), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_601), .A2(n_632), .B1(n_636), .B2(n_637), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_602), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_602), .Y(n_707) );
INVx1_ASAP7_75t_L g701 ( .A(n_604), .Y(n_701) );
INVx1_ASAP7_75t_SL g636 ( .A(n_605), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_607), .B(n_635), .Y(n_697) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_612), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g678 ( .A(n_612), .Y(n_678) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_621), .B1(n_623), .B2(n_624), .C(n_626), .Y(n_616) );
NOR2xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_620), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_618), .A2(n_636), .B1(n_682), .B2(n_683), .Y(n_681) );
CKINVDCx14_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_623), .A2(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR3xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_662), .C(n_686), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_631), .B(n_638), .C(n_646), .D(n_653), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g709 ( .A(n_634), .Y(n_709) );
INVx3_ASAP7_75t_SL g703 ( .A(n_635), .Y(n_703) );
OR2x2_ASAP7_75t_L g708 ( .A(n_635), .B(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_643), .B2(n_645), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_640), .B(n_658), .Y(n_699) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_648), .B(n_650), .Y(n_646) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_665), .B(n_668), .C(n_681), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g696 ( .A(n_667), .Y(n_696) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_673), .B1(n_674), .B2(n_677), .C1(n_679), .C2(n_680), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND4xp25_ASAP7_75t_SL g705 ( .A(n_678), .B(n_706), .C(n_707), .D(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_695), .C(n_704), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_704) );
INVx1_ASAP7_75t_L g724 ( .A(n_714), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_715), .Y(n_725) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx3_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
endmodule