module real_jpeg_27648_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_249;
wire n_292;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_299;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_0),
.B(n_52),
.Y(n_84)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_0),
.B(n_230),
.Y(n_235)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_30),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_30),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_44),
.B1(n_48),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_50),
.B1(n_52),
.B2(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_1),
.B(n_21),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_1),
.A2(n_10),
.B(n_44),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_1),
.A2(n_47),
.B(n_50),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_1),
.B(n_64),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_44),
.B1(n_48),
.B2(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_5),
.B1(n_30),
.B2(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_50),
.B1(n_52),
.B2(n_67),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_5),
.A2(n_7),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_6),
.B1(n_30),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_136),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_44),
.B1(n_48),
.B2(n_136),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_50),
.B1(n_52),
.B2(n_136),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_31),
.B1(n_44),
.B2(n_48),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_7),
.A2(n_31),
.B1(n_50),
.B2(n_52),
.Y(n_122)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_11),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_16),
.B(n_92),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_71),
.C(n_79),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_17),
.B(n_71),
.CI(n_79),
.CON(n_142),
.SN(n_142)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_38),
.B2(n_39),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_18),
.A2(n_19),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_57),
.C(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_20),
.B(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_21),
.B(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_23),
.B(n_30),
.C(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_22),
.A2(n_34),
.B(n_36),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_22),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_22),
.B(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_27),
.Y(n_172)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_25),
.A2(n_59),
.B(n_60),
.C(n_64),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_25),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_25),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_25),
.A2(n_56),
.B(n_59),
.C(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_34),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_33),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_34),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_35),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_36),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_37),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_57),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_40),
.A2(n_109),
.B1(n_158),
.B2(n_159),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_53),
.B(n_54),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_41),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_42),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_42),
.B(n_55),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_42),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_44),
.A2(n_46),
.B(n_56),
.C(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_49),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_52),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_77),
.B(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_53),
.B(n_56),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_56),
.B(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_65),
.B(n_68),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_58),
.B(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_58),
.B(n_161),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_58),
.Y(n_277)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_64),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_169),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_73),
.A2(n_104),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_74),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_76),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_77),
.B(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_81),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_82),
.A2(n_83),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_83),
.B(n_195),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_84),
.B(n_87),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_84),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_85),
.B(n_122),
.Y(n_152)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_88),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_90),
.B(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_91),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_107),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_99),
.B(n_157),
.Y(n_274)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_103),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_156),
.C(n_158),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_143),
.B(n_300),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_142),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_113),
.B(n_142),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_137),
.C(n_138),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_114),
.A2(n_115),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_125),
.C(n_128),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_116),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_117),
.B(n_124),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_118),
.B(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_119),
.A2(n_151),
.B(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_120),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_160),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_137),
.B(n_138),
.Y(n_298)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_142),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_294),
.B(n_299),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_281),
.B(n_293),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_189),
.B(n_264),
.C(n_280),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_177),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_147),
.B(n_177),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_162),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_149),
.B(n_155),
.C(n_162),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_150),
.B(n_153),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_152),
.B(n_229),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_154),
.B(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_170),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_164),
.B(n_167),
.C(n_170),
.Y(n_278)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_178),
.A2(n_179),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_263),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_256),
.B(n_262),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_214),
.B(n_255),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_204),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_193),
.B(n_204),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.C(n_200),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_194),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_211),
.C(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_250),
.B(n_254),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_231),
.B(n_249),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_238),
.B(n_248),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_242),
.B(n_247),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_266),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_278),
.B2(n_279),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_270),
.C(n_279),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_274),
.C(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_289),
.B2(n_290),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_290),
.C(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);


endmodule