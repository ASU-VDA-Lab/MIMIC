module fake_jpeg_31991_n_403 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_403);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_403;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_57),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_25),
.B1(n_41),
.B2(n_35),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_15),
.B(n_0),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_73),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_3),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_16),
.B(n_3),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_76),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_19),
.B(n_3),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_85),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_39),
.B1(n_23),
.B2(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_23),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_89),
.A2(n_93),
.B1(n_99),
.B2(n_110),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_42),
.B1(n_39),
.B2(n_30),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_42),
.B1(n_39),
.B2(n_32),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_34),
.B(n_41),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_47),
.B(n_82),
.C(n_22),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_103),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_34),
.B1(n_35),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_104),
.A2(n_114),
.B1(n_119),
.B2(n_120),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_112),
.A2(n_118),
.B1(n_22),
.B2(n_28),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_25),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_115),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_76),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_48),
.A2(n_22),
.B1(n_28),
.B2(n_11),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_62),
.B1(n_53),
.B2(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_52),
.B(n_8),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_8),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_57),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_151),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_134),
.Y(n_143)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_46),
.B1(n_44),
.B2(n_59),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_65),
.B1(n_50),
.B2(n_66),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_149),
.A2(n_159),
.B1(n_161),
.B2(n_169),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_56),
.C(n_69),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_150),
.B(n_164),
.C(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_64),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_28),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_152),
.B(n_160),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_174),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_90),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_60),
.B1(n_71),
.B2(n_68),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_87),
.C(n_85),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_28),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_47),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_171),
.Y(n_222)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_88),
.A2(n_54),
.B1(n_86),
.B2(n_84),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_22),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_74),
.B(n_80),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_123),
.A2(n_22),
.B1(n_28),
.B2(n_12),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_183),
.B1(n_91),
.B2(n_127),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_88),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_127),
.B1(n_102),
.B2(n_107),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_12),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_179),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_10),
.Y(n_178)
);

NOR2x1p5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_105),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_92),
.B(n_100),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_11),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_12),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_121),
.A2(n_124),
.B1(n_94),
.B2(n_108),
.Y(n_183)
);

BUFx4f_ASAP7_75t_SL g184 ( 
.A(n_105),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_97),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_137),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_215),
.B1(n_167),
.B2(n_178),
.C(n_152),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_193),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_168),
.B1(n_163),
.B2(n_158),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_167),
.A2(n_137),
.B1(n_124),
.B2(n_108),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_212),
.B(n_156),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_140),
.B(n_136),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_153),
.A2(n_97),
.B(n_105),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_173),
.C(n_164),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_159),
.B1(n_146),
.B2(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_225),
.B(n_228),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_227),
.A2(n_248),
.B(n_187),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_170),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_231),
.B1(n_188),
.B2(n_191),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_150),
.B1(n_142),
.B2(n_172),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_171),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_233),
.B(n_234),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_166),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_140),
.C(n_179),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_240),
.C(n_246),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_195),
.B1(n_189),
.B2(n_204),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_180),
.C(n_162),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_181),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_184),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_247),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_91),
.C(n_156),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_192),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_184),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_255),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_184),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_205),
.C(n_223),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_188),
.A2(n_143),
.B(n_158),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_201),
.B(n_204),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_143),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_260),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_215),
.B1(n_203),
.B2(n_206),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_266),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_206),
.B1(n_217),
.B2(n_200),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_271),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_251),
.B(n_227),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_213),
.B1(n_208),
.B2(n_187),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_272),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_284),
.C(n_240),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_251),
.A2(n_201),
.B(n_209),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_283),
.B(n_285),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_250),
.B(n_248),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_245),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_239),
.A2(n_205),
.B(n_195),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_239),
.A2(n_224),
.B(n_219),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_255),
.C(n_236),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_270),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_269),
.C(n_274),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_259),
.B(n_236),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_252),
.B(n_256),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_269),
.B(n_280),
.Y(n_313)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_242),
.B(n_234),
.C(n_232),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_273),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_266),
.B(n_231),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_267),
.B(n_278),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_228),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_233),
.Y(n_302)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_235),
.Y(n_306)
);

NOR4xp25_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_244),
.C(n_225),
.D(n_246),
.Y(n_308)
);

OAI322xp33_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_258),
.A3(n_271),
.B1(n_260),
.B2(n_278),
.C1(n_273),
.C2(n_281),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_263),
.A2(n_229),
.B1(n_257),
.B2(n_190),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_312),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_319),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_330),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_326),
.C(n_332),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_329),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_279),
.C(n_261),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_327),
.A2(n_304),
.B(n_296),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_295),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_295),
.C(n_291),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_325),
.A2(n_307),
.B(n_295),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_346),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_307),
.C(n_291),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_343),
.C(n_314),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_325),
.A2(n_311),
.B1(n_310),
.B2(n_309),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_342),
.A2(n_344),
.B1(n_349),
.B2(n_350),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_326),
.C(n_329),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_297),
.B1(n_299),
.B2(n_294),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_301),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_297),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_331),
.Y(n_357)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_318),
.A2(n_290),
.B1(n_289),
.B2(n_264),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_322),
.A2(n_290),
.B1(n_288),
.B2(n_308),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_322),
.A2(n_288),
.B1(n_264),
.B2(n_276),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_351),
.A2(n_323),
.B1(n_330),
.B2(n_276),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_352),
.B(n_357),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_331),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_359),
.C(n_364),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_321),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_361),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_339),
.Y(n_358)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_358),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_321),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_323),
.B1(n_333),
.B2(n_315),
.Y(n_360)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_335),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_334),
.B1(n_243),
.B2(n_257),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_245),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_345),
.A2(n_351),
.B1(n_341),
.B2(n_338),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_340),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_336),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_371),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_354),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_375),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_335),
.B(n_337),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_355),
.B(n_337),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_359),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_364),
.C(n_353),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_385),
.C(n_367),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_379),
.A2(n_380),
.B(n_383),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_357),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_334),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_224),
.B1(n_218),
.B2(n_194),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_384),
.A2(n_199),
.B1(n_158),
.B2(n_111),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_194),
.C(n_190),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_389),
.Y(n_393)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_388),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_366),
.C(n_199),
.Y(n_389)
);

AOI322xp5_ASAP7_75t_L g395 ( 
.A1(n_390),
.A2(n_392),
.A3(n_186),
.B1(n_135),
.B2(n_102),
.C1(n_131),
.C2(n_129),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_369),
.B(n_107),
.Y(n_391)
);

AOI31xp67_ASAP7_75t_SL g394 ( 
.A1(n_391),
.A2(n_186),
.A3(n_385),
.B(n_144),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_381),
.A2(n_144),
.B1(n_129),
.B2(n_131),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_395),
.A3(n_111),
.B1(n_139),
.B2(n_145),
.C1(n_186),
.C2(n_184),
.Y(n_399)
);

AOI322xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_387),
.A3(n_389),
.B1(n_392),
.B2(n_377),
.C1(n_386),
.C2(n_135),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_398),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g398 ( 
.A(n_393),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_399),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_139),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_401),
.Y(n_403)
);


endmodule