module fake_jpeg_15267_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx8_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_17),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_54),
.B1(n_58),
.B2(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_80),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_5),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_47),
.B1(n_57),
.B2(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_47),
.B1(n_46),
.B2(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_46),
.B1(n_44),
.B2(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_78),
.B1(n_79),
.B2(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_15),
.C(n_38),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_5),
.C(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_13),
.B1(n_36),
.B2(n_31),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_87),
.B1(n_93),
.B2(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_90),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_2),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_7),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_16),
.B1(n_29),
.B2(n_27),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_39),
.B1(n_25),
.B2(n_22),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_106),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_103),
.B(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_99),
.B1(n_87),
.B2(n_93),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_85),
.C(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_115),
.B1(n_116),
.B2(n_103),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_112),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_120),
.B1(n_128),
.B2(n_127),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_126),
.C(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_113),
.B1(n_105),
.B2(n_114),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_91),
.CI(n_18),
.CON(n_134),
.SN(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_21),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_20),
.A3(n_134),
.B1(n_109),
.B2(n_83),
.C1(n_8),
.C2(n_11),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_9),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_10),
.B(n_12),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_10),
.Y(n_139)
);


endmodule