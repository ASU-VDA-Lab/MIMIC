module fake_jpeg_27264_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_40),
.Y(n_95)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_40),
.Y(n_79)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_115)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_35),
.B1(n_18),
.B2(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_42),
.B1(n_62),
.B2(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_81),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_96),
.Y(n_99)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_24),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx9p33_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_95),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_86),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_123),
.B1(n_85),
.B2(n_60),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_35),
.B1(n_18),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_127),
.B1(n_20),
.B2(n_25),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_120),
.B1(n_52),
.B2(n_69),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_124),
.Y(n_130)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_48),
.B1(n_47),
.B2(n_39),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_80),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_45),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_82),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_46),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_153),
.C(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_94),
.B1(n_91),
.B2(n_59),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_139),
.B1(n_149),
.B2(n_152),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_135),
.Y(n_163)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_151),
.Y(n_156)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_126),
.B1(n_99),
.B2(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_68),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_68),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_146),
.Y(n_179)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_110),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_20),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_66),
.B1(n_73),
.B2(n_88),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_38),
.B(n_27),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_31),
.B(n_28),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_88),
.B1(n_73),
.B2(n_52),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_44),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_44),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_120),
.C(n_111),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_44),
.C(n_45),
.Y(n_154)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_162),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_124),
.B1(n_102),
.B2(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_182),
.B1(n_164),
.B2(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_167),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_106),
.C(n_103),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_133),
.C(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_172),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_173),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_102),
.B1(n_101),
.B2(n_106),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_176),
.B1(n_183),
.B2(n_155),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_101),
.B1(n_103),
.B2(n_25),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_110),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_36),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_125),
.B1(n_45),
.B2(n_44),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_125),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_32),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_45),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_69),
.B(n_30),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_153),
.B1(n_154),
.B2(n_148),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_199),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_148),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_194),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_210),
.B1(n_215),
.B2(n_2),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_1),
.C(n_2),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_133),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_203),
.Y(n_223)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_133),
.C(n_141),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_207),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_184),
.B(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_159),
.B(n_30),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_209),
.B(n_211),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_164),
.A2(n_161),
.B1(n_157),
.B2(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_178),
.B(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_214),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_32),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_162),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_21),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_218),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_32),
.C(n_19),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_221),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_232),
.B(n_200),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_165),
.B1(n_186),
.B2(n_169),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_240),
.B1(n_215),
.B2(n_190),
.Y(n_260)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_239),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_169),
.B1(n_3),
.B2(n_4),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_193),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_191),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_198),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_6),
.Y(n_284)
);

BUFx12_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_203),
.C(n_194),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_258),
.C(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_200),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_210),
.C(n_208),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_231),
.B1(n_230),
.B2(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_210),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_3),
.C(n_4),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_219),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_223),
.B(n_244),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_270),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_243),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_224),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_264),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_235),
.C(n_238),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_281),
.C(n_255),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_249),
.B1(n_262),
.B2(n_263),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_231),
.B1(n_222),
.B2(n_230),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_234),
.C(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_6),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_299),
.C(n_277),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_246),
.B1(n_262),
.B2(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_298),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_255),
.B(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_253),
.C(n_7),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_300),
.C(n_10),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_253),
.B1(n_7),
.B2(n_8),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_275),
.B1(n_11),
.B2(n_12),
.Y(n_307)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_6),
.C(n_7),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_296),
.B(n_291),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_270),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_275),
.B1(n_269),
.B2(n_274),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_293),
.C(n_287),
.Y(n_321)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_272),
.C(n_11),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_300),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_313),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_288),
.B(n_10),
.CI(n_13),
.CON(n_313),
.SN(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_285),
.B(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_321),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_292),
.C(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_314),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_13),
.B(n_14),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_313),
.B(n_320),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_310),
.Y(n_323)
);

OAI221xp5_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_305),
.B1(n_303),
.B2(n_319),
.C(n_14),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_327),
.B(n_328),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_311),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_304),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_302),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_330),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

OAI211xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_15),
.B(n_319),
.C(n_337),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_15),
.Y(n_340)
);


endmodule