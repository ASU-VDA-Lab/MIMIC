module fake_jpeg_2959_n_710 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_710);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_710;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_540;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_544;
wire n_455;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_650;
wire n_344;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_65),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_68),
.B(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_70),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_9),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_76),
.A2(n_77),
.B(n_83),
.C(n_113),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_19),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_78),
.Y(n_213)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_80),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_81),
.Y(n_204)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_85),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_89),
.Y(n_218)
);

BUFx12f_ASAP7_75t_SL g90 ( 
.A(n_20),
.Y(n_90)
);

NAND2x1_ASAP7_75t_SL g177 ( 
.A(n_90),
.B(n_57),
.Y(n_177)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_94),
.Y(n_192)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_103),
.Y(n_165)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_106),
.Y(n_217)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_22),
.B(n_19),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_26),
.Y(n_118)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_29),
.Y(n_125)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_25),
.Y(n_126)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_18),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_27),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_29),
.Y(n_128)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_77),
.B(n_49),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_133),
.B(n_152),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_37),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_136),
.B(n_155),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_42),
.B1(n_57),
.B2(n_34),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_139),
.A2(n_144),
.B1(n_186),
.B2(n_193),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_41),
.B1(n_22),
.B2(n_28),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_73),
.A2(n_48),
.B1(n_59),
.B2(n_42),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_149),
.B(n_0),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_68),
.B(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_46),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_81),
.B(n_46),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_157),
.B(n_176),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_116),
.C(n_128),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_167),
.B(n_211),
.C(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_118),
.B(n_28),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_170),
.B(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_43),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_177),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_102),
.B(n_49),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_125),
.A2(n_57),
.B1(n_34),
.B2(n_42),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_72),
.A2(n_48),
.B1(n_57),
.B2(n_42),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_122),
.B(n_33),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_194),
.B(n_40),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_66),
.A2(n_34),
.B1(n_41),
.B2(n_33),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_229),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_69),
.A2(n_34),
.B1(n_37),
.B2(n_43),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_71),
.A2(n_25),
.B1(n_54),
.B2(n_24),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_206),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_121),
.B(n_55),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_214),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_SL g211 ( 
.A1(n_129),
.A2(n_55),
.B(n_54),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_131),
.B(n_55),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_80),
.B(n_54),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_89),
.Y(n_222)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_222),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_224),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_96),
.A2(n_112),
.B1(n_109),
.B2(n_105),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_99),
.A2(n_48),
.B1(n_35),
.B2(n_24),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_231),
.B1(n_193),
.B2(n_144),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_103),
.A2(n_35),
.B1(n_24),
.B2(n_27),
.Y(n_231)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_234),
.B(n_252),
.Y(n_356)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_235),
.Y(n_344)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_35),
.B1(n_40),
.B2(n_27),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_238),
.A2(n_276),
.B1(n_196),
.B2(n_184),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_204),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_146),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_243),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_244),
.B(n_290),
.Y(n_347)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_248),
.Y(n_366)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_250),
.Y(n_353)
);

BUFx16f_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx13_ASAP7_75t_L g342 ( 
.A(n_251),
.Y(n_342)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_135),
.Y(n_253)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_253),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_146),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_265),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_198),
.B(n_40),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_280),
.Y(n_328)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_154),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_137),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_260),
.Y(n_332)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_164),
.Y(n_261)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_261),
.Y(n_376)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_150),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_262),
.Y(n_330)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_141),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_263),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_264),
.B(n_292),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_161),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_161),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_293),
.Y(n_327)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_267),
.Y(n_372)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_148),
.A2(n_51),
.B1(n_18),
.B2(n_15),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_278),
.B1(n_279),
.B2(n_282),
.Y(n_322)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_147),
.A2(n_51),
.B1(n_14),
.B2(n_13),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_140),
.A2(n_190),
.B1(n_204),
.B2(n_175),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_175),
.A2(n_51),
.B1(n_14),
.B2(n_13),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_178),
.B(n_172),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_220),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_281),
.Y(n_341)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_166),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_168),
.Y(n_283)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_283),
.Y(n_363)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_182),
.Y(n_284)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_156),
.B(n_0),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_286),
.B(n_307),
.Y(n_355)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_287),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_295),
.B1(n_301),
.B2(n_310),
.Y(n_338)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_168),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_202),
.A2(n_51),
.B1(n_2),
.B2(n_3),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_296),
.B1(n_300),
.B2(n_302),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_181),
.B(n_14),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_224),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_210),
.B(n_14),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_298),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_210),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_230),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_189),
.Y(n_297)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_192),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_142),
.B(n_10),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_304),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_145),
.A2(n_11),
.B1(n_10),
.B2(n_4),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_195),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_151),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_153),
.B(n_1),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_162),
.C(n_171),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_138),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_201),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_306),
.Y(n_350)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_166),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_183),
.B(n_1),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_134),
.B(n_1),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_213),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_311),
.A2(n_315),
.B1(n_134),
.B2(n_197),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_191),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_313),
.Y(n_359)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_165),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_138),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_314),
.B(n_197),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_213),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g319 ( 
.A1(n_289),
.A2(n_212),
.B1(n_216),
.B2(n_160),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_319),
.A2(n_357),
.B1(n_358),
.B2(n_362),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_271),
.A2(n_165),
.B1(n_226),
.B2(n_205),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_339),
.A2(n_232),
.B1(n_295),
.B2(n_304),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_345),
.B(n_361),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_259),
.A2(n_205),
.B1(n_226),
.B2(n_159),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_351),
.A2(n_232),
.B1(n_313),
.B2(n_276),
.Y(n_384)
);

AOI22x1_ASAP7_75t_SL g352 ( 
.A1(n_257),
.A2(n_195),
.B1(n_225),
.B2(n_218),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_352),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_252),
.A2(n_160),
.B1(n_158),
.B2(n_218),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_246),
.A2(n_158),
.B1(n_225),
.B2(n_215),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_244),
.A2(n_197),
.B1(n_196),
.B2(n_184),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_360),
.A2(n_264),
.B1(n_282),
.B2(n_291),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_247),
.A2(n_215),
.B1(n_173),
.B2(n_209),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_256),
.B(n_228),
.C(n_203),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_365),
.B(n_239),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_367),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_173),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_369),
.B(n_373),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_286),
.A2(n_220),
.B1(n_5),
.B2(n_6),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_371),
.A2(n_374),
.B1(n_241),
.B2(n_316),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_240),
.B(n_4),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_307),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_280),
.B(n_7),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_379),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_277),
.B(n_7),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_380),
.A2(n_394),
.B(n_420),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_327),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_387),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_384),
.A2(n_392),
.B1(n_398),
.B2(n_422),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_320),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_378),
.Y(n_388)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_303),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_391),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_359),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_390),
.B(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_303),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_328),
.A2(n_310),
.B(n_264),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_417),
.Y(n_442)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_397),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_338),
.A2(n_269),
.B1(n_258),
.B2(n_301),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_328),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

INVx13_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_404),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_319),
.A2(n_290),
.B(n_283),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_407),
.A2(n_384),
.B(n_402),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_236),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_408),
.B(n_413),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_243),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_SL g411 ( 
.A(n_347),
.B(n_251),
.C(n_309),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_411),
.B(n_335),
.C(n_324),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_326),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_350),
.Y(n_413)
);

INVx3_ASAP7_75t_SL g414 ( 
.A(n_337),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_348),
.B(n_254),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_415),
.B(n_416),
.Y(n_435)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_248),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_347),
.B(n_245),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_426),
.Y(n_451)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_419),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g420 ( 
.A(n_318),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_318),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_421),
.A2(n_429),
.B(n_251),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_341),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_361),
.A2(n_261),
.B1(n_275),
.B2(n_284),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_423),
.A2(n_425),
.B1(n_376),
.B2(n_343),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_352),
.A2(n_262),
.B1(n_249),
.B2(n_233),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_347),
.B(n_305),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_330),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_427),
.A2(n_376),
.B(n_323),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_334),
.B(n_298),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_394),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_434),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_365),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_440),
.C(n_462),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_363),
.C(n_333),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_424),
.A2(n_381),
.B1(n_349),
.B2(n_393),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_443),
.A2(n_460),
.B1(n_471),
.B2(n_399),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_424),
.A2(n_381),
.B1(n_395),
.B2(n_393),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_444),
.A2(n_456),
.B1(n_466),
.B2(n_467),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_445),
.A2(n_469),
.B(n_427),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_407),
.A2(n_322),
.B(n_349),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_447),
.A2(n_448),
.B(n_465),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_424),
.A2(n_351),
.B(n_332),
.Y(n_448)
);

OAI32xp33_ASAP7_75t_L g452 ( 
.A1(n_409),
.A2(n_334),
.A3(n_362),
.B1(n_357),
.B2(n_333),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_415),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_358),
.B1(n_371),
.B2(n_374),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_405),
.A2(n_325),
.B1(n_285),
.B2(n_297),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_396),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_330),
.C(n_363),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_385),
.A2(n_332),
.B(n_353),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_413),
.A2(n_353),
.B1(n_331),
.B2(n_335),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_398),
.A2(n_331),
.B1(n_324),
.B2(n_323),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_410),
.B1(n_401),
.B2(n_429),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_390),
.A2(n_364),
.B1(n_368),
.B2(n_317),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_431),
.B(n_448),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_473),
.A2(n_474),
.B(n_476),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_383),
.B(n_428),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_456),
.A2(n_391),
.B1(n_389),
.B2(n_387),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_477),
.A2(n_485),
.B1(n_500),
.B2(n_506),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_445),
.A2(n_383),
.B(n_420),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_478),
.A2(n_479),
.B(n_483),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_469),
.A2(n_385),
.B(n_382),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_480),
.A2(n_482),
.B1(n_493),
.B2(n_494),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_443),
.A2(n_420),
.B(n_422),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_400),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_484),
.B(n_490),
.C(n_439),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_457),
.A2(n_408),
.B1(n_386),
.B2(n_400),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_386),
.Y(n_486)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

XNOR2x1_ASAP7_75t_SL g487 ( 
.A(n_434),
.B(n_388),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_487),
.A2(n_496),
.B(n_497),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_440),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_442),
.B(n_397),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_430),
.Y(n_491)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_491),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_416),
.Y(n_492)
);

CKINVDCx14_ASAP7_75t_R g542 ( 
.A(n_492),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_447),
.A2(n_406),
.B1(n_419),
.B2(n_414),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_457),
.A2(n_420),
.B(n_385),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_436),
.A2(n_412),
.B(n_377),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_498),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_465),
.A2(n_421),
.B(n_377),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_499),
.A2(n_511),
.B(n_446),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_436),
.A2(n_414),
.B1(n_321),
.B2(n_337),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_435),
.B(n_451),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_503),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_435),
.B(n_321),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_450),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_505),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_450),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_437),
.A2(n_368),
.B1(n_364),
.B2(n_329),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_463),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_507),
.B(n_508),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_437),
.A2(n_329),
.B1(n_336),
.B2(n_272),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_459),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_432),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_366),
.Y(n_510)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_459),
.A2(n_268),
.B(n_274),
.Y(n_511)
);

FAx1_ASAP7_75t_SL g515 ( 
.A(n_487),
.B(n_439),
.CI(n_461),
.CON(n_515),
.SN(n_515)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_515),
.B(n_532),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_492),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_516),
.B(n_525),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_519),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_499),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_521),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_488),
.B(n_462),
.C(n_440),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_524),
.B(n_526),
.C(n_529),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_508),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_489),
.C(n_481),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_488),
.B(n_441),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_530),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_528),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_490),
.B(n_449),
.C(n_464),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_484),
.B(n_449),
.Y(n_530)
);

AOI211xp5_ASAP7_75t_SL g531 ( 
.A1(n_480),
.A2(n_452),
.B(n_467),
.C(n_470),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_531),
.A2(n_475),
.B1(n_509),
.B2(n_485),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_326),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g581 ( 
.A(n_534),
.Y(n_581)
);

OA22x2_ASAP7_75t_L g535 ( 
.A1(n_494),
.A2(n_466),
.B1(n_464),
.B2(n_453),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_535),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_503),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_536),
.B(n_541),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_484),
.B(n_477),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_538),
.B(n_545),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_490),
.B(n_460),
.Y(n_540)
);

XNOR2x1_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_538),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_508),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_487),
.B(n_453),
.C(n_432),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_478),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_547),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_486),
.B(n_242),
.C(n_454),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_550),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_549),
.A2(n_479),
.B(n_496),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_486),
.B(n_510),
.C(n_505),
.Y(n_550)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_544),
.Y(n_554)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_554),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_512),
.A2(n_475),
.B1(n_473),
.B2(n_476),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_555),
.A2(n_566),
.B1(n_574),
.B2(n_580),
.Y(n_593)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_544),
.Y(n_556)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_556),
.Y(n_591)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_520),
.Y(n_560)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_560),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_504),
.B1(n_472),
.B2(n_482),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_561),
.A2(n_582),
.B1(n_543),
.B2(n_549),
.Y(n_599)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_520),
.Y(n_562)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

XNOR2x1_ASAP7_75t_L g597 ( 
.A(n_564),
.B(n_540),
.Y(n_597)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_565),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_518),
.B(n_501),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_572),
.B(n_576),
.Y(n_603)
);

INVx13_ASAP7_75t_L g573 ( 
.A(n_535),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_573),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_522),
.A2(n_473),
.B1(n_476),
.B2(n_483),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_575),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_527),
.B(n_542),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_533),
.Y(n_577)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_577),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_530),
.B(n_529),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_578),
.Y(n_602)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_579),
.B(n_583),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_517),
.A2(n_483),
.B1(n_472),
.B2(n_478),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_517),
.A2(n_482),
.B1(n_494),
.B2(n_500),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_584),
.B(n_535),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_543),
.A2(n_496),
.B1(n_500),
.B2(n_506),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_585),
.A2(n_521),
.B1(n_528),
.B2(n_547),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_553),
.B(n_559),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_587),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_553),
.B(n_526),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_569),
.B(n_519),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_588),
.B(n_568),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_SL g590 ( 
.A(n_569),
.B(n_550),
.Y(n_590)
);

XNOR2x1_ASAP7_75t_L g637 ( 
.A(n_590),
.B(n_597),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_570),
.B(n_524),
.C(n_559),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_595),
.C(n_605),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_570),
.B(n_548),
.C(n_545),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_581),
.B(n_438),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_596),
.B(n_552),
.Y(n_628)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_598),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_599),
.A2(n_574),
.B1(n_551),
.B2(n_562),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_561),
.A2(n_546),
.B1(n_531),
.B2(n_539),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_555),
.B1(n_585),
.B2(n_560),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_523),
.C(n_546),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_564),
.B(n_523),
.C(n_539),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_608),
.C(n_575),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_571),
.B(n_474),
.C(n_535),
.Y(n_608)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_611),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_566),
.A2(n_493),
.B1(n_515),
.B2(n_502),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_580),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_601),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_614),
.B(n_627),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_616),
.B(n_634),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_617),
.A2(n_619),
.B1(n_620),
.B2(n_630),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_556),
.Y(n_621)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_621),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_589),
.B(n_554),
.Y(n_622)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_622),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_557),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_624),
.B(n_625),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_603),
.B(n_568),
.Y(n_626)
);

CKINVDCx14_ASAP7_75t_R g646 ( 
.A(n_626),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_594),
.B(n_587),
.C(n_595),
.Y(n_627)
);

OAI321xp33_ASAP7_75t_L g643 ( 
.A1(n_628),
.A2(n_629),
.A3(n_600),
.B1(n_605),
.B2(n_610),
.C(n_607),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_607),
.A2(n_571),
.B(n_558),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_604),
.A2(n_551),
.B1(n_583),
.B2(n_584),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_599),
.A2(n_567),
.B1(n_558),
.B2(n_573),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_631),
.A2(n_632),
.B1(n_636),
.B2(n_598),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_613),
.A2(n_567),
.B1(n_579),
.B2(n_577),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_590),
.B(n_582),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_497),
.C(n_511),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_635),
.B(n_606),
.C(n_588),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_592),
.A2(n_565),
.B1(n_498),
.B2(n_495),
.Y(n_636)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_641),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_623),
.A2(n_611),
.B1(n_591),
.B2(n_609),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_642),
.A2(n_648),
.B1(n_651),
.B2(n_656),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_643),
.A2(n_652),
.B(n_641),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_615),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_627),
.B(n_602),
.C(n_593),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_650),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_623),
.A2(n_593),
.B1(n_608),
.B2(n_600),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_619),
.A2(n_491),
.B1(n_471),
.B2(n_515),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_649),
.A2(n_654),
.B1(n_629),
.B2(n_621),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_618),
.B(n_597),
.C(n_454),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_633),
.A2(n_468),
.B1(n_446),
.B2(n_458),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_620),
.A2(n_468),
.B1(n_455),
.B2(n_433),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_625),
.B(n_404),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g674 ( 
.A(n_655),
.B(n_637),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_633),
.A2(n_433),
.B1(n_336),
.B2(n_372),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_433),
.C(n_344),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_657),
.B(n_615),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_660),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_647),
.B(n_628),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_661),
.B(n_662),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_645),
.B(n_622),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_663),
.A2(n_664),
.B1(n_667),
.B2(n_669),
.Y(n_678)
);

INVx11_ASAP7_75t_L g664 ( 
.A(n_646),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_655),
.B(n_634),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g677 ( 
.A(n_665),
.B(n_674),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_670),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_638),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_640),
.B(n_624),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_639),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_671),
.B(n_673),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_640),
.B(n_631),
.C(n_616),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_657),
.C(n_653),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_635),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_676),
.B(n_679),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_662),
.B(n_672),
.Y(n_679)
);

AOI321xp33_ASAP7_75t_L g681 ( 
.A1(n_664),
.A2(n_644),
.A3(n_650),
.B1(n_648),
.B2(n_637),
.C(n_649),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_681),
.B(n_685),
.Y(n_694)
);

XOR2xp5_ASAP7_75t_L g684 ( 
.A(n_673),
.B(n_639),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_684),
.B(n_665),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_671),
.B(n_642),
.Y(n_685)
);

NAND4xp25_ASAP7_75t_SL g686 ( 
.A(n_663),
.B(n_654),
.C(n_651),
.D(n_404),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_686),
.B(n_372),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_SL g687 ( 
.A1(n_678),
.A2(n_668),
.B(n_658),
.C(n_656),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_687),
.A2(n_689),
.B(n_690),
.Y(n_700)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_688),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_683),
.A2(n_658),
.B(n_659),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_SL g690 ( 
.A(n_680),
.B(n_674),
.Y(n_690)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_682),
.B(n_372),
.C(n_344),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_691),
.B(n_692),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_683),
.A2(n_306),
.B(n_253),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_SL g697 ( 
.A1(n_695),
.A2(n_260),
.B1(n_250),
.B2(n_237),
.Y(n_697)
);

A2O1A1O1Ixp25_ASAP7_75t_L g696 ( 
.A1(n_694),
.A2(n_675),
.B(n_684),
.C(n_677),
.D(n_686),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_696),
.Y(n_701)
);

MAJIxp5_ASAP7_75t_L g702 ( 
.A(n_697),
.B(n_699),
.C(n_689),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_702),
.A2(n_703),
.B(n_677),
.Y(n_704)
);

MAJIxp5_ASAP7_75t_L g703 ( 
.A(n_698),
.B(n_693),
.C(n_700),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_SL g706 ( 
.A(n_704),
.B(n_705),
.C(n_312),
.Y(n_706)
);

AOI21x1_ASAP7_75t_SL g705 ( 
.A1(n_701),
.A2(n_366),
.B(n_343),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_SL g707 ( 
.A1(n_706),
.A2(n_287),
.B(n_263),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_707),
.A2(n_267),
.B(n_235),
.Y(n_708)
);

MAJx2_ASAP7_75t_L g709 ( 
.A(n_708),
.B(n_270),
.C(n_7),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_709),
.A2(n_7),
.B1(n_8),
.B2(n_446),
.Y(n_710)
);


endmodule