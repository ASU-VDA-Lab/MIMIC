module real_jpeg_24104_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_19),
.B1(n_22),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_18)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_3),
.A2(n_21),
.B1(n_54),
.B2(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_19),
.B1(n_22),
.B2(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_25),
.C(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_40),
.B1(n_92),
.B2(n_98),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_19),
.B1(n_22),
.B2(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_74),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_51),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_15),
.B(n_51),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_34),
.C(n_39),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_16),
.A2(n_17),
.B1(n_34),
.B2(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_18),
.A2(n_23),
.B1(n_31),
.B2(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g22 ( 
.A(n_19),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g36 ( 
.A1(n_19),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g53 ( 
.A1(n_19),
.A2(n_37),
.A3(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_19),
.B(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_38),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_28),
.B(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_29),
.B(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_56),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_38),
.B1(n_54),
.B2(n_57),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_46),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_41),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_44),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_67),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_54),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_58),
.CON(n_56),
.SN(n_56)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_85),
.B(n_106),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_81),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_94),
.B(n_105),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_100),
.B(n_104),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);


endmodule