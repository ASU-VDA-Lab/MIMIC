module fake_netlist_1_11391_n_647 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_647);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_647;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_55), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_35), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_52), .Y(n_78) );
INVxp33_ASAP7_75t_SL g79 ( .A(n_67), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_40), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_11), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_42), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_34), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_7), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_11), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_32), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_9), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_72), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_51), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_30), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_31), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_5), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_29), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_56), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_12), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_20), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_2), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_21), .Y(n_101) );
BUFx5_ASAP7_75t_L g102 ( .A(n_70), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_9), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_3), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_41), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_43), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_54), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_27), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_4), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_53), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_14), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_0), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_118), .B(n_0), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_76), .B(n_1), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_78), .A2(n_39), .B(n_74), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_109), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_113), .B(n_1), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_102), .B(n_2), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_96), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_112), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_112), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_102), .B(n_3), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_109), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_116), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_88), .B(n_4), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_101), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_108), .A2(n_6), .B1(n_10), .B2(n_12), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_91), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_102), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
BUFx8_ASAP7_75t_L g148 ( .A(n_102), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_98), .Y(n_149) );
NOR2x1_ASAP7_75t_L g150 ( .A(n_82), .B(n_47), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_98), .B(n_10), .Y(n_151) );
NOR2xp33_ASAP7_75t_R g152 ( .A(n_77), .B(n_48), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_77), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_84), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_129), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_153), .B(n_89), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_149), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_153), .B(n_104), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_148), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_138), .B(n_124), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
NOR2x1p5_ASAP7_75t_L g165 ( .A(n_154), .B(n_87), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_154), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_135), .B(n_88), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_125), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_122), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_137), .B(n_89), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_127), .B(n_84), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_138), .B(n_124), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_138), .A2(n_79), .B1(n_80), .B2(n_114), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_124), .B(n_117), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_137), .B(n_87), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_148), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_144), .B(n_92), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
BUFx10_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_148), .B(n_92), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_150), .B(n_99), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_141), .A2(n_100), .B1(n_86), .B2(n_94), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_140), .B(n_105), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_151), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_136), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_122), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_178), .B(n_147), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_192), .Y(n_199) );
INVx5_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_192), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_163), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_180), .B(n_147), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_178), .B(n_145), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_180), .B(n_142), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_162), .B(n_145), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_162), .B(n_143), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_180), .B(n_143), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_180), .B(n_120), .Y(n_210) );
INVx5_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_157), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_195), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_163), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_196), .B(n_119), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_170), .B(n_110), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_195), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_173), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_174), .A2(n_79), .B1(n_80), .B2(n_132), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_172), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_159), .Y(n_225) );
AO22x1_ASAP7_75t_L g226 ( .A1(n_166), .A2(n_93), .B1(n_105), .B2(n_115), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_195), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_191), .B(n_136), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_195), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_171), .B(n_93), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
INVxp33_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
NOR2xp33_ASAP7_75t_R g234 ( .A(n_181), .B(n_131), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_185), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_177), .B(n_131), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_172), .Y(n_238) );
NOR3xp33_ASAP7_75t_SL g239 ( .A(n_186), .B(n_103), .C(n_128), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_170), .B(n_111), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_190), .B(n_130), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_176), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_170), .B(n_107), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_176), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_197), .A2(n_106), .B(n_126), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_167), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_167), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_174), .A2(n_130), .B1(n_126), .B2(n_121), .Y(n_249) );
OAI21xp33_ASAP7_75t_L g250 ( .A1(n_233), .A2(n_156), .B(n_179), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_236), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_224), .B(n_165), .Y(n_252) );
INVxp67_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_206), .A2(n_199), .B1(n_201), .B2(n_238), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_233), .B(n_166), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_234), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_242), .B(n_206), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_228), .Y(n_258) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_211), .B(n_170), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_242), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_203), .B(n_165), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_209), .B(n_187), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_211), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_247), .B(n_187), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_206), .A2(n_182), .B1(n_197), .B2(n_170), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_217), .A2(n_197), .B(n_170), .Y(n_269) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_232), .B(n_96), .Y(n_270) );
BUFx8_ASAP7_75t_SL g271 ( .A(n_212), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_248), .B(n_184), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_211), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_236), .Y(n_274) );
AND3x1_ASAP7_75t_SL g275 ( .A(n_226), .B(n_121), .C(n_14), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_220), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_213), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_232), .B(n_181), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_223), .B(n_13), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_217), .A2(n_193), .B(n_185), .Y(n_281) );
CKINVDCx6p67_ASAP7_75t_R g282 ( .A(n_200), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_220), .A2(n_183), .B1(n_184), .B2(n_188), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_232), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_213), .Y(n_285) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_220), .B(n_183), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_219), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_244), .A2(n_184), .B1(n_161), .B2(n_188), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_202), .Y(n_290) );
INVx8_ASAP7_75t_L g291 ( .A(n_200), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_246), .A2(n_168), .B1(n_161), .B2(n_175), .Y(n_292) );
OAI22x1_ASAP7_75t_L g293 ( .A1(n_216), .A2(n_13), .B1(n_15), .B2(n_181), .Y(n_293) );
INVx5_ASAP7_75t_L g294 ( .A(n_200), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_227), .Y(n_295) );
NAND2x1_ASAP7_75t_L g296 ( .A(n_251), .B(n_229), .Y(n_296) );
AO31x2_ASAP7_75t_L g297 ( .A1(n_293), .A2(n_245), .A3(n_231), .B(n_235), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_269), .A2(n_243), .B(n_240), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_259), .A2(n_243), .B(n_240), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_259), .A2(n_241), .B(n_237), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_258), .B(n_214), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_253), .B(n_198), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_270), .A2(n_210), .B1(n_204), .B2(n_215), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_255), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_255), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_256), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_281), .A2(n_205), .B(n_198), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_257), .B(n_205), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g313 ( .A1(n_267), .A2(n_230), .B1(n_249), .B2(n_218), .Y(n_313) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_292), .A2(n_239), .B(n_207), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_259), .A2(n_207), .B(n_208), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_254), .B(n_222), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_266), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_257), .B(n_221), .Y(n_321) );
OR2x2_ASAP7_75t_SL g322 ( .A(n_260), .B(n_96), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_257), .A2(n_208), .B1(n_181), .B2(n_200), .Y(n_323) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_295), .A2(n_168), .B(n_175), .Y(n_324) );
OAI21x1_ASAP7_75t_L g325 ( .A1(n_289), .A2(n_183), .B(n_193), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_270), .B(n_193), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
NOR2x1_ASAP7_75t_L g328 ( .A(n_324), .B(n_280), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_313), .A2(n_257), .B1(n_252), .B2(n_250), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_320), .B(n_263), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_324), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_307), .A2(n_252), .B1(n_293), .B2(n_272), .C(n_264), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_308), .B(n_252), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_324), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_305), .A2(n_314), .B1(n_311), .B2(n_309), .Y(n_335) );
BUFx2_ASAP7_75t_SL g336 ( .A(n_324), .Y(n_336) );
OAI221xp5_ASAP7_75t_L g337 ( .A1(n_318), .A2(n_268), .B1(n_283), .B2(n_261), .C(n_284), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_303), .Y(n_338) );
OAI211xp5_ASAP7_75t_L g339 ( .A1(n_303), .A2(n_286), .B(n_275), .C(n_276), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_310), .A2(n_285), .B(n_278), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_317), .B(n_284), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_302), .A2(n_279), .B(n_265), .C(n_288), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_327), .Y(n_343) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_306), .B(n_96), .C(n_279), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_299), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_309), .A2(n_291), .B1(n_273), .B2(n_271), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_299), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_314), .A2(n_271), .B1(n_282), .B2(n_291), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_302), .A2(n_285), .B(n_288), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_312), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_314), .A2(n_282), .B1(n_291), .B2(n_265), .Y(n_352) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_325), .A2(n_287), .B(n_185), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_322), .A2(n_287), .B1(n_294), .B2(n_273), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_334), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_334), .B(n_301), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_330), .B(n_317), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_345), .B(n_327), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_345), .B(n_316), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_345), .B(n_316), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_347), .B(n_319), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_347), .B(n_348), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_347), .B(n_319), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_331), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_348), .B(n_297), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_348), .B(n_297), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_351), .B(n_297), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_331), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_351), .B(n_297), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_353), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_353), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_343), .B(n_297), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_301), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_328), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_335), .B(n_321), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_378), .B(n_350), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_378), .B(n_342), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_358), .A2(n_344), .B(n_332), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_372), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_357), .B(n_338), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_355), .B(n_322), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_381), .A2(n_344), .B1(n_354), .B2(n_339), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_357), .B(n_329), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_383), .A2(n_346), .B1(n_349), .B2(n_333), .C(n_321), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_381), .B(n_325), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_374), .B(n_352), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_368), .B(n_96), .Y(n_401) );
AO21x2_ASAP7_75t_L g402 ( .A1(n_379), .A2(n_340), .B(n_298), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_368), .B(n_301), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_382), .B(n_341), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_370), .B(n_298), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_370), .B(n_15), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_362), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_364), .B(n_315), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_362), .B(n_300), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_373), .B(n_300), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_383), .A2(n_304), .B1(n_337), .B2(n_323), .C(n_326), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_367), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_373), .B(n_315), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_379), .B(n_296), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_380), .B(n_359), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_371), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_374), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_364), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_356), .B(n_296), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_380), .B(n_294), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_407), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_397), .B(n_382), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_403), .B(n_384), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_396), .A2(n_384), .B1(n_377), .B2(n_376), .C(n_375), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_403), .B(n_377), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_421), .B(n_360), .Y(n_433) );
INVx3_ASAP7_75t_SL g434 ( .A(n_407), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_397), .B(n_382), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_407), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_398), .B(n_376), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_409), .B(n_361), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_424), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_403), .B(n_375), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_409), .B(n_361), .Y(n_442) );
AND3x2_ASAP7_75t_L g443 ( .A(n_409), .B(n_360), .C(n_365), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_398), .B(n_371), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_408), .B(n_371), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_408), .B(n_371), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_389), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_408), .B(n_356), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_424), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g451 ( .A(n_396), .B(n_359), .C(n_356), .D(n_363), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_390), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_356), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_391), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_389), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_425), .B(n_365), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_389), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_414), .B(n_363), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_425), .B(n_294), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_16), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_419), .B(n_401), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_405), .B(n_277), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_388), .B(n_405), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_419), .B(n_18), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_419), .B(n_19), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_401), .B(n_22), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_406), .A2(n_277), .B1(n_262), .B2(n_291), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_401), .B(n_23), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_420), .B(n_24), .Y(n_471) );
NOR3xp33_ASAP7_75t_SL g472 ( .A(n_416), .B(n_26), .C(n_28), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_420), .B(n_33), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_420), .B(n_38), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_390), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_411), .B(n_44), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_390), .B(n_277), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_387), .B(n_294), .C(n_273), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_411), .B(n_415), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_415), .B(n_45), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_415), .B(n_46), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_417), .Y(n_483) );
NAND4xp25_ASAP7_75t_SL g484 ( .A(n_469), .B(n_479), .C(n_438), .D(n_442), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_465), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_460), .B(n_426), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
NAND2xp33_ASAP7_75t_SL g490 ( .A(n_434), .B(n_392), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_436), .B(n_386), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_480), .B(n_386), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_433), .B(n_394), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_480), .B(n_394), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_460), .B(n_386), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_479), .A2(n_393), .B(n_387), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_392), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_430), .B(n_426), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_430), .B(n_426), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_454), .B(n_394), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_454), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_476), .B(n_418), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_455), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_468), .B(n_406), .Y(n_504) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_439), .B(n_450), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_455), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_457), .B(n_406), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_459), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_449), .B(n_386), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_476), .B(n_418), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_473), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_483), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_483), .B(n_418), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_437), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_437), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_443), .B(n_395), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_463), .B(n_395), .Y(n_520) );
OR2x2_ASAP7_75t_SL g521 ( .A(n_451), .B(n_395), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_463), .B(n_386), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_432), .B(n_410), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_432), .Y(n_524) );
AND2x2_ASAP7_75t_SL g525 ( .A(n_428), .B(n_397), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_453), .B(n_423), .Y(n_526) );
AND3x2_ASAP7_75t_L g527 ( .A(n_471), .B(n_427), .C(n_397), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_434), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_453), .B(n_423), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_441), .B(n_410), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_441), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_451), .A2(n_416), .B(n_400), .C(n_385), .Y(n_532) );
BUFx2_ASAP7_75t_SL g533 ( .A(n_436), .Y(n_533) );
NAND2x1_ASAP7_75t_SL g534 ( .A(n_434), .B(n_397), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_449), .B(n_410), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_444), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_444), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_462), .B(n_413), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_464), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_487), .B(n_445), .Y(n_540) );
AOI211x1_ASAP7_75t_L g541 ( .A1(n_484), .A2(n_431), .B(n_471), .C(n_474), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_521), .A2(n_469), .B1(n_428), .B2(n_448), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_493), .B(n_461), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_505), .B(n_428), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_517), .B(n_445), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_505), .Y(n_546) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_528), .A2(n_428), .B1(n_448), .B2(n_474), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_490), .A2(n_472), .B(n_448), .C(n_475), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_435), .B1(n_429), .B2(n_475), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_518), .B(n_446), .Y(n_550) );
NOR2xp67_ASAP7_75t_SL g551 ( .A(n_533), .B(n_468), .Y(n_551) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_496), .A2(n_393), .B(n_435), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_532), .A2(n_462), .B(n_466), .C(n_467), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_525), .B(n_466), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_490), .A2(n_435), .B1(n_429), .B2(n_467), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_515), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_488), .B(n_477), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_524), .B(n_477), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_492), .B(n_495), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_532), .A2(n_470), .B(n_481), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_525), .B(n_470), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_531), .B(n_494), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_504), .A2(n_478), .B1(n_435), .B2(n_429), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_486), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_489), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_519), .B(n_482), .C(n_481), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_501), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_503), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_511), .A2(n_464), .B(n_458), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_511), .A2(n_422), .B(n_385), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_536), .B(n_446), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_537), .B(n_429), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_491), .A2(n_447), .B1(n_456), .B2(n_458), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_539), .B(n_456), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_534), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_491), .A2(n_385), .B1(n_413), .B2(n_478), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_491), .B(n_447), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_540), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_560), .B(n_495), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_556), .Y(n_584) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_541), .B(n_527), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_551), .Y(n_586) );
OAI322xp33_ASAP7_75t_L g587 ( .A1(n_566), .A2(n_497), .A3(n_507), .B1(n_502), .B2(n_512), .C1(n_500), .C2(n_535), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_564), .B(n_492), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_557), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_546), .B(n_504), .Y(n_590) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_566), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_553), .A2(n_482), .B(n_522), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_553), .A2(n_527), .B(n_510), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_546), .B(n_510), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_543), .B(n_529), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_563), .A2(n_520), .B1(n_530), .B2(n_523), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_562), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_567), .Y(n_598) );
AOI322xp5_ASAP7_75t_L g599 ( .A1(n_552), .A2(n_498), .A3(n_499), .B1(n_526), .B2(n_514), .C1(n_513), .C2(n_509), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_555), .A2(n_538), .B1(n_516), .B2(n_485), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_542), .B(n_485), .C(n_404), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_545), .B(n_385), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g603 ( .A1(n_561), .A2(n_385), .B1(n_413), .B2(n_422), .C1(n_399), .C2(n_404), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_550), .B(n_413), .Y(n_604) );
NAND2xp33_ASAP7_75t_SL g605 ( .A(n_581), .B(n_422), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_573), .B(n_404), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_569), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_597), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_599), .B(n_580), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_587), .A2(n_571), .B1(n_549), .B2(n_547), .C(n_559), .Y(n_610) );
CKINVDCx20_ASAP7_75t_L g611 ( .A(n_586), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_593), .A2(n_548), .B1(n_544), .B2(n_575), .C(n_554), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_598), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_SL g614 ( .A1(n_601), .A2(n_568), .B(n_572), .C(n_565), .Y(n_614) );
OAI222xp33_ASAP7_75t_L g615 ( .A1(n_596), .A2(n_578), .B1(n_558), .B2(n_572), .C1(n_574), .C2(n_579), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_585), .A2(n_576), .B1(n_570), .B2(n_577), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g617 ( .A1(n_603), .A2(n_404), .B1(n_399), .B2(n_413), .C(n_402), .Y(n_617) );
AOI221x1_ASAP7_75t_L g618 ( .A1(n_605), .A2(n_399), .B1(n_402), .B2(n_277), .C(n_262), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g619 ( .A1(n_585), .A2(n_399), .B1(n_294), .B2(n_277), .C1(n_262), .C2(n_273), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_592), .A2(n_273), .B1(n_262), .B2(n_402), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_589), .B(n_402), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_590), .A2(n_169), .B1(n_164), .B2(n_189), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_611), .A2(n_600), .B1(n_590), .B2(n_582), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_608), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_617), .A2(n_600), .B1(n_591), .B2(n_584), .C(n_607), .Y(n_625) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_622), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_614), .A2(n_605), .B(n_595), .Y(n_627) );
AO22x1_ASAP7_75t_L g628 ( .A1(n_609), .A2(n_588), .B1(n_594), .B2(n_583), .Y(n_628) );
AOI221x1_ASAP7_75t_L g629 ( .A1(n_613), .A2(n_621), .B1(n_620), .B2(n_619), .C(n_615), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_616), .A2(n_602), .B1(n_604), .B2(n_583), .C(n_606), .Y(n_630) );
OAI21xp33_ASAP7_75t_SL g631 ( .A1(n_610), .A2(n_49), .B(n_50), .Y(n_631) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_627), .B(n_612), .Y(n_632) );
NAND4xp75_ASAP7_75t_L g633 ( .A(n_629), .B(n_618), .C(n_617), .D(n_61), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_631), .A2(n_57), .B1(n_58), .B2(n_62), .C(n_63), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_624), .B(n_64), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_626), .B(n_65), .Y(n_636) );
OAI22x1_ASAP7_75t_L g637 ( .A1(n_632), .A2(n_623), .B1(n_628), .B2(n_625), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_633), .B(n_630), .C(n_624), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_634), .B(n_160), .C(n_155), .D(n_158), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_637), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_638), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_640), .A2(n_636), .B1(n_635), .B2(n_639), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_641), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_643), .A2(n_635), .B1(n_160), .B2(n_155), .C1(n_158), .C2(n_73), .Y(n_644) );
OA22x2_ASAP7_75t_L g645 ( .A1(n_644), .A2(n_642), .B1(n_155), .B2(n_158), .Y(n_645) );
AOI211x1_ASAP7_75t_L g646 ( .A1(n_645), .A2(n_66), .B(n_68), .C(n_69), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_646), .A2(n_164), .B1(n_169), .B2(n_189), .C(n_75), .Y(n_647) );
endmodule