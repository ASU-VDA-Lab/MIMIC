module fake_jpeg_12034_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_56),
.Y(n_98)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_61),
.B(n_68),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_16),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_80),
.C(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_30),
.B1(n_15),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_64),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_30),
.B1(n_15),
.B2(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_30),
.B1(n_19),
.B2(n_32),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_78),
.B1(n_23),
.B2(n_22),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_85),
.B1(n_23),
.B2(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_33),
.B1(n_21),
.B2(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_0),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_24),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_32),
.B1(n_17),
.B2(n_29),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_95),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_20),
.C(n_25),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_82),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_46),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_118),
.B(n_103),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_74),
.B1(n_76),
.B2(n_18),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_122),
.Y(n_142)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_20),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_31),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_31),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_46),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_52),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_62),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_0),
.B(n_1),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_63),
.B(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_125),
.A2(n_150),
.B(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_80),
.C(n_60),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_130),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_65),
.B1(n_55),
.B2(n_75),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_127),
.A2(n_128),
.B1(n_140),
.B2(n_155),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_55),
.B1(n_54),
.B2(n_66),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_133),
.B1(n_136),
.B2(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_132),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_54),
.B1(n_66),
.B2(n_52),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_89),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_138),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_53),
.B1(n_59),
.B2(n_86),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_11),
.B(n_10),
.C(n_9),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_137),
.A2(n_10),
.B(n_13),
.C(n_12),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_139),
.B(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_74),
.B1(n_76),
.B2(n_18),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_31),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_31),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_102),
.A2(n_103),
.B1(n_92),
.B2(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_159),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_0),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_1),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_99),
.B1(n_110),
.B2(n_119),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_161),
.A2(n_190),
.B1(n_126),
.B2(n_142),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_164),
.B(n_173),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_195),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_114),
.B1(n_99),
.B2(n_113),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_178),
.B1(n_180),
.B2(n_184),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_114),
.B1(n_113),
.B2(n_104),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_117),
.B1(n_96),
.B2(n_97),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_145),
.B1(n_160),
.B2(n_143),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_97),
.B(n_121),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_156),
.B(n_130),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_121),
.B1(n_9),
.B2(n_10),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_194),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_2),
.B(n_3),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_4),
.B(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_14),
.C(n_5),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_221),
.B(n_162),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_130),
.B(n_155),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_202),
.B(n_211),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_168),
.B(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_183),
.Y(n_246)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_137),
.A3(n_134),
.B1(n_158),
.B2(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_218),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_135),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_208),
.C(n_210),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_140),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_128),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_128),
.B(n_132),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_159),
.B(n_154),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_217),
.B(n_199),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_193),
.B(n_4),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_223),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_7),
.B(n_161),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_SL g223 ( 
.A(n_172),
.B(n_179),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_166),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_202),
.C(n_223),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_192),
.B(n_217),
.Y(n_257)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_195),
.B1(n_189),
.B2(n_171),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_162),
.B1(n_180),
.B2(n_178),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_208),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_187),
.B1(n_177),
.B2(n_171),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_243),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_200),
.B1(n_211),
.B2(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_177),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_205),
.B(n_222),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_255),
.C(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_264),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_258),
.B(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_220),
.C(n_183),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_231),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_245),
.B(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_214),
.C(n_181),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_214),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_244),
.B(n_238),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_252),
.A2(n_241),
.B1(n_244),
.B2(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_268),
.A2(n_278),
.B1(n_261),
.B2(n_259),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_240),
.C(n_237),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_277),
.C(n_272),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_257),
.B(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_239),
.B1(n_227),
.B2(n_243),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_274),
.B(n_248),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_227),
.C(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_249),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_285),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_255),
.C(n_253),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_290),
.C(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_251),
.C(n_247),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_270),
.B(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_297),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_295),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_280),
.B1(n_283),
.B2(n_270),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_265),
.B1(n_277),
.B2(n_269),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_267),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_278),
.B1(n_275),
.B2(n_228),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_285),
.B1(n_286),
.B2(n_212),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_292),
.C(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_212),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_294),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_301),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_301),
.B1(n_300),
.B2(n_304),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_312),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_309),
.B1(n_302),
.B2(n_181),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_163),
.B(n_174),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_176),
.B(n_169),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_191),
.Y(n_318)
);


endmodule