module fake_jpeg_15749_n_349 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_0),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_24),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_53),
.B(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_37),
.B1(n_26),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_70),
.B1(n_51),
.B2(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_24),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_76),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_22),
.B1(n_37),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_73),
.B1(n_36),
.B2(n_21),
.Y(n_96)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_37),
.B1(n_22),
.B2(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_32),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_37),
.B1(n_33),
.B2(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_29),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_34),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_34),
.B(n_32),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_83),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_96),
.B1(n_77),
.B2(n_51),
.Y(n_124)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_70),
.C(n_60),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_107),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_109),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_78),
.Y(n_103)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_36),
.B(n_34),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_77),
.B(n_19),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_51),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_115),
.B(n_86),
.Y(n_143)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_64),
.B1(n_105),
.B2(n_71),
.Y(n_146)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_57),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_125),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_55),
.B1(n_64),
.B2(n_54),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_115),
.B1(n_124),
.B2(n_55),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_78),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_50),
.C(n_49),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_50),
.C(n_49),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_146),
.B1(n_152),
.B2(n_103),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_147),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_97),
.C(n_83),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_162),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_69),
.B1(n_66),
.B2(n_58),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_69),
.B1(n_59),
.B2(n_102),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_69),
.B1(n_102),
.B2(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_86),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_155),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_40),
.B1(n_135),
.B2(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_101),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_40),
.B1(n_128),
.B2(n_84),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_113),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_44),
.B1(n_45),
.B2(n_42),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_123),
.B1(n_126),
.B2(n_111),
.Y(n_184)
);

XOR2x2_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_113),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_172),
.B(n_190),
.Y(n_192)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_122),
.A3(n_137),
.B1(n_97),
.B2(n_62),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_150),
.B1(n_142),
.B2(n_144),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_132),
.B1(n_130),
.B2(n_129),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_180),
.B1(n_184),
.B2(n_187),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_137),
.B(n_47),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_47),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_160),
.C(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_62),
.B1(n_123),
.B2(n_121),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_28),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_151),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_29),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_45),
.B1(n_44),
.B2(n_42),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_0),
.B(n_1),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_28),
.B(n_19),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_142),
.B(n_164),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_157),
.B(n_154),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_199),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_205),
.B1(n_185),
.B2(n_167),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_164),
.B(n_149),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_210),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_166),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_207),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_159),
.B1(n_160),
.B2(n_116),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_89),
.C(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_30),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_47),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_78),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_213),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_131),
.B(n_27),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_30),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_45),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_217),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_131),
.C(n_44),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_98),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_229),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_177),
.B1(n_178),
.B2(n_173),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_223),
.B1(n_228),
.B2(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_177),
.B1(n_190),
.B2(n_167),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_236),
.B1(n_214),
.B2(n_206),
.Y(n_250)
);

XNOR2x2_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_191),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_225),
.B(n_192),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_242),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_184),
.B1(n_175),
.B2(n_114),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_114),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_194),
.A2(n_112),
.B1(n_106),
.B2(n_104),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_197),
.B1(n_205),
.B2(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_112),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_204),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_257),
.B1(n_236),
.B2(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_252),
.B(n_263),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_249),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_201),
.B1(n_192),
.B2(n_202),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_193),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_211),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.C(n_265),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_213),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_235),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_273),
.C(n_274),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_229),
.B1(n_240),
.B2(n_228),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_250),
.B1(n_248),
.B2(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_216),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_238),
.C(n_215),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_223),
.C(n_216),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_282),
.C(n_25),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_31),
.B1(n_12),
.B2(n_13),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_259),
.B1(n_244),
.B2(n_264),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_287),
.B1(n_267),
.B2(n_282),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_25),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_293),
.C(n_299),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_25),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_12),
.B(n_17),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_11),
.B(n_16),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_8),
.B(n_15),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_10),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_31),
.C(n_23),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_31),
.B1(n_10),
.B2(n_11),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_303),
.B(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_280),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_267),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_295),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_290),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_286),
.A2(n_283),
.B1(n_269),
.B2(n_31),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_293),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_297),
.B1(n_292),
.B2(n_287),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_283),
.C(n_23),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_23),
.C(n_18),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_8),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_15),
.B(n_9),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_320),
.C(n_322),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_27),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_298),
.CI(n_299),
.CON(n_319),
.SN(n_319)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_301),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_302),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_18),
.C(n_27),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_18),
.C(n_27),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_314),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_326),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_302),
.B(n_3),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_0),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_317),
.A2(n_313),
.B(n_312),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_329),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_331),
.A2(n_333),
.B(n_330),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_334),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_2),
.B(n_3),
.Y(n_335)
);

OAI211xp5_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_321),
.B(n_318),
.C(n_320),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_319),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_336),
.A2(n_338),
.B(n_340),
.C(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_323),
.B(n_322),
.Y(n_341)
);

AOI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_339),
.A2(n_3),
.B(n_4),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_343),
.A2(n_344),
.B(n_4),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_4),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_342),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_5),
.B(n_6),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_347),
.A2(n_5),
.B(n_6),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_6),
.B(n_27),
.Y(n_349)
);


endmodule