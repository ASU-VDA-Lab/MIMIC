module fake_jpeg_24937_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

CKINVDCx11_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_28),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_53)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_85),
.B1(n_34),
.B2(n_36),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_35),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_74),
.Y(n_103)
);

CKINVDCx9p33_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_69),
.B1(n_17),
.B2(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_35),
.B1(n_23),
.B2(n_27),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_20),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_46),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_27),
.C(n_33),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_1),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_34),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_104),
.B1(n_30),
.B2(n_17),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_116),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_36),
.B1(n_23),
.B2(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_105),
.B1(n_69),
.B2(n_26),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_77),
.B1(n_29),
.B2(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_108),
.B1(n_28),
.B2(n_32),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_84),
.B1(n_26),
.B2(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_24),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_120),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_55),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_119),
.B(n_122),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_63),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_92),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_128),
.B1(n_104),
.B2(n_88),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_94),
.B1(n_117),
.B2(n_90),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_60),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_102),
.B1(n_103),
.B2(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_128),
.B1(n_132),
.B2(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_60),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_87),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_144),
.C(n_145),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_32),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_88),
.B1(n_111),
.B2(n_90),
.Y(n_149)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_115),
.B(n_104),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_75),
.B(n_67),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_22),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_54),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_94),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_146),
.B1(n_101),
.B2(n_107),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_151),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.C(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_22),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_176),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_22),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_144),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_22),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_127),
.A2(n_130),
.B1(n_137),
.B2(n_136),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_174),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_176),
.B1(n_168),
.B2(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_188),
.B1(n_191),
.B2(n_164),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_154),
.B(n_175),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_166),
.B(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_180),
.B(n_8),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_135),
.B1(n_141),
.B2(n_101),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_186),
.B1(n_189),
.B2(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_195),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_1),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_2),
.B(n_4),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_159),
.B(n_160),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_156),
.C(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_2),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_168),
.B1(n_169),
.B2(n_152),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_6),
.B(n_7),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_205),
.B(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_206),
.C(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_202),
.Y(n_224)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_208),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_173),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_153),
.C(n_7),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_183),
.B(n_153),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_212),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_164),
.C(n_171),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_171),
.C(n_9),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_197),
.C(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_198),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_209),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_184),
.C(n_185),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_225),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_178),
.B(n_181),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_209),
.B(n_10),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_185),
.C(n_196),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_181),
.B(n_193),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_239),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_207),
.C(n_211),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_187),
.B(n_179),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_233),
.Y(n_245)
);

AOI31xp67_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_209),
.A3(n_179),
.B(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_227),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_216),
.C(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_246),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_239),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_225),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_238),
.A3(n_235),
.B1(n_230),
.B2(n_232),
.C1(n_231),
.C2(n_228),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_254),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_251),
.A2(n_246),
.B1(n_248),
.B2(n_244),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_255),
.Y(n_259)
);

AOI21x1_ASAP7_75t_SL g260 ( 
.A1(n_256),
.A2(n_242),
.B(n_250),
.Y(n_260)
);

OAI322xp33_ASAP7_75t_L g263 ( 
.A1(n_260),
.A2(n_258),
.A3(n_242),
.B1(n_247),
.B2(n_241),
.C1(n_216),
.C2(n_11),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_258),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_259),
.Y(n_265)
);


endmodule