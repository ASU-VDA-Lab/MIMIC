module real_aes_12030_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_905;
wire n_357;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_523;
wire n_298;
wire n_781;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g556 ( .A(n_0), .B(n_148), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_1), .A2(n_84), .B1(n_555), .B2(n_585), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g923 ( .A1(n_2), .A2(n_529), .B(n_924), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_3), .B(n_182), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_4), .B(n_164), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_5), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_6), .A2(n_36), .B1(n_138), .B2(n_572), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_7), .B(n_86), .Y(n_517) );
INVx1_ASAP7_75t_L g934 ( .A(n_7), .Y(n_934) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_8), .B(n_140), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_9), .B(n_121), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_10), .A2(n_63), .B1(n_138), .B2(n_258), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_11), .B(n_138), .C(n_141), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_12), .B(n_121), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_13), .B(n_179), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_14), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_15), .B(n_606), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_16), .B(n_128), .Y(n_633) );
AND2x2_ASAP7_75t_L g257 ( .A(n_17), .B(n_258), .Y(n_257) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_18), .B(n_134), .C(n_140), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_19), .A2(n_26), .B1(n_140), .B2(n_572), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_20), .B(n_606), .Y(n_618) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_21), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_22), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_23), .B(n_147), .Y(n_215) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_24), .B(n_197), .Y(n_196) );
NAND2xp33_ASAP7_75t_L g245 ( .A(n_25), .B(n_197), .Y(n_245) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_27), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_28), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_29), .B(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_30), .A2(n_50), .B1(n_197), .B2(n_258), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_31), .B(n_134), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_32), .B(n_163), .Y(n_200) );
INVx1_ASAP7_75t_L g516 ( .A(n_33), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_33), .B(n_936), .Y(n_935) );
OAI21x1_ASAP7_75t_L g123 ( .A1(n_34), .A2(n_66), .B(n_124), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_35), .A2(n_133), .B(n_263), .C(n_264), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_37), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_38), .B(n_138), .Y(n_157) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_39), .B(n_177), .Y(n_183) );
AND2x6_ASAP7_75t_L g144 ( .A(n_40), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g596 ( .A(n_41), .B(n_168), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_42), .B(n_168), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_43), .A2(n_53), .B1(n_905), .B2(n_906), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_43), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_44), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_45), .B(n_244), .Y(n_243) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_46), .B(n_177), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_47), .B(n_128), .Y(n_620) );
INVx1_ASAP7_75t_L g145 ( .A(n_48), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_49), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_51), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_52), .B(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g906 ( .A(n_53), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_54), .A2(n_105), .B1(n_929), .B2(n_940), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_55), .B(n_168), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_56), .B(n_140), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_57), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_58), .B(n_140), .Y(n_664) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_59), .Y(n_520) );
NAND2x1_ASAP7_75t_L g625 ( .A(n_59), .B(n_168), .Y(n_625) );
AND2x2_ASAP7_75t_L g266 ( .A(n_60), .B(n_147), .Y(n_266) );
AND2x2_ASAP7_75t_L g937 ( .A(n_61), .B(n_938), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_62), .B(n_141), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_64), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_65), .B(n_658), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_67), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_68), .Y(n_661) );
NAND2xp33_ASAP7_75t_L g127 ( .A(n_69), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_70), .B(n_141), .Y(n_636) );
OAI22xp5_ASAP7_75t_SL g908 ( .A1(n_71), .A2(n_102), .B1(n_909), .B2(n_910), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_71), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_72), .A2(n_77), .B1(n_140), .B2(n_572), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_73), .B(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_74), .A2(n_520), .B1(n_521), .B2(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_74), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_75), .Y(n_564) );
BUFx10_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_78), .B(n_156), .Y(n_241) );
INVx1_ASAP7_75t_SL g587 ( .A(n_79), .Y(n_587) );
NAND2xp33_ASAP7_75t_L g139 ( .A(n_80), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_81), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_82), .B(n_197), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_83), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_85), .Y(n_265) );
AND2x2_ASAP7_75t_L g933 ( .A(n_86), .B(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_88), .B(n_141), .Y(n_609) );
OR2x2_ASAP7_75t_L g513 ( .A(n_89), .B(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g540 ( .A(n_89), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_89), .B(n_515), .Y(n_928) );
INVx1_ASAP7_75t_L g939 ( .A(n_89), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_90), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_91), .B(n_177), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_92), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_93), .B(n_168), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_94), .Y(n_209) );
INVx1_ASAP7_75t_L g938 ( .A(n_95), .Y(n_938) );
INVx1_ASAP7_75t_L g256 ( .A(n_96), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_97), .Y(n_225) );
AND2x2_ASAP7_75t_L g235 ( .A(n_98), .B(n_121), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_99), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_100), .B(n_232), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_101), .B(n_147), .Y(n_146) );
INVxp67_ASAP7_75t_L g910 ( .A(n_102), .Y(n_910) );
AO22x1_ASAP7_75t_L g505 ( .A1(n_103), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_103), .Y(n_508) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_532), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx12f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_L g538 ( .A(n_110), .Y(n_538) );
INVx2_ASAP7_75t_SL g927 ( .A(n_110), .Y(n_927) );
OAI21xp33_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_518), .B(n_523), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_510), .Y(n_112) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_113), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_505), .B(n_509), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp33_ASAP7_75t_L g509 ( .A(n_115), .B(n_505), .Y(n_509) );
INVx2_ASAP7_75t_L g921 ( .A(n_115), .Y(n_921) );
NAND4xp75_ASAP7_75t_L g115 ( .A(n_116), .B(n_361), .C(n_426), .D(n_476), .Y(n_115) );
NOR3x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_292), .C(n_329), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_186), .B(n_202), .C(n_267), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_118), .A2(n_307), .B(n_494), .Y(n_493) );
OR2x6_ASAP7_75t_SL g118 ( .A(n_119), .B(n_149), .Y(n_118) );
AND2x2_ASAP7_75t_L g379 ( .A(n_119), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g383 ( .A(n_119), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2x1_ASAP7_75t_L g390 ( .A(n_120), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_120), .Y(n_458) );
INVx2_ASAP7_75t_L g474 ( .A(n_120), .Y(n_474) );
OA21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_146), .Y(n_120) );
BUFx4f_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
INVx3_ASAP7_75t_L g173 ( .A(n_121), .Y(n_173) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_121), .A2(n_125), .B(n_146), .Y(n_188) );
INVx4_ASAP7_75t_L g219 ( .A(n_121), .Y(n_219) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_121), .A2(n_125), .B(n_146), .Y(n_283) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_121), .Y(n_645) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g169 ( .A(n_122), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_122), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_135), .B(n_142), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B(n_132), .Y(n_126) );
INVx2_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
INVx1_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
INVx2_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
INVx2_ASAP7_75t_L g555 ( .A(n_128), .Y(n_555) );
INVx2_ASAP7_75t_L g562 ( .A(n_128), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_128), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g622 ( .A(n_128), .Y(n_622) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_129), .Y(n_138) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
INVx2_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_129), .Y(n_232) );
INVx1_ASAP7_75t_L g260 ( .A(n_129), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_132), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_132), .A2(n_213), .B(n_214), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_132), .A2(n_234), .B1(n_571), .B2(n_573), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_132), .A2(n_165), .B1(n_583), .B2(n_584), .Y(n_582) );
OA22x2_ASAP7_75t_L g592 ( .A1(n_132), .A2(n_165), .B1(n_593), .B2(n_594), .Y(n_592) );
CKINVDCx6p67_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_SL g226 ( .A(n_133), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_133), .A2(n_558), .B(n_563), .Y(n_557) );
AOI21x1_ASAP7_75t_L g616 ( .A1(n_133), .A2(n_617), .B(n_618), .Y(n_616) );
AOI21x1_ASAP7_75t_L g632 ( .A1(n_133), .A2(n_633), .B(n_634), .Y(n_632) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx5_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_134), .A2(n_154), .B(n_155), .C(n_157), .Y(n_153) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
OAI321xp33_ASAP7_75t_L g552 ( .A1(n_134), .A2(n_140), .A3(n_553), .B1(n_554), .B2(n_555), .C(n_556), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_134), .A2(n_636), .B1(n_637), .B2(n_638), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B(n_141), .Y(n_135) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_137), .B(n_225), .Y(n_224) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g161 ( .A(n_140), .Y(n_161) );
INVx2_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_140), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_SL g244 ( .A(n_140), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_140), .A2(n_141), .B(n_661), .C(n_662), .Y(n_660) );
AOI21x1_ASAP7_75t_L g175 ( .A1(n_141), .A2(n_176), .B(n_178), .Y(n_175) );
INVx1_ASAP7_75t_L g246 ( .A(n_141), .Y(n_246) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_142), .A2(n_153), .B(n_158), .Y(n_152) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_142), .A2(n_194), .B(n_198), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_142), .A2(n_208), .B(n_212), .Y(n_207) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_142), .A2(n_239), .B(n_242), .Y(n_238) );
AND2x2_ASAP7_75t_L g569 ( .A(n_142), .B(n_173), .Y(n_569) );
AO31x2_ASAP7_75t_L g581 ( .A1(n_142), .A2(n_219), .A3(n_582), .B(n_586), .Y(n_581) );
INVx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_143), .A2(n_221), .B(n_227), .Y(n_220) );
NOR2xp67_ASAP7_75t_L g251 ( .A(n_143), .B(n_252), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_143), .A2(n_556), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g591 ( .A(n_143), .Y(n_591) );
INVx8_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx2_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_144), .A2(n_603), .B(n_608), .Y(n_602) );
OAI21x1_ASAP7_75t_L g631 ( .A1(n_144), .A2(n_632), .B(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g668 ( .A(n_144), .Y(n_668) );
INVx2_ASAP7_75t_L g590 ( .A(n_147), .Y(n_590) );
BUFx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_148), .Y(n_566) );
INVx1_ASAP7_75t_L g576 ( .A(n_148), .Y(n_576) );
INVx2_ASAP7_75t_L g337 ( .A(n_149), .Y(n_337) );
OR2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_170), .Y(n_149) );
AND2x2_ASAP7_75t_L g271 ( .A(n_150), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g386 ( .A(n_150), .Y(n_386) );
AND2x2_ASAP7_75t_L g393 ( .A(n_150), .B(n_275), .Y(n_393) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_167), .Y(n_150) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_151), .A2(n_193), .B(n_201), .Y(n_192) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_151), .A2(n_207), .B(n_215), .Y(n_206) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_151), .A2(n_152), .B(n_167), .Y(n_279) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_151), .A2(n_193), .B(n_201), .Y(n_285) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .C(n_165), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g198 ( .A1(n_160), .A2(n_165), .B(n_199), .C(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g177 ( .A(n_164), .Y(n_177) );
INVx2_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_L g208 ( .A1(n_165), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_166), .A2(n_181), .B(n_183), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_166), .Y(n_234) );
BUFx2_ASAP7_75t_L g261 ( .A(n_166), .Y(n_261) );
AOI21x1_ASAP7_75t_L g619 ( .A1(n_166), .A2(n_620), .B(n_621), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_166), .A2(n_664), .B(n_665), .Y(n_663) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g190 ( .A(n_170), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g306 ( .A(n_170), .Y(n_306) );
AND2x2_ASAP7_75t_L g355 ( .A(n_170), .B(n_192), .Y(n_355) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_185), .Y(n_171) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_172), .A2(n_238), .B(n_247), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_172), .A2(n_174), .B(n_185), .Y(n_272) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_172), .A2(n_602), .B(n_611), .Y(n_601) );
OAI21x1_ASAP7_75t_L g649 ( .A1(n_172), .A2(n_602), .B(n_611), .Y(n_649) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_180), .B(n_184), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_177), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g210 ( .A(n_179), .Y(n_210) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_184), .A2(n_616), .B(n_619), .Y(n_615) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
OR2x2_ASAP7_75t_L g346 ( .A(n_187), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g398 ( .A(n_187), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g408 ( .A(n_187), .B(n_402), .Y(n_408) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_SL g274 ( .A(n_188), .Y(n_274) );
BUFx2_ASAP7_75t_L g319 ( .A(n_188), .Y(n_319) );
INVx1_ASAP7_75t_SL g437 ( .A(n_188), .Y(n_437) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g317 ( .A(n_190), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g468 ( .A(n_190), .B(n_353), .Y(n_468) );
INVx2_ASAP7_75t_L g275 ( .A(n_191), .Y(n_275) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_197), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI221xp5_ASAP7_75t_SL g459 ( .A1(n_203), .A2(n_460), .B1(n_463), .B2(n_465), .C(n_466), .Y(n_459) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_216), .Y(n_203) );
INVxp67_ASAP7_75t_L g394 ( .A(n_204), .Y(n_394) );
AND2x4_ASAP7_75t_L g397 ( .A(n_204), .B(n_374), .Y(n_397) );
OR2x2_ASAP7_75t_L g419 ( .A(n_204), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_205), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g359 ( .A(n_205), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_205), .B(n_314), .Y(n_376) );
AND2x2_ASAP7_75t_L g387 ( .A(n_205), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_205), .B(n_374), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_205), .B(n_217), .Y(n_456) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
AND2x2_ASAP7_75t_L g471 ( .A(n_206), .B(n_297), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_216), .A2(n_352), .B1(n_379), .B2(n_381), .Y(n_378) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_236), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_217), .B(n_299), .Y(n_484) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_SL g328 ( .A(n_218), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_218), .B(n_335), .Y(n_334) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_235), .Y(n_218) );
INVx3_ASAP7_75t_L g252 ( .A(n_219), .Y(n_252) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_219), .A2(n_220), .B(n_235), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_226), .Y(n_221) );
OAI21xp33_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_230), .B(n_234), .Y(n_227) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_231), .B(n_233), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_231), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g572 ( .A(n_232), .Y(n_572) );
INVx2_ASAP7_75t_L g606 ( .A(n_232), .Y(n_606) );
INVx2_ASAP7_75t_L g666 ( .A(n_232), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_234), .A2(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g457 ( .A(n_236), .Y(n_457) );
AND2x4_ASAP7_75t_L g470 ( .A(n_236), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_248), .Y(n_236) );
AND2x2_ASAP7_75t_L g287 ( .A(n_237), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
OR2x2_ASAP7_75t_L g310 ( .A(n_237), .B(n_297), .Y(n_310) );
INVx1_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_237), .Y(n_360) );
INVx1_ASAP7_75t_L g388 ( .A(n_237), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B(n_246), .Y(n_242) );
INVx2_ASAP7_75t_L g263 ( .A(n_244), .Y(n_263) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g291 ( .A(n_249), .Y(n_291) );
AND2x2_ASAP7_75t_L g296 ( .A(n_249), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g369 ( .A(n_249), .B(n_328), .Y(n_369) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g314 ( .A(n_250), .Y(n_314) );
AOI21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B(n_266), .Y(n_250) );
OAI21x1_ASAP7_75t_L g614 ( .A1(n_252), .A2(n_615), .B(n_625), .Y(n_614) );
OAI21x1_ASAP7_75t_L g630 ( .A1(n_252), .A2(n_631), .B(n_639), .Y(n_630) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_252), .A2(n_615), .B(n_625), .Y(n_677) );
OAI21x1_ASAP7_75t_L g702 ( .A1(n_252), .A2(n_631), .B(n_639), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_262), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_257), .B(n_261), .Y(n_254) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g585 ( .A(n_260), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_263), .A2(n_609), .B(n_610), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_276), .B(n_286), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_273), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NOR2x1_ASAP7_75t_SL g366 ( .A(n_270), .B(n_273), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_270), .A2(n_453), .B(n_455), .C(n_458), .Y(n_452) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g340 ( .A(n_271), .Y(n_340) );
BUFx2_ASAP7_75t_L g487 ( .A(n_272), .Y(n_487) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_273), .Y(n_315) );
INVx1_ASAP7_75t_L g431 ( .A(n_273), .Y(n_431) );
OR2x2_ASAP7_75t_L g446 ( .A(n_273), .B(n_447), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_273), .A2(n_470), .B(n_487), .C(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_274), .B(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g303 ( .A(n_275), .B(n_283), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_275), .B(n_306), .Y(n_323) );
INVx1_ASAP7_75t_L g348 ( .A(n_275), .Y(n_348) );
AND2x2_ASAP7_75t_L g497 ( .A(n_275), .B(n_283), .Y(n_497) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
AND2x2_ASAP7_75t_L g496 ( .A(n_277), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_SL g304 ( .A(n_278), .B(n_305), .Y(n_304) );
NAND2x1_ASAP7_75t_L g347 ( .A(n_278), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_278), .B(n_284), .Y(n_399) );
BUFx2_ASAP7_75t_L g461 ( .A(n_278), .Y(n_461) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_279), .Y(n_322) );
INVx1_ASAP7_75t_L g354 ( .A(n_279), .Y(n_354) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_280), .Y(n_336) );
AND2x2_ASAP7_75t_L g491 ( .A(n_280), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_283), .B(n_386), .Y(n_418) );
INVx1_ASAP7_75t_L g339 ( .A(n_284), .Y(n_339) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g380 ( .A(n_285), .B(n_306), .Y(n_380) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
AND2x2_ASAP7_75t_L g324 ( .A(n_287), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g344 ( .A(n_287), .B(n_296), .Y(n_344) );
AND2x4_ASAP7_75t_L g368 ( .A(n_287), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_287), .B(n_357), .Y(n_479) );
OR2x2_ASAP7_75t_L g299 ( .A(n_288), .B(n_300), .Y(n_299) );
BUFx3_ASAP7_75t_L g425 ( .A(n_288), .Y(n_425) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g342 ( .A(n_290), .B(n_310), .Y(n_342) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g421 ( .A(n_291), .B(n_297), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_301), .B1(n_307), .B2(n_315), .C(n_316), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_294), .A2(n_484), .B(n_495), .C(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_295), .A2(n_467), .B1(n_469), .B2(n_472), .Y(n_466) );
OR2x2_ASAP7_75t_L g504 ( .A(n_295), .B(n_359), .Y(n_504) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g412 ( .A(n_296), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_296), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_298), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g413 ( .A(n_299), .Y(n_413) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_299), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
AND2x4_ASAP7_75t_L g433 ( .A(n_302), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g462 ( .A(n_303), .Y(n_462) );
INVx1_ASAP7_75t_L g392 ( .A(n_305), .Y(n_392) );
AND2x4_ASAP7_75t_L g438 ( .A(n_305), .B(n_353), .Y(n_438) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g374 ( .A(n_310), .Y(n_374) );
OR2x2_ASAP7_75t_L g451 ( .A(n_310), .B(n_332), .Y(n_451) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g488 ( .A(n_312), .B(n_334), .Y(n_488) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g332 ( .A(n_314), .Y(n_332) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_314), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B(n_324), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g411 ( .A(n_319), .B(n_355), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_320), .A2(n_445), .B1(n_448), .B2(n_450), .C(n_452), .Y(n_444) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_322), .Y(n_434) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_322), .Y(n_447) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g404 ( .A(n_326), .Y(n_404) );
AOI322xp5_ASAP7_75t_L g428 ( .A1(n_326), .A2(n_344), .A3(n_429), .B1(n_432), .B2(n_433), .C1(n_435), .C2(n_439), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_326), .B(n_387), .Y(n_464) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_343), .C(n_349), .Y(n_329) );
AOI32xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .A3(n_337), .B1(n_338), .B2(n_341), .Y(n_330) );
OAI21xp33_ASAP7_75t_SL g343 ( .A1(n_331), .A2(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g454 ( .A(n_332), .Y(n_454) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g449 ( .A(n_334), .B(n_376), .Y(n_449) );
NAND2x1_ASAP7_75t_SL g430 ( .A(n_337), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g485 ( .A(n_339), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g409 ( .A(n_340), .Y(n_409) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g381 ( .A(n_342), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_344), .A2(n_433), .B1(n_438), .B2(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g465 ( .A(n_347), .Y(n_465) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp67_ASAP7_75t_SL g350 ( .A(n_351), .B(n_356), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g480 ( .A(n_352), .B(n_458), .Y(n_480) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx2_ASAP7_75t_L g492 ( .A(n_353), .Y(n_492) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_355), .B(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g475 ( .A(n_355), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_356), .A2(n_410), .B1(n_467), .B2(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_382), .C(n_405), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_377), .Y(n_363) );
OAI21xp33_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_367), .B(n_370), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x2_ASAP7_75t_L g416 ( .A(n_371), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g489 ( .A(n_371), .Y(n_489) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g402 ( .A(n_380), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_387), .B(n_389), .Y(n_382) );
INVx1_ASAP7_75t_L g401 ( .A(n_385), .Y(n_401) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_387), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g495 ( .A(n_387), .Y(n_495) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_394), .A3(n_395), .B1(n_396), .B2(n_398), .C1(n_400), .C2(n_403), .Y(n_389) );
INVx1_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g407 ( .A(n_393), .Y(n_407) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g501 ( .A(n_398), .Y(n_501) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_412), .B(n_414), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .C(n_409), .D(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_419), .B1(n_422), .B2(n_423), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g442 ( .A(n_421), .B(n_424), .Y(n_442) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g473 ( .A(n_425), .B(n_474), .Y(n_473) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_443), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_441), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_459), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g502 ( .A(n_453), .Y(n_502) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
NAND2xp33_ASAP7_75t_SL g472 ( .A(n_473), .B(n_475), .Y(n_472) );
AND3x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .C(n_498), .Y(n_476) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_SL g481 ( .A(n_482), .B(n_493), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B1(n_488), .B2(n_489), .C(n_490), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g500 ( .A(n_486), .Y(n_500) );
INVx2_ASAP7_75t_L g499 ( .A(n_488), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_501), .B2(n_502), .C(n_503), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx5_ASAP7_75t_L g531 ( .A(n_511), .Y(n_531) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_512), .Y(n_528) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g539 ( .A(n_514), .B(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g916 ( .A(n_514), .B(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_519), .B(n_526), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_520), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_529), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp67_ASAP7_75t_R g529 ( .A(n_530), .B(n_531), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_541), .B1(n_913), .B2(n_918), .C(n_923), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x6_ASAP7_75t_SL g915 ( .A(n_537), .B(n_916), .Y(n_915) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_540), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_908), .B1(n_911), .B2(n_912), .Y(n_541) );
INVx2_ASAP7_75t_L g911 ( .A(n_542), .Y(n_911) );
OA22x2_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_903), .B1(n_904), .B2(n_907), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVxp67_ASAP7_75t_L g907 ( .A(n_544), .Y(n_907) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_794), .Y(n_544) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_546), .B(n_696), .C(n_733), .D(n_767), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_650), .Y(n_546) );
OAI32xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_577), .A3(n_597), .B1(n_626), .B2(n_642), .Y(n_547) );
OAI222xp33_ASAP7_75t_L g833 ( .A1(n_548), .A2(n_834), .B1(n_837), .B2(n_840), .C1(n_841), .C2(n_843), .Y(n_833) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_549), .B(n_847), .Y(n_846) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g752 ( .A(n_550), .Y(n_752) );
AND2x2_ASAP7_75t_L g766 ( .A(n_550), .B(n_738), .Y(n_766) );
AND2x2_ASAP7_75t_L g774 ( .A(n_550), .B(n_765), .Y(n_774) );
AND2x2_ASAP7_75t_L g901 ( .A(n_550), .B(n_739), .Y(n_901) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_567), .Y(n_550) );
INVx1_ASAP7_75t_L g681 ( .A(n_551), .Y(n_681) );
INVx2_ASAP7_75t_L g701 ( .A(n_551), .Y(n_701) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_557), .B(n_565), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g641 ( .A(n_567), .B(n_613), .Y(n_641) );
INVx2_ASAP7_75t_L g678 ( .A(n_567), .Y(n_678) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_567), .Y(n_771) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g695 ( .A(n_568), .Y(n_695) );
AOI21x1_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_574), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_576), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g658 ( .A(n_576), .Y(n_658) );
OAI332xp33_ASAP7_75t_L g858 ( .A1(n_577), .A2(n_648), .A3(n_859), .B1(n_860), .B2(n_861), .B3(n_863), .C1(n_865), .C2(n_867), .Y(n_858) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g777 ( .A(n_579), .B(n_778), .Y(n_777) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g689 ( .A(n_580), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_580), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_588), .Y(n_580) );
AND2x2_ASAP7_75t_L g643 ( .A(n_581), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g672 ( .A(n_581), .Y(n_672) );
INVx1_ASAP7_75t_L g687 ( .A(n_581), .Y(n_687) );
INVx1_ASAP7_75t_L g706 ( .A(n_581), .Y(n_706) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_581), .Y(n_732) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_588), .Y(n_711) );
INVx1_ASAP7_75t_L g792 ( .A(n_588), .Y(n_792) );
INVx1_ASAP7_75t_L g813 ( .A(n_588), .Y(n_813) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_588), .Y(n_850) );
INVx1_ASAP7_75t_L g878 ( .A(n_588), .Y(n_878) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B(n_595), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OA21x2_ASAP7_75t_L g644 ( .A1(n_592), .A2(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g646 ( .A(n_596), .Y(n_646) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_612), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_599), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_600), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g778 ( .A(n_600), .B(n_654), .Y(n_778) );
AND2x2_ASAP7_75t_L g857 ( .A(n_600), .B(n_672), .Y(n_857) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g836 ( .A(n_601), .B(n_644), .Y(n_836) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_607), .Y(n_603) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g682 ( .A(n_612), .Y(n_682) );
BUFx2_ASAP7_75t_L g742 ( .A(n_612), .Y(n_742) );
OR2x2_ASAP7_75t_L g750 ( .A(n_612), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_613), .Y(n_830) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g755 ( .A(n_614), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g637 ( .A(n_622), .Y(n_637) );
INVx4_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g734 ( .A(n_626), .B(n_735), .C(n_740), .Y(n_734) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_640), .Y(n_627) );
AND2x2_ASAP7_75t_L g864 ( .A(n_628), .B(n_799), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_628), .B(n_675), .Y(n_872) );
AND2x4_ASAP7_75t_L g885 ( .A(n_628), .B(n_785), .Y(n_885) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g751 ( .A(n_629), .Y(n_751) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g693 ( .A(n_630), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_640), .B(n_720), .Y(n_840) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g775 ( .A(n_641), .B(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
AND2x2_ASAP7_75t_L g748 ( .A(n_643), .B(n_648), .Y(n_748) );
AND2x2_ASAP7_75t_L g653 ( .A(n_644), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_647), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g802 ( .A(n_647), .B(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g831 ( .A(n_647), .B(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp67_ASAP7_75t_L g669 ( .A(n_648), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_648), .B(n_687), .Y(n_686) );
BUFx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g709 ( .A(n_649), .B(n_656), .Y(n_709) );
AND2x2_ASAP7_75t_L g758 ( .A(n_649), .B(n_655), .Y(n_758) );
OAI322xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_673), .A3(n_679), .B1(n_682), .B2(n_683), .C1(n_688), .C2(n_690), .Y(n_650) );
AOI21xp5_ASAP7_75t_SL g712 ( .A1(n_651), .A2(n_713), .B(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_652), .A2(n_768), .B1(n_777), .B2(n_779), .C(n_783), .Y(n_767) );
AND2x4_ASAP7_75t_L g652 ( .A(n_653), .B(n_669), .Y(n_652) );
INVx2_ASAP7_75t_L g685 ( .A(n_653), .Y(n_685) );
AND2x2_ASAP7_75t_L g856 ( .A(n_653), .B(n_857), .Y(n_856) );
AND2x2_ASAP7_75t_L g811 ( .A(n_654), .B(n_706), .Y(n_811) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g716 ( .A(n_656), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_667), .Y(n_659) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g793 ( .A(n_671), .B(n_716), .Y(n_793) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g803 ( .A(n_672), .B(n_716), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_673), .A2(n_884), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g699 ( .A(n_674), .Y(n_699) );
OR2x2_ASAP7_75t_L g822 ( .A(n_674), .B(n_789), .Y(n_822) );
AND2x2_ASAP7_75t_L g894 ( .A(n_674), .B(n_700), .Y(n_894) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx2_ASAP7_75t_L g780 ( .A(n_676), .Y(n_780) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g816 ( .A(n_677), .B(n_681), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_678), .B(n_693), .Y(n_741) );
INVx1_ASAP7_75t_L g786 ( .A(n_678), .Y(n_786) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_678), .Y(n_815) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g737 ( .A(n_680), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g694 ( .A(n_681), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_681), .B(n_755), .Y(n_772) );
OR2x2_ASAP7_75t_L g723 ( .A(n_682), .B(n_721), .Y(n_723) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2x1p5_ASAP7_75t_SL g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_687), .B(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_687), .Y(n_866) );
AND2x2_ASAP7_75t_L g743 ( .A(n_689), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx2_ASAP7_75t_L g720 ( .A(n_692), .Y(n_720) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g826 ( .A(n_694), .B(n_798), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_694), .B(n_864), .Y(n_863) );
OR2x2_ASAP7_75t_L g721 ( .A(n_695), .B(n_701), .Y(n_721) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_695), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_695), .B(n_739), .Y(n_782) );
AOI211xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_703), .B(n_712), .C(n_722), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_700), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g808 ( .A(n_700), .Y(n_808) );
AND2x2_ASAP7_75t_L g883 ( .A(n_700), .B(n_815), .Y(n_883) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g726 ( .A(n_701), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g776 ( .A(n_701), .B(n_751), .Y(n_776) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_701), .Y(n_869) );
INVx1_ASAP7_75t_L g727 ( .A(n_702), .Y(n_727) );
INVx2_ASAP7_75t_L g739 ( .A(n_702), .Y(n_739) );
AND2x4_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .Y(n_703) );
OAI322xp33_ASAP7_75t_L g817 ( .A1(n_704), .A2(n_818), .A3(n_822), .B1(n_823), .B2(n_827), .C1(n_828), .C2(n_831), .Y(n_817) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_705), .B(n_820), .Y(n_827) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g762 ( .A(n_707), .Y(n_762) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g730 ( .A(n_709), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g745 ( .A(n_709), .Y(n_745) );
AND2x2_ASAP7_75t_L g884 ( .A(n_709), .B(n_878), .Y(n_884) );
INVx1_ASAP7_75t_L g759 ( .A(n_710), .Y(n_759) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g842 ( .A(n_715), .Y(n_842) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g805 ( .A(n_720), .B(n_806), .Y(n_805) );
OR2x2_ASAP7_75t_L g854 ( .A(n_721), .B(n_780), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B(n_729), .Y(n_722) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_724), .A2(n_877), .B1(n_879), .B2(n_881), .C(n_882), .Y(n_876) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVx2_ASAP7_75t_L g789 ( .A(n_726), .Y(n_789) );
AND2x2_ASAP7_75t_L g855 ( .A(n_726), .B(n_799), .Y(n_855) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI211x1_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_743), .B(n_746), .C(n_760), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g829 ( .A(n_737), .B(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
O2A1O1Ixp33_ASAP7_75t_SL g783 ( .A1(n_740), .A2(n_784), .B(n_787), .C(n_790), .Y(n_783) );
OR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_741), .B(n_869), .Y(n_868) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_741), .Y(n_892) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B1(n_753), .B2(n_756), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
AND2x2_ASAP7_75t_L g824 ( .A(n_751), .B(n_825), .Y(n_824) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
BUFx2_ASAP7_75t_L g765 ( .A(n_755), .Y(n_765) );
AND2x2_ASAP7_75t_L g825 ( .A(n_755), .B(n_786), .Y(n_825) );
INVx1_ASAP7_75t_L g801 ( .A(n_756), .Y(n_801) );
OR2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g859 ( .A(n_757), .Y(n_859) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g839 ( .A(n_758), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_759), .B(n_842), .Y(n_841) );
NOR2xp67_ASAP7_75t_SL g760 ( .A(n_761), .B(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVxp67_ASAP7_75t_L g902 ( .A(n_765), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_766), .A2(n_810), .B1(n_812), .B2(n_814), .Y(n_809) );
INVx2_ASAP7_75t_SL g843 ( .A(n_766), .Y(n_843) );
NAND3xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_773), .C(n_775), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g806 ( .A(n_771), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_773), .A2(n_841), .B1(n_871), .B2(n_873), .Y(n_870) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI21xp33_ASAP7_75t_SL g804 ( .A1(n_777), .A2(n_805), .B(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g821 ( .A(n_778), .Y(n_821) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
AND2x2_ASAP7_75t_L g785 ( .A(n_780), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g799 ( .A(n_780), .Y(n_799) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
OR2x2_ASAP7_75t_L g797 ( .A(n_782), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
AND2x2_ASAP7_75t_L g810 ( .A(n_792), .B(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g862 ( .A(n_792), .Y(n_862) );
AND2x4_ASAP7_75t_L g835 ( .A(n_793), .B(n_836), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_844), .C(n_875), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_817), .C(n_833), .Y(n_795) );
OAI211xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_800), .B(n_804), .C(n_809), .Y(n_796) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
AND2x2_ASAP7_75t_L g812 ( .A(n_803), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g832 ( .A(n_803), .Y(n_832) );
INVx2_ASAP7_75t_L g851 ( .A(n_803), .Y(n_851) );
BUFx2_ASAP7_75t_L g896 ( .A(n_803), .Y(n_896) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_812), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g889 ( .A(n_816), .Y(n_889) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_820), .B(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_SL g823 ( .A(n_824), .B(n_826), .Y(n_823) );
INVx1_ASAP7_75t_L g860 ( .A(n_824), .Y(n_860) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g880 ( .A(n_832), .Y(n_880) );
OAI211xp5_ASAP7_75t_L g886 ( .A1(n_834), .A2(n_887), .B(n_890), .C(n_893), .Y(n_886) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_836), .B(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g895 ( .A(n_836), .B(n_896), .Y(n_895) );
INVxp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g874 ( .A(n_838), .B(n_862), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_858), .C(n_870), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_852), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
OR2x6_ASAP7_75t_L g877 ( .A(n_851), .B(n_878), .Y(n_877) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_855), .B(n_856), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g881 ( .A(n_855), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_856), .B(n_891), .Y(n_890) );
INVxp67_ASAP7_75t_L g898 ( .A(n_859), .Y(n_898) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NOR3xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_886), .C(n_897), .Y(n_875) );
INVxp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
AO22x2_ASAP7_75t_L g920 ( .A1(n_903), .A2(n_904), .B1(n_921), .B2(n_922), .Y(n_920) );
INVxp33_ASAP7_75t_SL g903 ( .A(n_904), .Y(n_903) );
INVxp33_ASAP7_75t_SL g912 ( .A(n_908), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_908), .A2(n_912), .B1(n_919), .B2(n_920), .Y(n_918) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
BUFx4_ASAP7_75t_SL g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_SL g922 ( .A(n_921), .Y(n_922) );
INVx5_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
BUFx12f_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
BUFx4f_ASAP7_75t_SL g929 ( .A(n_930), .Y(n_929) );
BUFx3_ASAP7_75t_L g941 ( .A(n_930), .Y(n_941) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx4_ASAP7_75t_SL g931 ( .A(n_932), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_933), .B(n_935), .Y(n_932) );
NAND2xp5_ASAP7_75t_SL g936 ( .A(n_937), .B(n_939), .Y(n_936) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
endmodule