module fake_jpeg_19556_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_16),
.B1(n_24),
.B2(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_49),
.B1(n_24),
.B2(n_18),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_16),
.B1(n_24),
.B2(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_18),
.B1(n_31),
.B2(n_20),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_19),
.C(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_40),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_35),
.B1(n_40),
.B2(n_39),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_71),
.B1(n_72),
.B2(n_77),
.Y(n_97)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_43),
.C(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_39),
.B1(n_34),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_55),
.B1(n_51),
.B2(n_52),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_23),
.B(n_25),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_74),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_31),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_33),
.B1(n_38),
.B2(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_22),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_78),
.A3(n_79),
.B1(n_59),
.B2(n_74),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_33),
.B1(n_38),
.B2(n_20),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_38),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_38),
.B(n_23),
.C(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_21),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_82),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_25),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_43),
.C(n_53),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_93),
.C(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_94),
.B1(n_79),
.B2(n_75),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_53),
.C(n_55),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_68),
.B1(n_67),
.B2(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_46),
.B1(n_21),
.B2(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_29),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_63),
.B1(n_81),
.B2(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_112),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_70),
.B1(n_79),
.B2(n_75),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_132),
.B1(n_91),
.B2(n_94),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_123),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_88),
.B1(n_85),
.B2(n_17),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_122),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_61),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_87),
.B(n_92),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_32),
.C(n_28),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_109),
.C(n_112),
.Y(n_148)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_129),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_1),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_139),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_161),
.B1(n_5),
.B2(n_7),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_142),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_108),
.B1(n_100),
.B2(n_92),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_147),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_102),
.C(n_92),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_1),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_121),
.C(n_101),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_125),
.C(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_97),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_160),
.A2(n_134),
.B(n_133),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_124),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_168),
.C(n_169),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_121),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_116),
.B(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_184),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_120),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_173),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_4),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_149),
.B(n_160),
.C(n_150),
.D(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_179),
.A2(n_152),
.B1(n_140),
.B2(n_9),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_7),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_194),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_145),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_189),
.B1(n_172),
.B2(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_139),
.B1(n_157),
.B2(n_156),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_142),
.B1(n_138),
.B2(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_153),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_152),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_169),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_208),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_178),
.B1(n_170),
.B2(n_179),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_162),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_192),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_193),
.C(n_177),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_164),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_173),
.C(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_186),
.B1(n_198),
.B2(n_195),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_198),
.B(n_188),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_223),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_189),
.C(n_184),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_212),
.C(n_213),
.Y(n_234)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_200),
.B1(n_211),
.B2(n_215),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_176),
.B1(n_217),
.B2(n_140),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_209),
.B(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_171),
.C(n_165),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_7),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_218),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_176),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_236),
.B1(n_230),
.B2(n_9),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_218),
.C(n_8),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_8),
.C(n_9),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.C(n_243),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_250),
.B1(n_246),
.B2(n_11),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_237),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_248),
.B(n_242),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_253),
.B(n_8),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_249),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_13),
.Y(n_257)
);


endmodule