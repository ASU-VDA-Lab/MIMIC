module fake_jpeg_2542_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_5),
.B(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_44),
.Y(n_68)
);

OR2x4_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_42),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_38),
.B1(n_36),
.B2(n_42),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_46),
.B1(n_41),
.B2(n_35),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_66),
.B(n_47),
.C(n_1),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_48),
.C(n_38),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_46),
.C(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_41),
.B1(n_35),
.B2(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_76),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_15),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_6),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_58),
.B(n_64),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_57),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_88),
.C(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_27),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_75),
.B1(n_69),
.B2(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_102),
.Y(n_111)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_101),
.C(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_103),
.Y(n_113)
);

NAND5xp2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_75),
.C(n_24),
.D(n_25),
.E(n_34),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_9),
.B(n_11),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_79),
.B1(n_88),
.B2(n_91),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_9),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_89),
.C(n_23),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_19),
.A3(n_30),
.B1(n_32),
.B2(n_33),
.C1(n_116),
.C2(n_113),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_99),
.A3(n_101),
.B1(n_14),
.B2(n_26),
.C1(n_28),
.C2(n_22),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.C(n_122),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_99),
.C(n_29),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_110),
.C(n_106),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_115),
.B(n_114),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_120),
.B(n_109),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_126),
.C(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_108),
.Y(n_131)
);


endmodule