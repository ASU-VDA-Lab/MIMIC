module fake_netlist_6_2472_n_108 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_108);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_108;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_1),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_31),
.B1(n_25),
.B2(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_42),
.Y(n_55)
);

OR2x6_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_R g57 ( 
.A(n_46),
.B(n_37),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_43),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_50),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_56),
.B(n_55),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_35),
.B1(n_37),
.B2(n_53),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_60),
.B1(n_68),
.B2(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_68),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_R g75 ( 
.A(n_73),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_76),
.B1(n_74),
.B2(n_47),
.C(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_53),
.B(n_67),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_14),
.Y(n_83)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_78),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OR2x6_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

O2A1O1Ixp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_40),
.B(n_80),
.C(n_47),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_41),
.B(n_39),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_84),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_88),
.Y(n_95)
);

OAI322xp33_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_84),
.A3(n_6),
.B1(n_8),
.B2(n_4),
.C1(n_39),
.C2(n_41),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_91),
.B1(n_90),
.B2(n_39),
.C(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_87),
.B1(n_83),
.B2(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_87),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_45),
.C(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_98),
.Y(n_102)
);

NOR4xp25_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_6),
.C(n_52),
.D(n_45),
.Y(n_103)
);

AND3x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_52),
.C(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

NOR2x1p5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_102),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_41),
.B(n_45),
.Y(n_108)
);


endmodule