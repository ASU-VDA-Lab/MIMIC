module fake_jpeg_3746_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_20),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_32),
.B1(n_24),
.B2(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_72),
.B1(n_24),
.B2(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_66),
.Y(n_82)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_60),
.B1(n_18),
.B2(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_84),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_32),
.B1(n_67),
.B2(n_40),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_44),
.C(n_37),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_90),
.C(n_20),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_94),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_98),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g98 ( 
.A(n_57),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_59),
.A2(n_46),
.B(n_43),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_28),
.B(n_19),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_108),
.B1(n_124),
.B2(n_83),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_23),
.B(n_29),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_27),
.Y(n_131)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_117),
.B1(n_118),
.B2(n_122),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_121),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_67),
.B1(n_59),
.B2(n_31),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_37),
.C(n_69),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_119),
.C(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_37),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_95),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_42),
.C(n_51),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_125),
.Y(n_147)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_128),
.B1(n_42),
.B2(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_96),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_74),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_87),
.B1(n_31),
.B2(n_83),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_142),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_147),
.C(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_79),
.B1(n_32),
.B2(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_150),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_34),
.B(n_28),
.C(n_19),
.D(n_22),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_23),
.B1(n_94),
.B2(n_25),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_110),
.B(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_172),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_179),
.B(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_171),
.Y(n_194)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_174),
.C(n_177),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_178),
.B(n_137),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_121),
.B1(n_128),
.B2(n_123),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_151),
.B1(n_146),
.B2(n_127),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_22),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_81),
.B(n_22),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_81),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_22),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_183),
.C(n_25),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_117),
.B(n_122),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_22),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_155),
.B1(n_137),
.B2(n_144),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_191),
.B1(n_200),
.B2(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_207),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_149),
.B(n_131),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_190),
.B(n_163),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_150),
.B1(n_132),
.B2(n_153),
.Y(n_191)
);

AOI21x1_ASAP7_75t_SL g195 ( 
.A1(n_159),
.A2(n_152),
.B(n_132),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_140),
.B1(n_109),
.B2(n_118),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_55),
.B1(n_50),
.B2(n_88),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_25),
.A3(n_34),
.B1(n_28),
.B2(n_50),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_183),
.C(n_176),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_165),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_218),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_188),
.B(n_208),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_174),
.CI(n_198),
.CON(n_243),
.SN(n_243)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_180),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_177),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_224),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_169),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_209),
.C(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_171),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_234),
.B(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_164),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_232),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_185),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_179),
.B1(n_34),
.B2(n_10),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_245),
.C(n_219),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_187),
.B1(n_196),
.B2(n_185),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_238),
.A2(n_247),
.B1(n_250),
.B2(n_255),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_198),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_216),
.A2(n_184),
.B1(n_200),
.B2(n_197),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_186),
.B1(n_191),
.B2(n_172),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_257),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_206),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_178),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_161),
.B1(n_204),
.B2(n_207),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_256),
.A2(n_223),
.B1(n_225),
.B2(n_222),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_230),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_211),
.A2(n_179),
.B1(n_9),
.B2(n_11),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_264),
.C(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_229),
.C(n_215),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_243),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_214),
.C(n_211),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_227),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_273),
.B(n_274),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_214),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_225),
.Y(n_273)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_277),
.B(n_1),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_241),
.C(n_245),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_292),
.C(n_293),
.Y(n_306)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_242),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_5),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_248),
.B1(n_222),
.B2(n_223),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_287),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_253),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_250),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_267),
.A2(n_255),
.B1(n_244),
.B2(n_256),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_226),
.C(n_2),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_1),
.C(n_2),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_6),
.B(n_7),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_302),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_272),
.CI(n_278),
.CON(n_297),
.SN(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_304),
.Y(n_313)
);

OAI31xp67_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_269),
.A3(n_275),
.B(n_3),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_299),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_4),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_7),
.C(n_8),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_305),
.B(n_293),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_280),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_11),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_286),
.B(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_314),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_279),
.B(n_8),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_297),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_7),
.C(n_9),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_12),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_307),
.B(n_302),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_322),
.B(n_325),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_327),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_12),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_309),
.B1(n_315),
.B2(n_14),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_332),
.Y(n_335)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_12),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_333),
.B(n_13),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_330),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_335),
.B1(n_328),
.B2(n_16),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_16),
.B(n_13),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_15),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_15),
.Y(n_340)
);


endmodule