module fake_jpeg_31417_n_172 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_53),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_16),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_32),
.B1(n_22),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_39),
.B1(n_35),
.B2(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_32),
.B1(n_18),
.B2(n_15),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_29),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_20),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_68),
.Y(n_89)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_73),
.B1(n_71),
.B2(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_84),
.B1(n_57),
.B2(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_36),
.B1(n_41),
.B2(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_58),
.B1(n_54),
.B2(n_63),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_42),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_15),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_19),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_48),
.B(n_52),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_105),
.B(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_87),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_68),
.B(n_64),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_47),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_98),
.C(n_94),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_82),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_19),
.B(n_28),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_114),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.C(n_88),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_89),
.C(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_120),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_94),
.B(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

OAI322xp33_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_116),
.A3(n_107),
.B1(n_70),
.B2(n_122),
.C1(n_19),
.C2(n_0),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_1),
.C(n_3),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_91),
.B(n_84),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_118),
.B1(n_109),
.B2(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_134),
.B1(n_121),
.B2(n_118),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_65),
.B1(n_80),
.B2(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_28),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_142),
.Y(n_149)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_125),
.A3(n_11),
.B1(n_13),
.B2(n_8),
.C(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_136),
.C(n_127),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_150),
.B(n_153),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_131),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_136),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_133),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_160),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_156),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_140),
.B1(n_152),
.B2(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_167),
.C(n_163),
.Y(n_169)
);

AOI31xp67_ASAP7_75t_SL g168 ( 
.A1(n_166),
.A2(n_162),
.A3(n_134),
.B(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);

O2A1O1Ixp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_159),
.B(n_155),
.C(n_137),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_13),
.Y(n_172)
);


endmodule