module fake_jpeg_18494_n_237 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_33),
.Y(n_61)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_29),
.Y(n_57)
);

NAND2x1p5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_22),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_34),
.B(n_38),
.C(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_48),
.B(n_15),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_32),
.B1(n_19),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_51),
.B1(n_53),
.B2(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_32),
.B1(n_18),
.B2(n_20),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_23),
.B1(n_19),
.B2(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_44),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_18),
.B1(n_30),
.B2(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_45),
.Y(n_86)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_23),
.B1(n_27),
.B2(n_16),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_38),
.B1(n_33),
.B2(n_28),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_98),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_42),
.B1(n_44),
.B2(n_38),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_97),
.B1(n_68),
.B2(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_28),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_45),
.B(n_44),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_28),
.B(n_25),
.C(n_4),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_99),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_55),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_15),
.C(n_2),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_1),
.C(n_3),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_17),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_72),
.B1(n_74),
.B2(n_52),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_132),
.B1(n_92),
.B2(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_7),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_70),
.C(n_65),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_67),
.C(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_75),
.B1(n_49),
.B2(n_56),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_118),
.B1(n_131),
.B2(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_67),
.B1(n_58),
.B2(n_33),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_124),
.Y(n_140)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_126),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_93),
.B(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_25),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_105),
.B1(n_80),
.B2(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_1),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_13),
.B1(n_8),
.B2(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_139),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_153),
.B(n_157),
.Y(n_159)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_96),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_144),
.C(n_125),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_109),
.B(n_91),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_152),
.C(n_131),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_116),
.B1(n_107),
.B2(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_82),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_114),
.B(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_169),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_171),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_124),
.B(n_118),
.C(n_109),
.D(n_113),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_142),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_122),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_110),
.B(n_106),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_176),
.B(n_147),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_106),
.C(n_88),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_137),
.C(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_129),
.B(n_102),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_173),
.C(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_161),
.A2(n_145),
.B1(n_140),
.B2(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_145),
.B1(n_156),
.B2(n_140),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_164),
.B1(n_172),
.B2(n_176),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_156),
.B1(n_158),
.B2(n_143),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_136),
.B(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_191),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_168),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_146),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_112),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_141),
.B(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_139),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_194),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_162),
.C(n_166),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_170),
.C(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_183),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_81),
.C(n_12),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_179),
.B1(n_186),
.B2(n_190),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_198),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_205),
.A2(n_187),
.B1(n_181),
.B2(n_191),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_192),
.B1(n_196),
.B2(n_195),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_200),
.B(n_202),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_184),
.B(n_193),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_193),
.B(n_201),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_222),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_210),
.C(n_216),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_221),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_211),
.B(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_227),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_212),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_213),
.B1(n_209),
.B2(n_210),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_225),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_232),
.A2(n_234),
.B(n_81),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_81),
.C(n_189),
.Y(n_233)
);

NAND2x1_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_12),
.Y(n_236)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);


endmodule