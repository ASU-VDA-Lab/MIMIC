module real_jpeg_16533_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_413),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_0),
.B(n_414),
.Y(n_413)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.A3(n_28),
.B1(n_34),
.B2(n_38),
.Y(n_24)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_1),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_1),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_37),
.B1(n_235),
.B2(n_239),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_3),
.A2(n_95),
.B1(n_123),
.B2(n_127),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_3),
.A2(n_95),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_95),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_4),
.Y(n_117)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_5),
.A2(n_277),
.B1(n_316),
.B2(n_409),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_6),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_8),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_9),
.A2(n_299),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_9),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g323 ( 
.A1(n_9),
.A2(n_303),
.B1(n_324),
.B2(n_327),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_10),
.Y(n_217)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_10),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_13),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_13),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_13),
.Y(n_257)
);

XOR2x2_ASAP7_75t_R g15 ( 
.A(n_16),
.B(n_392),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

AO221x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_282),
.B1(n_284),
.B2(n_385),
.C(n_391),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_222),
.B(n_281),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_199),
.B(n_221),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_149),
.B(n_198),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_131),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_22),
.B(n_131),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_65),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_23),
.B(n_98),
.C(n_129),
.Y(n_220)
);

XOR2x2_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_24),
.B(n_43),
.Y(n_202)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_26),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_108)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_33),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_33),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_36),
.A2(n_315),
.B1(n_317),
.B2(n_320),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_37),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_38),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_44),
.A2(n_135),
.B1(n_136),
.B2(n_143),
.Y(n_134)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_45),
.B(n_54),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_100),
.B(n_104),
.Y(n_99)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_49),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_49),
.Y(n_304)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_53),
.B(n_298),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_57),
.A2(n_104),
.A3(n_153),
.B1(n_157),
.B2(n_161),
.Y(n_152)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_61),
.Y(n_181)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_98),
.B1(n_129),
.B2(n_130),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_66),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_66),
.A2(n_129),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_66),
.B(n_287),
.C(n_288),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_66),
.A2(n_129),
.B1(n_287),
.B2(n_347),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_76),
.B1(n_83),
.B2(n_92),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_67),
.A2(n_76),
.B1(n_83),
.B2(n_92),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g358 ( 
.A1(n_67),
.A2(n_76),
.B(n_83),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_67),
.Y(n_406)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_72),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_72),
.B(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_74),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_212)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_75),
.Y(n_214)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_76),
.Y(n_407)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

OA22x2_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_SL g409 ( 
.A(n_93),
.Y(n_409)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_98),
.A2(n_130),
.B1(n_152),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_98),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_98),
.A2(n_130),
.B1(n_352),
.B2(n_378),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_107),
.B1(n_116),
.B2(n_122),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_107),
.B1(n_116),
.B2(n_122),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_99),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_99),
.B(n_230),
.Y(n_342)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_107),
.Y(n_230)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_107),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_110),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_118),
.Y(n_297)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_126),
.Y(n_330)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_129),
.B(n_228),
.C(n_232),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_147),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_132),
.A2(n_133),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_202),
.C(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_132),
.A2(n_133),
.B1(n_289),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_133),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_187),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_134),
.A2(n_168),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_135),
.A2(n_290),
.B1(n_298),
.B2(n_305),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_183),
.B(n_185),
.Y(n_182)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_142),
.Y(n_293)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_148),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.Y(n_405)
);

AOI21x1_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_171),
.B(n_197),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_167),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_SL g197 ( 
.A(n_151),
.B(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_168),
.B(n_262),
.Y(n_366)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_192),
.B(n_196),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_186),
.B(n_191),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_193),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_182),
.B(n_206),
.C(n_210),
.Y(n_259)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_185),
.A2(n_290),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_189),
.A2(n_313),
.B1(n_321),
.B2(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21x1_ASAP7_75t_SL g228 ( 
.A1(n_190),
.A2(n_229),
.B(n_231),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_190),
.A2(n_314),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_190),
.B(n_322),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_220),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_220),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_219),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_218),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_206),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_206),
.A2(n_312),
.B(n_331),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_206),
.B(n_312),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_206),
.B(n_287),
.C(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_206),
.A2(n_218),
.B1(n_287),
.B2(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_234),
.B1(n_242),
.B2(n_254),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_212),
.A2(n_243),
.B(n_249),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g287 ( 
.A1(n_212),
.A2(n_234),
.B1(n_242),
.B2(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_212),
.B(n_242),
.Y(n_337)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_224),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_258),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_225),
.B(n_259),
.C(n_260),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_232),
.Y(n_356)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_233),
.B(n_358),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_233),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_234),
.Y(n_336)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_272),
.B1(n_276),
.B2(n_277),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_369),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_359),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_343),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_285),
.B(n_343),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_310),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_286),
.B(n_311),
.C(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_287),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_332),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_323),
.B(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_331),
.A2(n_400),
.B1(n_401),
.B2(n_410),
.Y(n_399)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_332),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_340),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_338),
.B2(n_339),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_334),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_334),
.A2(n_338),
.B1(n_341),
.B2(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_334),
.A2(n_339),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_341),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_341),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_348),
.C(n_350),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_348),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.C(n_357),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_367),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_367),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.C(n_365),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_363),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_381),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_372),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_377),
.C(n_379),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_379),
.B2(n_380),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_384),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B(n_389),
.C(n_390),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_411),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_396),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);


endmodule