module fake_jpeg_25348_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_46),
.B1(n_49),
.B2(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_56),
.Y(n_67)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_36),
.B1(n_50),
.B2(n_47),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_66),
.B1(n_48),
.B2(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_4),
.Y(n_87)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_83),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_39),
.B1(n_43),
.B2(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_1),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_79),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_62),
.B(n_70),
.C(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_2),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_3),
.C(n_4),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_7),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_77),
.B1(n_79),
.B2(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_13),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_82),
.B1(n_74),
.B2(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_99),
.Y(n_109)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_88),
.B1(n_80),
.B2(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_93),
.B(n_96),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_110),
.B(n_14),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_88),
.C(n_91),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_15),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_114),
.A2(n_115),
.B(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_107),
.C(n_109),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_16),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_18),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_19),
.C(n_20),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_22),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_29),
.B(n_30),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_32),
.Y(n_123)
);


endmodule