module fake_jpeg_10498_n_123 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_20),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_18),
.Y(n_28)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_17),
.B1(n_16),
.B2(n_12),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_14),
.B1(n_12),
.B2(n_25),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_14),
.C(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_41),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_19),
.B(n_21),
.C(n_23),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_20),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_36),
.B1(n_43),
.B2(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_15),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_45),
.B(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_23),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_33),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI22x1_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_53),
.B1(n_37),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_21),
.B1(n_26),
.B2(n_20),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_28),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_40),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_55),
.C(n_51),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_8),
.Y(n_77)
);

XNOR2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_37),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_67),
.B(n_54),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_56),
.B(n_63),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_73),
.C(n_13),
.Y(n_85)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_74),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_13),
.B1(n_11),
.B2(n_22),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_77),
.B(n_13),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_8),
.C(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_22),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_35),
.C(n_22),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_78),
.B1(n_11),
.B2(n_35),
.Y(n_94)
);

OA21x2_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_72),
.B(n_71),
.Y(n_90)
);

OA21x2_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_82),
.B(n_83),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_95),
.C(n_96),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_35),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_35),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_84),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_105),
.C(n_98),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_91),
.C(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_104),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_82),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_104),
.B(n_99),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_108),
.B(n_5),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_110),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_96),
.C(n_1),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_4),
.C(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_2),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_5),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_3),
.C(n_4),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_115),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_112),
.B(n_7),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_3),
.B(n_4),
.C(n_7),
.D(n_8),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_9),
.B(n_0),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_120),
.B(n_9),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_118),
.B(n_9),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_0),
.Y(n_123)
);


endmodule