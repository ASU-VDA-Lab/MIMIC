module real_jpeg_19773_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_346, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_346;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_24),
.B1(n_26),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_0),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_0),
.A2(n_71),
.B1(n_72),
.B2(n_95),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_0),
.A2(n_53),
.B1(n_55),
.B2(n_95),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_95),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_1),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_1),
.A2(n_53),
.B1(n_55),
.B2(n_64),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_2),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_2),
.A2(n_23),
.B1(n_53),
.B2(n_55),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_36),
.B1(n_53),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_36),
.B1(n_71),
.B2(n_72),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_71),
.B1(n_72),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_53),
.B1(n_55),
.B2(n_131),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_131),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_131),
.Y(n_267)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_6),
.A2(n_55),
.B(n_67),
.C(n_111),
.D(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_6),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_6),
.B(n_52),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_6),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_6),
.A2(n_132),
.B(n_134),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_6),
.A2(n_33),
.B(n_49),
.C(n_170),
.D(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_33),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_37),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_150),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_32),
.B(n_34),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_24),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_62),
.B1(n_71),
.B2(n_72),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_7),
.A2(n_53),
.B1(n_55),
.B2(n_62),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_62),
.Y(n_283)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_8),
.A2(n_143),
.B1(n_180),
.B2(n_195),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_53),
.B1(n_55),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_10),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_114),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_114),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_53),
.B1(n_55),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_12),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_12),
.A2(n_71),
.B1(n_72),
.B2(n_126),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_126),
.Y(n_238)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_21),
.B(n_43),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_22),
.A2(n_27),
.B1(n_37),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_24),
.A2(n_29),
.B(n_150),
.C(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_35),
.B(n_37),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_27),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_28),
.A2(n_31),
.B1(n_238),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_28),
.A2(n_216),
.B(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_31),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_31),
.A2(n_94),
.B(n_239),
.Y(n_309)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_37),
.B(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21x1_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_81),
.B(n_343),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_76),
.C(n_78),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_45),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_59),
.C(n_65),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_47),
.B1(n_65),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_48),
.A2(n_57),
.B1(n_189),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_48),
.A2(n_211),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_52),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_49),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_49),
.A2(n_52),
.B1(n_264),
.B2(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_49),
.A2(n_52),
.B1(n_100),
.B2(n_283),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_51),
.Y(n_178)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_53),
.B(n_54),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_55),
.A2(n_170),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_57),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_57),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_57),
.A2(n_190),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_60),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_65),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B(n_75),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_66),
.A2(n_74),
.B1(n_125),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_66),
.A2(n_168),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_66),
.A2(n_74),
.B1(n_208),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_66),
.A2(n_74),
.B1(n_249),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_66),
.A2(n_74),
.B1(n_258),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_67),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_67),
.A2(n_70),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_68),
.B(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_71),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_71),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_72),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_74),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_74),
.A2(n_127),
.B(n_208),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_75),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_101),
.B(n_342),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_83),
.B(n_87),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_96),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.C(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_93),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_93),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_96),
.B(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_325),
.A3(n_335),
.B1(n_340),
.B2(n_341),
.C(n_345),
.Y(n_101)
);

AOI321xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_275),
.A3(n_313),
.B1(n_319),
.B2(n_324),
.C(n_346),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_232),
.C(n_271),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_202),
.B(n_231),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_183),
.B(n_201),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_162),
.B(n_182),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_138),
.B(n_161),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_112),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_129),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_124),
.C(n_129),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_132),
.B(n_134),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_132),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_132),
.A2(n_226),
.B1(n_227),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_132),
.A2(n_152),
.B1(n_247),
.B2(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_132),
.A2(n_152),
.B(n_256),
.Y(n_288)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_154),
.B(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_147),
.B(n_160),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_145),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_155),
.B(n_159),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_152),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_164),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_175),
.B2(n_181),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_174),
.C(n_181),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_171),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_185),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_198),
.C(n_199),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_196),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_193),
.C(n_194),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_218),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_219),
.C(n_230),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_224),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_228),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_233),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_251),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_234),
.B(n_251),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_245),
.C(n_250),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_244),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_250),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_248),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_269),
.B2(n_270),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_259),
.C(n_270),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_257),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_265),
.C(n_268),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_262),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_273),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_293),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_276),
.B(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.C(n_292),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_277),
.A2(n_278),
.B1(n_286),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_286),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_288),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_287),
.A2(n_305),
.B(n_309),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_289),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_290),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_311),
.B2(n_312),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_304),
.C(n_312),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_301),
.B(n_302),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_301),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_302),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_302),
.A2(n_327),
.B1(n_331),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_307),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_333),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_327),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);


endmodule