module real_jpeg_12309_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_28),
.B1(n_31),
.B2(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_3),
.A2(n_49),
.B1(n_54),
.B2(n_69),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_37),
.B1(n_39),
.B2(n_69),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_62),
.B(n_65),
.C(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_5),
.B(n_104),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_37),
.B1(n_39),
.B2(n_130),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_5),
.A2(n_87),
.B1(n_90),
.B2(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_84),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_28),
.B1(n_31),
.B2(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_132),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_6),
.A2(n_49),
.B1(n_54),
.B2(n_132),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_136),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_37),
.B1(n_39),
.B2(n_136),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_10),
.A2(n_49),
.B1(n_54),
.B2(n_136),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_30),
.B1(n_65),
.B2(n_66),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_30),
.B1(n_49),
.B2(n_54),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_12),
.A2(n_28),
.B1(n_31),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_12),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_12),
.A2(n_37),
.B1(n_39),
.B2(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_12),
.A2(n_44),
.B1(n_49),
.B2(n_54),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_13),
.A2(n_49),
.B1(n_54),
.B2(n_59),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_59),
.B1(n_65),
.B2(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_59),
.Y(n_115)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_15),
.A2(n_28),
.B1(n_31),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_15),
.A2(n_37),
.B1(n_39),
.B2(n_138),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_15),
.A2(n_49),
.B1(n_54),
.B2(n_138),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_138),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_105),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_85),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_21),
.B(n_75),
.CI(n_85),
.CON(n_307),
.SN(n_307)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_60),
.B2(n_74),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_46),
.C(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_27),
.A2(n_33),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_28),
.A2(n_31),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g191 ( 
.A(n_28),
.B(n_130),
.CON(n_191),
.SN(n_191)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_31),
.A2(n_63),
.B(n_130),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_31),
.B(n_36),
.C(n_37),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_32),
.A2(n_34),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_32),
.A2(n_114),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_33),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_33),
.A2(n_84),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_33),
.A2(n_84),
.B1(n_158),
.B2(n_191),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_33),
.A2(n_42),
.B(n_115),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_34),
.A2(n_83),
.B(n_116),
.Y(n_285)
);

OA22x2_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_35),
.A2(n_39),
.B(n_190),
.C(n_192),
.Y(n_189)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_39),
.B1(n_52),
.B2(n_55),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_39),
.B(n_212),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_45),
.A2(n_46),
.B1(n_113),
.B2(n_118),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_56),
.B(n_58),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_58),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_47),
.A2(n_56),
.B1(n_197),
.B2(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_47),
.A2(n_56),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_47),
.A2(n_56),
.B1(n_205),
.B2(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_47),
.A2(n_56),
.B1(n_96),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_80),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_48),
.A2(n_78),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_48),
.B(n_130),
.Y(n_231)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_SL g55 ( 
.A(n_52),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_52),
.B(n_54),
.C(n_130),
.Y(n_212)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_54),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_56),
.A2(n_58),
.B(n_97),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_56),
.Y(n_195)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_74),
.B1(n_108),
.B2(n_119),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_70),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_61),
.A2(n_100),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_64),
.Y(n_110)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_104),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_104),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_71),
.A2(n_104),
.B1(n_168),
.B2(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_75),
.A2(n_76),
.B(n_81),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_77),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_115),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_93),
.B(n_98),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_86),
.A2(n_94),
.B1(n_95),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_86),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_86),
.A2(n_98),
.B1(n_99),
.B2(n_279),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_91),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_87),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_87),
.A2(n_90),
.B1(n_220),
.B2(n_228),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_87),
.A2(n_222),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_88),
.A2(n_89),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_88),
.B(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_88),
.A2(n_92),
.B(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_88),
.A2(n_89),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_89),
.B(n_92),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_90),
.A2(n_143),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_90),
.B(n_130),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_93),
.B(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_103),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_100),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_102),
.B(n_104),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_304),
.B(n_308),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_293),
.B(n_303),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_274),
.B(n_292),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_181),
.B(n_256),
.C(n_273),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_160),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_126),
.B(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_140),
.C(n_149),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_127),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_134),
.C(n_139),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_140),
.B(n_149),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_147),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.C(n_156),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_150),
.A2(n_154),
.B1(n_155),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_151),
.B(n_238),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_172),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_161),
.B(n_173),
.C(n_180),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_171),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_165),
.B(n_169),
.C(n_171),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_174),
.B(n_178),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_251),
.B(n_255),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_206),
.B(n_250),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_201),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_201),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_198),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_194),
.C(n_198),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_189),
.B(n_193),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.C(n_204),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_204),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_245),
.B(n_249),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_234),
.B(n_244),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_223),
.B(n_233),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_216),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_229),
.B(n_232),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_240),
.C(n_243),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_254),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_272),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_272),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_260),
.C(n_266),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_265),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_263),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_269),
.C(n_270),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_291),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_280),
.B1(n_289),
.B2(n_290),
.Y(n_277)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_290),
.C(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_285),
.C(n_286),
.Y(n_296)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_302),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_302),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);


endmodule