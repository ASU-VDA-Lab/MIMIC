module fake_jpeg_3618_n_619 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_619);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_619;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_14),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_58),
.B(n_64),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_70),
.Y(n_122)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_9),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_76),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_9),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_72),
.B(n_96),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_77),
.B(n_80),
.Y(n_162)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_87),
.Y(n_136)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g177 ( 
.A(n_93),
.Y(n_177)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_10),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_29),
.B(n_36),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_113),
.Y(n_134)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_10),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_102),
.B(n_106),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_22),
.B(n_10),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

BUFx16f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_10),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_115),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_51),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_29),
.B1(n_36),
.B2(n_74),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_117),
.A2(n_123),
.B1(n_137),
.B2(n_165),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_38),
.B1(n_40),
.B2(n_55),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_118),
.A2(n_143),
.B1(n_170),
.B2(n_188),
.Y(n_195)
);

HAxp5_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_29),
.CON(n_120),
.SN(n_120)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_120),
.A2(n_0),
.B(n_42),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_40),
.B1(n_55),
.B2(n_34),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_131),
.A2(n_186),
.B1(n_35),
.B2(n_86),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_55),
.B1(n_40),
.B2(n_57),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_138),
.A2(n_99),
.B1(n_114),
.B2(n_116),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_141),
.B(n_154),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_68),
.A2(n_55),
.B1(n_57),
.B2(n_33),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_142),
.A2(n_24),
.B1(n_49),
.B2(n_27),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_38),
.B1(n_56),
.B2(n_27),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_61),
.B(n_38),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_63),
.B(n_41),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_100),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_62),
.A2(n_20),
.B1(n_42),
.B2(n_41),
.Y(n_170)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_67),
.A2(n_20),
.B1(n_42),
.B2(n_41),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_34),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_65),
.B(n_56),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_84),
.B(n_53),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_65),
.B(n_53),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_78),
.B(n_43),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_97),
.B(n_43),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_92),
.B(n_26),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_69),
.A2(n_33),
.B1(n_49),
.B2(n_24),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_105),
.A2(n_34),
.B1(n_20),
.B2(n_19),
.Y(n_188)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_193),
.Y(n_290)
);

OR2x4_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_93),
.Y(n_194)
);

MAJx3_ASAP7_75t_L g271 ( 
.A(n_194),
.B(n_148),
.C(n_158),
.Y(n_271)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_79),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_198),
.B(n_208),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_199),
.B(n_204),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_147),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_200),
.Y(n_263)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_201),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_202),
.A2(n_248),
.B1(n_249),
.B2(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_85),
.B1(n_94),
.B2(n_101),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_203),
.A2(n_230),
.B1(n_246),
.B2(n_155),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_147),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g206 ( 
.A(n_161),
.B(n_66),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_206),
.A2(n_207),
.B(n_220),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_120),
.B(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_110),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_103),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_211),
.B(n_215),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_180),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_212),
.B(n_227),
.Y(n_318)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_135),
.B(n_103),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_216),
.Y(n_299)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_218),
.Y(n_302)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_219),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_134),
.B(n_98),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_122),
.B(n_109),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_223),
.B(n_224),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_124),
.B(n_98),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_134),
.B(n_113),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_225),
.B(n_2),
.Y(n_315)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_156),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_157),
.B(n_26),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_228),
.B(n_238),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_236),
.Y(n_285)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_237),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_153),
.B(n_175),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_136),
.B(n_35),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_242),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_121),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_241),
.A2(n_251),
.B1(n_173),
.B2(n_166),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_153),
.B(n_35),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_128),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_175),
.B(n_186),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_252),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_148),
.B(n_177),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_174),
.A2(n_104),
.B1(n_91),
.B2(n_90),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_247),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_131),
.A2(n_75),
.B1(n_73),
.B2(n_113),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_134),
.B(n_83),
.C(n_51),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_220),
.C(n_225),
.Y(n_264)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_121),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_140),
.B(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_129),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_138),
.A2(n_83),
.B1(n_51),
.B2(n_0),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_174),
.B(n_0),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_139),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_258),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_189),
.A2(n_164),
.B1(n_160),
.B2(n_169),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_261),
.A2(n_281),
.B1(n_294),
.B2(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_264),
.B(n_266),
.C(n_280),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_148),
.C(n_150),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_SL g328 ( 
.A1(n_271),
.A2(n_245),
.B(n_200),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_274),
.B(n_314),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_199),
.A2(n_128),
.B1(n_130),
.B2(n_150),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_279),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_206),
.B(n_164),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_144),
.B1(n_169),
.B2(n_155),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_205),
.B(n_130),
.CI(n_139),
.CON(n_289),
.SN(n_289)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_289),
.B(n_297),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_195),
.A2(n_173),
.B1(n_132),
.B2(n_166),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_296),
.B(n_191),
.Y(n_332)
);

INVxp67_ASAP7_75t_R g297 ( 
.A(n_194),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_238),
.B(n_158),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_308),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_190),
.B(n_171),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_319),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_232),
.A2(n_171),
.B1(n_125),
.B2(n_132),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_218),
.B1(n_234),
.B2(n_212),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_197),
.B(n_125),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_248),
.A2(n_133),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_207),
.B(n_133),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_251),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_249),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_314),
.A2(n_320),
.B1(n_241),
.B2(n_11),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_315),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_220),
.B(n_5),
.C(n_6),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_256),
.A2(n_17),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_253),
.C(n_225),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_340),
.C(n_367),
.Y(n_378)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_275),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_335),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_328),
.B(n_315),
.Y(n_385)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_267),
.A2(n_213),
.B1(n_233),
.B2(n_204),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_331),
.A2(n_356),
.B1(n_359),
.B2(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_332),
.B(n_346),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_222),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_333),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_334),
.A2(n_352),
.B1(n_354),
.B2(n_302),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_260),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_287),
.B(n_226),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_336),
.B(n_343),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_308),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_337),
.B(n_338),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_287),
.B(n_229),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_239),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_339),
.B(n_342),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_264),
.B(n_209),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_239),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_296),
.B(n_192),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_289),
.B(n_305),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_231),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_217),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_347),
.B(n_364),
.Y(n_397)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_263),
.Y(n_348)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_282),
.B(n_196),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_350),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_219),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_237),
.Y(n_351)
);

A2O1A1O1Ixp25_ASAP7_75t_L g415 ( 
.A1(n_351),
.A2(n_272),
.B(n_278),
.C(n_270),
.D(n_269),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_312),
.A2(n_221),
.B1(n_201),
.B2(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_267),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g359 ( 
.A1(n_271),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_259),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_366),
.Y(n_406)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_265),
.Y(n_362)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_362),
.Y(n_404)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_271),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_285),
.B(n_12),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_365),
.B(n_368),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_259),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_266),
.B(n_280),
.C(n_315),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_283),
.B(n_15),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_272),
.Y(n_369)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_284),
.Y(n_371)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_268),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_374),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_268),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_292),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_376),
.B(n_385),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_325),
.A2(n_292),
.B1(n_289),
.B2(n_297),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_377),
.A2(n_398),
.B(n_409),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_329),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_387),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_345),
.A2(n_317),
.B(n_292),
.C(n_258),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_415),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_341),
.B(n_299),
.C(n_276),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_392),
.C(n_400),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_349),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_391),
.B(n_399),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_261),
.C(n_277),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_395),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_330),
.A2(n_303),
.B(n_290),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_346),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_319),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g402 ( 
.A1(n_330),
.A2(n_284),
.B(n_320),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_402),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_290),
.B(n_286),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_412),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_332),
.A2(n_286),
.B(n_288),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_370),
.B(n_343),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_327),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_417),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_350),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_418),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_373),
.A2(n_273),
.B1(n_302),
.B2(n_262),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_419),
.A2(n_322),
.B1(n_356),
.B2(n_348),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_393),
.B(n_338),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_423),
.B(n_436),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_400),
.C(n_384),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_424),
.B(n_431),
.C(n_447),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_425),
.A2(n_433),
.B1(n_443),
.B2(n_451),
.Y(n_464)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_430),
.A2(n_383),
.B(n_414),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_378),
.B(n_376),
.C(n_323),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_373),
.B1(n_357),
.B2(n_331),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_387),
.A2(n_344),
.B1(n_322),
.B2(n_351),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_434),
.A2(n_421),
.B1(n_389),
.B2(n_390),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_406),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_407),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_438),
.B(n_442),
.Y(n_480)
);

AO22x1_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_359),
.B1(n_370),
.B2(n_369),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_439),
.B(n_450),
.Y(n_472)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_380),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_382),
.A2(n_355),
.B1(n_361),
.B2(n_366),
.Y(n_443)
);

NOR3xp33_ASAP7_75t_SL g444 ( 
.A(n_411),
.B(n_344),
.C(n_355),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_SL g485 ( 
.A(n_444),
.B(n_383),
.C(n_402),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_395),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_445),
.B(n_412),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_323),
.C(n_324),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_385),
.B(n_353),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_452),
.C(n_456),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_398),
.Y(n_449)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_409),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_417),
.A2(n_354),
.B1(n_372),
.B2(n_374),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_363),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_399),
.A2(n_360),
.B1(n_362),
.B2(n_371),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_454),
.A2(n_455),
.B1(n_416),
.B2(n_419),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_410),
.A2(n_288),
.B1(n_262),
.B2(n_278),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_397),
.B(n_269),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_458),
.Y(n_495)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_460),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_381),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_467),
.Y(n_500)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_466),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_422),
.B(n_381),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_468),
.A2(n_478),
.B1(n_481),
.B2(n_485),
.Y(n_515)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_435),
.Y(n_470)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_427),
.A2(n_410),
.B1(n_421),
.B2(n_391),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_451),
.B1(n_439),
.B2(n_433),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_444),
.Y(n_477)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_427),
.A2(n_382),
.B1(n_383),
.B2(n_394),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_437),
.B(n_383),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_479),
.B(n_492),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_428),
.A2(n_450),
.B1(n_446),
.B2(n_459),
.Y(n_481)
);

XNOR2x1_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_452),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_484),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_422),
.B(n_447),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_486),
.B(n_488),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_434),
.B(n_389),
.Y(n_487)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_487),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_402),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_428),
.A2(n_411),
.B1(n_379),
.B2(n_396),
.Y(n_489)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_396),
.C(n_408),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_426),
.C(n_441),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_432),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_454),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_448),
.B(n_401),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_446),
.A2(n_408),
.B1(n_405),
.B2(n_404),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_493),
.A2(n_401),
.B1(n_420),
.B2(n_413),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_413),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_494),
.B(n_430),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_470),
.B(n_461),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_499),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_479),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_502),
.B(n_506),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_503),
.B(n_524),
.Y(n_549)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_474),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_504),
.B(n_510),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_480),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_507),
.B(n_520),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_512),
.B1(n_523),
.B2(n_496),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_468),
.B(n_461),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_509),
.Y(n_550)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_482),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_426),
.C(n_455),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_521),
.C(n_525),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_464),
.A2(n_439),
.B1(n_404),
.B2(n_405),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_415),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_513),
.B(n_514),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_420),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_516),
.A2(n_514),
.B1(n_497),
.B2(n_526),
.Y(n_539)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_495),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_519),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_462),
.B(n_293),
.C(n_316),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_472),
.A2(n_429),
.B(n_457),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_467),
.B(n_465),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_462),
.B(n_316),
.C(n_311),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_508),
.A2(n_481),
.B1(n_478),
.B2(n_483),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_528),
.A2(n_512),
.B1(n_523),
.B2(n_498),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_488),
.C(n_490),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_530),
.B(n_532),
.Y(n_567)
);

OA22x2_ASAP7_75t_L g531 ( 
.A1(n_497),
.A2(n_475),
.B1(n_472),
.B2(n_485),
.Y(n_531)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_476),
.C(n_492),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_540),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_476),
.C(n_473),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_534),
.B(n_538),
.C(n_542),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_536),
.A2(n_551),
.B1(n_516),
.B2(n_515),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_469),
.C(n_463),
.Y(n_538)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_539),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_471),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_469),
.C(n_311),
.Y(n_542)
);

FAx1_ASAP7_75t_SL g543 ( 
.A(n_505),
.B(n_313),
.CI(n_270),
.CON(n_543),
.SN(n_543)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_548),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_544),
.B(n_547),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_517),
.A2(n_307),
.B1(n_518),
.B2(n_498),
.Y(n_545)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_545),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_506),
.B(n_499),
.Y(n_547)
);

FAx1_ASAP7_75t_SL g548 ( 
.A(n_505),
.B(n_307),
.CI(n_501),
.CON(n_548),
.SN(n_548)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_523),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_549),
.B(n_509),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_552),
.B(n_554),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_553),
.A2(n_555),
.B1(n_543),
.B2(n_548),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_549),
.B(n_538),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_522),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_569),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_513),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_560),
.B(n_565),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_504),
.Y(n_562)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_562),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_527),
.B(n_510),
.C(n_519),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_527),
.B(n_530),
.C(n_542),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_568),
.B(n_570),
.C(n_548),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_535),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_534),
.B(n_532),
.C(n_528),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_533),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_531),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_SL g593 ( 
.A(n_572),
.B(n_584),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_563),
.A2(n_551),
.B1(n_550),
.B2(n_537),
.Y(n_573)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_573),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_550),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_574),
.B(n_576),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_558),
.A2(n_546),
.B(n_531),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_566),
.A2(n_546),
.B1(n_531),
.B2(n_535),
.Y(n_577)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_577),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g595 ( 
.A(n_578),
.Y(n_595)
);

NOR2x1_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_543),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_581),
.A2(n_585),
.B(n_570),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_541),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_582),
.B(n_564),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_583),
.B(n_587),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_555),
.A2(n_557),
.B(n_567),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_568),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_557),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_561),
.B(n_571),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_588),
.B(n_561),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_579),
.B(n_585),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_591),
.B(n_592),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_564),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_600),
.Y(n_603)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_596),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_598),
.A2(n_599),
.B(n_595),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_SL g599 ( 
.A(n_583),
.B(n_556),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_586),
.B(n_575),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_584),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_604),
.B(n_593),
.C(n_590),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_589),
.B(n_580),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_605),
.B(n_609),
.Y(n_612)
);

NAND4xp25_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_576),
.C(n_574),
.D(n_577),
.Y(n_607)
);

AO221x1_ASAP7_75t_L g611 ( 
.A1(n_607),
.A2(n_608),
.B1(n_573),
.B2(n_597),
.C(n_593),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_595),
.B(n_580),
.Y(n_608)
);

AOI31xp33_ASAP7_75t_L g615 ( 
.A1(n_610),
.A2(n_611),
.A3(n_613),
.B(n_605),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_588),
.C(n_572),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_612),
.B(n_606),
.C(n_603),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_614),
.A2(n_615),
.B(n_612),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_581),
.Y(n_617)
);

BUFx24_ASAP7_75t_SL g618 ( 
.A(n_617),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_618),
.B(n_578),
.Y(n_619)
);


endmodule