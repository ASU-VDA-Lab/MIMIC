module fake_jpeg_2030_n_548 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_548);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_548;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_60),
.Y(n_204)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_84),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_65),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_76),
.Y(n_153)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_71),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_72),
.Y(n_165)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_49),
.Y(n_80)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_82),
.B(n_85),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_32),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_15),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_91),
.Y(n_189)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_46),
.B(n_15),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_15),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_94),
.B(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_95),
.B(n_98),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_99),
.B(n_102),
.Y(n_197)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_45),
.B(n_14),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_12),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_106),
.B(n_107),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_22),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_42),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_109),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_12),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_114),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_30),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_118),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_31),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_119),
.B(n_120),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_19),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_123),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_126),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_33),
.B1(n_50),
.B2(n_37),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_42),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_33),
.B1(n_50),
.B2(n_37),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_142),
.A2(n_155),
.B1(n_183),
.B2(n_213),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_27),
.B1(n_36),
.B2(n_31),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_146),
.A2(n_147),
.B1(n_158),
.B2(n_214),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_74),
.A2(n_93),
.B1(n_83),
.B2(n_92),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_64),
.A2(n_67),
.B1(n_126),
.B2(n_80),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_150),
.A2(n_151),
.B1(n_162),
.B2(n_185),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_64),
.A2(n_54),
.B1(n_52),
.B2(n_51),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_154),
.B(n_159),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_69),
.A2(n_36),
.B1(n_54),
.B2(n_25),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_72),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_156),
.B(n_170),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_96),
.A2(n_23),
.B1(n_51),
.B2(n_47),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_87),
.B(n_23),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_52),
.B1(n_47),
.B2(n_44),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_70),
.B(n_43),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_163),
.B(n_167),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_111),
.A2(n_43),
.B(n_39),
.C(n_25),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_152),
.B(n_130),
.C(n_197),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_44),
.B1(n_39),
.B2(n_3),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g271 ( 
.A1(n_166),
.A2(n_169),
.B1(n_178),
.B2(n_196),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_88),
.B(n_0),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_0),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_168),
.B(n_176),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_58),
.B(n_1),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_59),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_71),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_90),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_103),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_186),
.B(n_192),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_122),
.A2(n_11),
.B1(n_90),
.B2(n_101),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_187),
.A2(n_195),
.B1(n_211),
.B2(n_150),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_11),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_118),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_193),
.B(n_200),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_122),
.A2(n_101),
.B1(n_60),
.B2(n_119),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_120),
.B(n_99),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_199),
.B(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_84),
.B(n_94),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_102),
.B(n_85),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_64),
.A2(n_67),
.B1(n_49),
.B2(n_126),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_61),
.B(n_62),
.C(n_75),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_148),
.C(n_140),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_110),
.A2(n_104),
.B1(n_94),
.B2(n_84),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_104),
.A2(n_62),
.B1(n_61),
.B2(n_94),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_169),
.B1(n_178),
.B2(n_205),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_219),
.B(n_224),
.C(n_230),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_189),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_220),
.B(n_234),
.Y(n_293)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_131),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_222),
.B(n_223),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_131),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_228),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_132),
.B(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_231),
.B(n_278),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_148),
.B(n_135),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g334 ( 
.A1(n_232),
.A2(n_233),
.B(n_235),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_153),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_149),
.C(n_161),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_160),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_243),
.B(n_244),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_131),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_191),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_245),
.B(n_246),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_137),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_182),
.C(n_137),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_249),
.B(n_256),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_164),
.A2(n_211),
.B(n_162),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_273),
.B(n_253),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g330 ( 
.A1(n_253),
.A2(n_279),
.B(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_171),
.B(n_191),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_134),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_134),
.Y(n_259)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_136),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_210),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_263),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_204),
.Y(n_265)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_266),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_203),
.A2(n_184),
.B1(n_202),
.B2(n_128),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_267),
.A2(n_271),
.B1(n_275),
.B2(n_282),
.Y(n_318)
);

CKINVDCx9p33_ASAP7_75t_R g268 ( 
.A(n_147),
.Y(n_268)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_127),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_270),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_202),
.B(n_196),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_274),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_133),
.A2(n_151),
.B(n_195),
.C(n_128),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_203),
.A2(n_136),
.B1(n_143),
.B2(n_145),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_281),
.Y(n_307)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_138),
.B(n_139),
.Y(n_278)
);

HB1xp67_ASAP7_75t_SL g279 ( 
.A(n_185),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_139),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_190),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_143),
.A2(n_145),
.B1(n_190),
.B2(n_179),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_175),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_278),
.B(n_285),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_141),
.Y(n_284)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_270),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_187),
.A2(n_177),
.B1(n_209),
.B2(n_141),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_286),
.A2(n_232),
.B1(n_283),
.B2(n_253),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_177),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_225),
.B1(n_271),
.B2(n_252),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_295),
.A2(n_318),
.B(n_303),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_251),
.A2(n_271),
.B1(n_231),
.B2(n_225),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_303),
.B1(n_325),
.B2(n_236),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_236),
.B1(n_253),
.B2(n_242),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_306),
.A2(n_309),
.B(n_236),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_246),
.A2(n_243),
.B(n_219),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g316 ( 
.A(n_250),
.B(n_262),
.C(n_227),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_228),
.C(n_288),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g317 ( 
.A(n_233),
.B(n_255),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_232),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_237),
.A2(n_229),
.B1(n_247),
.B2(n_216),
.Y(n_325)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_257),
.B(n_235),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_257),
.B(n_250),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_216),
.A2(n_221),
.B1(n_274),
.B2(n_276),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_283),
.B1(n_281),
.B2(n_269),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_236),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_348),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_327),
.B(n_224),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_338),
.B(n_347),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_360),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_230),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_341),
.C(n_343),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_215),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_254),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_344),
.A2(n_361),
.B(n_372),
.Y(n_390)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_332),
.B(n_249),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_346),
.B(n_367),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_327),
.B(n_239),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_355),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_331),
.B(n_248),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_289),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_354),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_218),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_241),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_357),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_306),
.A2(n_280),
.B1(n_259),
.B2(n_258),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_313),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_359),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_265),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_307),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_309),
.A2(n_244),
.B(n_260),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_362),
.A2(n_296),
.B(n_320),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_226),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_364),
.Y(n_395)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_368),
.B(n_369),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_310),
.B(n_238),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_312),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_370),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_336),
.A2(n_266),
.B1(n_277),
.B2(n_294),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_378),
.B1(n_337),
.B2(n_361),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_297),
.B(n_291),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_302),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_324),
.C(n_326),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_298),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_374),
.A2(n_376),
.B(n_377),
.Y(n_402)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_375),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_291),
.B(n_326),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_294),
.A2(n_295),
.B1(n_330),
.B2(n_290),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_365),
.B(n_317),
.CI(n_316),
.CON(n_382),
.SN(n_382)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_382),
.B(n_409),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_SL g437 ( 
.A1(n_383),
.A2(n_363),
.B(n_372),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_348),
.A2(n_295),
.B1(n_290),
.B2(n_307),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_384),
.A2(n_410),
.B1(n_357),
.B2(n_376),
.Y(n_425)
);

XOR2x2_ASAP7_75t_SL g388 ( 
.A(n_365),
.B(n_304),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_397),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_356),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_289),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_399),
.C(n_404),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_328),
.C(n_300),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_344),
.A2(n_298),
.B(n_296),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_400),
.A2(n_411),
.B(n_402),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_305),
.B1(n_335),
.B2(n_322),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_401),
.A2(n_376),
.B1(n_354),
.B2(n_352),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_328),
.C(n_301),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_301),
.C(n_299),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_362),
.C(n_375),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_359),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_337),
.A2(n_322),
.B1(n_335),
.B2(n_321),
.Y(n_410)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_411),
.A2(n_377),
.B(n_369),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_360),
.Y(n_413)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_342),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_415),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_385),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_390),
.A2(n_361),
.B(n_337),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_416),
.A2(n_431),
.B(n_433),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_405),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_417),
.B(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_342),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_361),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_430),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_438),
.C(n_439),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_424),
.A2(n_425),
.B1(n_442),
.B2(n_391),
.Y(n_451)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_405),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_428),
.B(n_436),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_407),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_370),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_435),
.Y(n_452)
);

NAND2x1_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_378),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_371),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_434),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_379),
.B(n_340),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_351),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_384),
.B1(n_408),
.B2(n_386),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_346),
.C(n_339),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_358),
.C(n_343),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_440),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_381),
.B(n_341),
.Y(n_441)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_403),
.B(n_380),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_425),
.A2(n_386),
.B1(n_380),
.B2(n_387),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_444),
.A2(n_451),
.B1(n_453),
.B2(n_454),
.Y(n_484)
);

AOI322xp5_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_403),
.A3(n_382),
.B1(n_386),
.B2(n_408),
.C1(n_402),
.C2(n_390),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_447),
.B(n_415),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_450),
.A2(n_465),
.B(n_431),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_422),
.A2(n_428),
.B1(n_430),
.B2(n_387),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_422),
.A2(n_391),
.B1(n_395),
.B2(n_389),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_392),
.C(n_404),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_458),
.C(n_464),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_414),
.A2(n_401),
.B1(n_395),
.B2(n_389),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_457),
.A2(n_436),
.B1(n_442),
.B2(n_434),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_394),
.C(n_388),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_427),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_406),
.C(n_347),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_434),
.A2(n_398),
.B1(n_406),
.B2(n_374),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_364),
.C(n_367),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_423),
.C(n_458),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_462),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_480),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_420),
.Y(n_470)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_452),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_471),
.A2(n_485),
.B1(n_487),
.B2(n_488),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_472),
.A2(n_475),
.B(n_476),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_439),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_478),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_463),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_481),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_431),
.B(n_416),
.C(n_418),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_466),
.A2(n_433),
.B(n_418),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_460),
.C(n_467),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_482),
.C(n_483),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_462),
.Y(n_480)
);

OA21x2_ASAP7_75t_SL g481 ( 
.A1(n_446),
.A2(n_413),
.B(n_382),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_427),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g485 ( 
.A(n_457),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_443),
.Y(n_486)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_486),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_433),
.C(n_440),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_443),
.C(n_461),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_485),
.A2(n_444),
.B1(n_461),
.B2(n_453),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_494),
.A2(n_498),
.B1(n_504),
.B2(n_484),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_SL g496 ( 
.A(n_478),
.B(n_450),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_469),
.A2(n_461),
.B1(n_448),
.B2(n_454),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_501),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_503),
.Y(n_510)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_486),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_476),
.A2(n_461),
.B(n_468),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_468),
.B1(n_459),
.B2(n_463),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_491),
.A2(n_484),
.B1(n_487),
.B2(n_475),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_506),
.A2(n_495),
.B1(n_494),
.B2(n_474),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_504),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_481),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_509),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_505),
.B(n_479),
.C(n_473),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_488),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_512),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_492),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_489),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_493),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_493),
.B(n_477),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_517),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_502),
.B(n_482),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_483),
.C(n_477),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_502),
.A2(n_472),
.B(n_465),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_519),
.A2(n_526),
.B(n_509),
.Y(n_531)
);

AO21x1_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_492),
.B(n_498),
.Y(n_520)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_520),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_510),
.A2(n_503),
.B(n_490),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_523),
.A2(n_518),
.B(n_515),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g530 ( 
.A(n_524),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_528),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_516),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_520),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_533),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_531),
.A2(n_534),
.B(n_522),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_513),
.C(n_510),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_527),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_535),
.B(n_398),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_539),
.B(n_540),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_533),
.A2(n_518),
.B(n_523),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_534),
.A2(n_524),
.B(n_449),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_445),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_530),
.C(n_532),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_542),
.Y(n_546)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_543),
.Y(n_545)
);

AOI321xp33_ASAP7_75t_SL g547 ( 
.A1(n_546),
.A2(n_544),
.A3(n_536),
.B1(n_545),
.B2(n_426),
.C(n_421),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_374),
.Y(n_548)
);


endmodule