module fake_jpeg_9521_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_52),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_46),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_19),
.B1(n_32),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_65),
.B1(n_34),
.B2(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_35),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_19),
.B1(n_32),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_18),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_19),
.B1(n_17),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_66),
.B1(n_23),
.B2(n_28),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_57),
.Y(n_80)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_69),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_17),
.B1(n_31),
.B2(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_1),
.Y(n_86)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_72),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_83),
.B1(n_92),
.B2(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_74),
.B(n_82),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_58),
.B1(n_69),
.B2(n_54),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_88),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_41),
.B(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_103),
.B1(n_51),
.B2(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_84),
.B(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_16),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_37),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_97),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_37),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_44),
.CI(n_43),
.CON(n_129),
.SN(n_129)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_58),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_51),
.A2(n_44),
.B1(n_43),
.B2(n_36),
.Y(n_103)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_111),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_117),
.B1(n_81),
.B2(n_93),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_114),
.B1(n_131),
.B2(n_70),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_41),
.B(n_49),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_44),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_100),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_41),
.B(n_44),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_49),
.B(n_41),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_101),
.B(n_97),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_146),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_90),
.B(n_84),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_149),
.B(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_77),
.B1(n_90),
.B2(n_86),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_143),
.B1(n_110),
.B2(n_114),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_76),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_144),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_77),
.B1(n_87),
.B2(n_98),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_87),
.B(n_71),
.C(n_86),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_94),
.C(n_103),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_112),
.C(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_155),
.B1(n_163),
.B2(n_116),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_132),
.C(n_108),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_124),
.C(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_92),
.B1(n_50),
.B2(n_44),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_92),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_159),
.B(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_125),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_41),
.B(n_49),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_43),
.A3(n_36),
.B1(n_41),
.B2(n_7),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_43),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_129),
.A2(n_50),
.B1(n_78),
.B2(n_6),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_165),
.B(n_168),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_157),
.A2(n_117),
.B1(n_131),
.B2(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_171),
.Y(n_197)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_180),
.C(n_183),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_177),
.B(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_188),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_115),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_150),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_116),
.C(n_111),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_118),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_186),
.C(n_189),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_50),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_107),
.C(n_5),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_1),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_5),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_186),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_160),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_204),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.C(n_174),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_159),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_156),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_144),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_211),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_173),
.A2(n_142),
.B(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_136),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_141),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_177),
.B1(n_164),
.B2(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_225),
.C(n_230),
.Y(n_241)
);

XOR2x1_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_212),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_228),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_173),
.B1(n_172),
.B2(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_180),
.C(n_184),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_197),
.B1(n_198),
.B2(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_215),
.B1(n_210),
.B2(n_209),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_170),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_154),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_221),
.C(n_225),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_202),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_242),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_218),
.B1(n_214),
.B2(n_230),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_229),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_205),
.B(n_156),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_222),
.B1(n_220),
.B2(n_202),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_249),
.C(n_162),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_191),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_216),
.C(n_199),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_227),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_265),
.C(n_241),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_239),
.B(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_232),
.B1(n_228),
.B2(n_235),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_239),
.B1(n_252),
.B2(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_263),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_247),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_264),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_138),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_6),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_246),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_10),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_140),
.B1(n_241),
.B2(n_107),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_7),
.C(n_9),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_10),
.C(n_11),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_10),
.B(n_12),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_258),
.B(n_260),
.C(n_13),
.D(n_15),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_280),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_268),
.B(n_277),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_276),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_271),
.B(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_281),
.B(n_278),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_289),
.B(n_283),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_269),
.C(n_272),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_288),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_294),
.B(n_291),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_15),
.Y(n_297)
);


endmodule