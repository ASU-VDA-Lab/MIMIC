module fake_jpeg_19448_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx2_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx3_ASAP7_75t_SL g71 ( 
.A(n_3),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_0),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_2),
.B(n_3),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_56),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_93),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_63),
.B1(n_48),
.B2(n_56),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_97),
.B1(n_15),
.B2(n_16),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_63),
.B1(n_48),
.B2(n_57),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_106),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_52),
.B(n_59),
.C(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_5),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_74),
.B1(n_67),
.B2(n_68),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_62),
.B1(n_70),
.B2(n_64),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_61),
.B1(n_60),
.B2(n_54),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_75),
.B1(n_53),
.B2(n_5),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_28),
.B1(n_11),
.B2(n_12),
.Y(n_115)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_120),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_124),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_25),
.B(n_26),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_45),
.B(n_34),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_30),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_32),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_132),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_108),
.B1(n_124),
.B2(n_40),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_131),
.C(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_146),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_142),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_129),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_145),
.B1(n_137),
.B2(n_130),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_139),
.C(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_156),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_140),
.C(n_39),
.Y(n_158)
);


endmodule