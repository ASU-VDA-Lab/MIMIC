module fake_netlist_1_2924_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_1), .B(n_0), .Y(n_4) );
AND2x2_ASAP7_75t_L g5 ( .A(n_2), .B(n_0), .Y(n_5) );
INVx4_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
OR2x2_ASAP7_75t_L g7 ( .A(n_3), .B(n_2), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_6), .B(n_5), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_0), .Y(n_10) );
OAI221xp5_ASAP7_75t_SL g11 ( .A1(n_10), .A2(n_9), .B1(n_3), .B2(n_2), .C(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_11), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_12), .B(n_1), .Y(n_13) );
NAND2x1p5_ASAP7_75t_SL g14 ( .A(n_13), .B(n_2), .Y(n_14) );
endmodule