module fake_ibex_837_n_4719 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4719);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4719;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_4688;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4687;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_4632;
wire n_1080;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_4514;
wire n_3838;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_4668;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3653;
wire n_3458;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_3904;
wire n_4378;
wire n_4239;
wire n_3175;
wire n_3729;
wire n_4169;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_4418;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4708;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_4652;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_4673;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_4690;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_3242;
wire n_3395;
wire n_4403;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_4672;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3668;
wire n_3699;
wire n_1955;
wire n_3197;
wire n_4312;
wire n_4567;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_4014;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_3030;
wire n_3097;
wire n_2906;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_4667;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_4711;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_4671;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_4499;
wire n_2957;
wire n_4676;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_4714;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_4258;
wire n_3874;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_4252;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_3909;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_4692;
wire n_4713;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_4615;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3963;
wire n_3887;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_4710;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_4680;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_4693;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4549;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_4098;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_4700;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4523;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_4712;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3634;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3788;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_4571;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4681;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_4374;
wire n_4501;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_3815;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3529;
wire n_1711;
wire n_3222;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_4033;
wire n_4485;
wire n_3855;
wire n_4608;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_1990;
wire n_1179;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_2935;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1566;
wire n_1464;
wire n_4362;
wire n_3568;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_4706;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4674;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4679;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_1115;
wire n_1729;
wire n_1395;
wire n_998;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4660;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_4664;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_4709;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3948;
wire n_3719;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_4077;
wire n_3897;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4255;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_4683;
wire n_3557;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_4694;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_4717;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1683;
wire n_1185;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_2728;
wire n_3772;
wire n_4685;
wire n_2948;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_3657;
wire n_4716;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1997;
wire n_1162;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_2997;
wire n_3314;
wire n_991;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_1349;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_4704;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4142;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1694;
wire n_1458;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_4066;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4123;
wire n_3154;
wire n_4000;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_4007;
wire n_3960;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_4707;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_4695;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1860;
wire n_1491;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_4638;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_4319;
wire n_3760;
wire n_4637;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4212;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_3162;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_4697;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1642;
wire n_1871;
wire n_1455;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_4715;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_4410;
wire n_3574;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_4698;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4162;
wire n_4111;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_4666;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_4663;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_1622;
wire n_2757;
wire n_4611;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_4670;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1542;
wire n_1586;
wire n_1547;
wire n_1362;
wire n_3497;
wire n_4696;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_3586;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2593;
wire n_3899;
wire n_1623;
wire n_2911;
wire n_4279;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_4345;
wire n_4281;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_4675;
wire n_3083;
wire n_2083;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_3844;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_4045;
wire n_4432;
wire n_2405;
wire n_3380;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3742;
wire n_3655;
wire n_4552;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_3791;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_1285;
wire n_3042;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_4686;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4682;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_4705;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_4301;
wire n_3176;
wire n_4471;
wire n_4107;
wire n_3297;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_4684;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_1193;
wire n_2928;
wire n_3225;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3483;
wire n_1074;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3823;
wire n_3369;
wire n_4718;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1904;
wire n_1262;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_1022;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_999;
wire n_2634;
wire n_2982;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1027;
wire n_1516;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2303;
wire n_2618;
wire n_2357;
wire n_2855;
wire n_4354;
wire n_3938;
wire n_4448;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_4701;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_4544;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2961;
wire n_2770;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_4689;
wire n_3613;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_4702;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_4506;
wire n_2073;
wire n_4093;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_1551;
wire n_4153;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3988;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3406;
wire n_4327;
wire n_2656;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_4703;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_4691;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_450),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_708),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_592),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_445),
.Y(n_977)
);

INVxp33_ASAP7_75t_L g978 ( 
.A(n_91),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_971),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_190),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_683),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_653),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_473),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_815),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_634),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_642),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_591),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_184),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_621),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_473),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_820),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_69),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_640),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_130),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_897),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_947),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_182),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_549),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_27),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_911),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_282),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_768),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_814),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_955),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_960),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_566),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_753),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_260),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_746),
.Y(n_1009)
);

CKINVDCx14_ASAP7_75t_R g1010 ( 
.A(n_306),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_954),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_654),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_854),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_873),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_831),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_312),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_829),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_482),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_929),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_965),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_760),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_508),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_821),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_467),
.Y(n_1024)
);

BUFx10_ASAP7_75t_L g1025 ( 
.A(n_427),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_928),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_529),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_514),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_832),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_165),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_687),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_819),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_319),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_731),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_210),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_662),
.Y(n_1036)
);

BUFx5_ASAP7_75t_L g1037 ( 
.A(n_175),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_520),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_218),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_141),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_943),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_160),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_903),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_743),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_935),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_731),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_576),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_286),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_313),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_248),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_937),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_935),
.Y(n_1052)
);

CKINVDCx16_ASAP7_75t_R g1053 ( 
.A(n_693),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_43),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_683),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_550),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_177),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_644),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_628),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_562),
.Y(n_1060)
);

BUFx8_ASAP7_75t_SL g1061 ( 
.A(n_344),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_298),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_373),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_567),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_515),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_18),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_636),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_667),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_239),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_144),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_284),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_76),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_878),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_121),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_26),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_451),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_930),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_14),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_279),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_428),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_340),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_255),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_856),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_913),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_500),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_476),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_18),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_908),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_368),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_296),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_196),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_931),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_258),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_406),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_89),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_912),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_181),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_809),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_813),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_946),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_280),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_701),
.Y(n_1102)
);

BUFx10_ASAP7_75t_L g1103 ( 
.A(n_566),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_797),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_884),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_765),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_396),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_815),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_831),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_34),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_926),
.Y(n_1111)
);

CKINVDCx14_ASAP7_75t_R g1112 ( 
.A(n_916),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_647),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_488),
.Y(n_1114)
);

CKINVDCx16_ASAP7_75t_R g1115 ( 
.A(n_517),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_519),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_14),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_940),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_547),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_812),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_80),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_247),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_345),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_910),
.Y(n_1124)
);

CKINVDCx16_ASAP7_75t_R g1125 ( 
.A(n_688),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_208),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_909),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_453),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_715),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_81),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_294),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_150),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_118),
.Y(n_1133)
);

CKINVDCx14_ASAP7_75t_R g1134 ( 
.A(n_358),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_956),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_735),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_854),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_415),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_712),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_472),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_900),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_956),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_372),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_101),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_973),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_155),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_501),
.Y(n_1147)
);

BUFx5_ASAP7_75t_L g1148 ( 
.A(n_519),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_844),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_53),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_158),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_535),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_847),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_955),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_361),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_68),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_722),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_612),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_905),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_870),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_214),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_545),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_549),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_281),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_514),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_655),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_653),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_902),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_886),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_950),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_225),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_806),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_88),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_425),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_74),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_149),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_209),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_154),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_777),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_835),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_946),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_405),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_690),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_98),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_582),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_684),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_351),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_926),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_873),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_482),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_529),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_282),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_588),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_747),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_786),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_601),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_323),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_680),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_658),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_145),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_789),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_63),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_631),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_637),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_148),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_927),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_370),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_884),
.Y(n_1208)
);

BUFx5_ASAP7_75t_L g1209 ( 
.A(n_932),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_907),
.Y(n_1210)
);

CKINVDCx16_ASAP7_75t_R g1211 ( 
.A(n_941),
.Y(n_1211)
);

CKINVDCx16_ASAP7_75t_R g1212 ( 
.A(n_501),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_207),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_899),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_811),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_596),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_959),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_853),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_599),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_585),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_70),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_662),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_82),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_37),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_225),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_185),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_575),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_941),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_53),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_664),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_634),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_936),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_686),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_713),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_508),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_670),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_432),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_592),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_852),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_661),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_641),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_356),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_548),
.Y(n_1243)
);

BUFx10_ASAP7_75t_L g1244 ( 
.A(n_617),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_198),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_313),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_769),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_587),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_132),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_573),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_715),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_412),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_75),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_708),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_906),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_340),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_329),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_57),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_217),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_137),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_921),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_670),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_966),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_787),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_701),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_668),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_958),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_856),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_456),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_184),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_898),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_744),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_627),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_680),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_86),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_271),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_320),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_575),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_917),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_522),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_819),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_539),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_925),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_937),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_172),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_844),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_874),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_698),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_484),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_350),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_830),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_81),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_404),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_618),
.Y(n_1294)
);

BUFx5_ASAP7_75t_L g1295 ( 
.A(n_720),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_312),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_738),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_554),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_207),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_147),
.Y(n_1300)
);

CKINVDCx14_ASAP7_75t_R g1301 ( 
.A(n_358),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_952),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_743),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_939),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_127),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_41),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_589),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_202),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_909),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_412),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_759),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_934),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_671),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_180),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_945),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_389),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_6),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_287),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_370),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_326),
.Y(n_1320)
);

BUFx10_ASAP7_75t_L g1321 ( 
.A(n_586),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_276),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_580),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_260),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_264),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_15),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_933),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_399),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_787),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_918),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_377),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_466),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_923),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_151),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_206),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_804),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_407),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_289),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_250),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_230),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_66),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_948),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_124),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_841),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_866),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_763),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_924),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_838),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_792),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_124),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_735),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_203),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_176),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_717),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_25),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_938),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_919),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_957),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_435),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_539),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_277),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_953),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_632),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_53),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_951),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_132),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_694),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_879),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_668),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_175),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_839),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_392),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_882),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_460),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_87),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_465),
.Y(n_1376)
);

CKINVDCx16_ASAP7_75t_R g1377 ( 
.A(n_534),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_555),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_771),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_807),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_389),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_643),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_724),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_824),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_52),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_703),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_163),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_244),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_922),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_376),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_204),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_409),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_601),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_418),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_174),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_312),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_716),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_887),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_137),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_880),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_949),
.Y(n_1401)
);

CKINVDCx14_ASAP7_75t_R g1402 ( 
.A(n_600),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_223),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_118),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_276),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_497),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_944),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_964),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_85),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_493),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_452),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_915),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_712),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_904),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_890),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_439),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_158),
.Y(n_1417)
);

CKINVDCx16_ASAP7_75t_R g1418 ( 
.A(n_597),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_916),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_229),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_448),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_729),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_902),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_449),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_942),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_177),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_451),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_600),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_713),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_528),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_261),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_72),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_824),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_781),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_652),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_51),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_822),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_480),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_323),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_710),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_877),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_613),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_276),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_825),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_848),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_901),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_36),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_591),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_26),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_657),
.Y(n_1450)
);

BUFx5_ASAP7_75t_L g1451 ( 
.A(n_718),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_781),
.Y(n_1452)
);

BUFx10_ASAP7_75t_L g1453 ( 
.A(n_292),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_545),
.Y(n_1454)
);

BUFx10_ASAP7_75t_L g1455 ( 
.A(n_859),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_544),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_144),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_837),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_129),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_914),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_98),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_920),
.Y(n_1462)
);

BUFx10_ASAP7_75t_L g1463 ( 
.A(n_528),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_445),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_915),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_495),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_597),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_943),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_542),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_431),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_315),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_806),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_441),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_19),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_113),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_421),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_101),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_965),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_372),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_896),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_807),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_784),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_966),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_864),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_602),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_358),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_307),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_274),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_569),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_773),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_359),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_823),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_678),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_338),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_396),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_82),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1010),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1061),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1100),
.B(n_1027),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_1139),
.B(n_0),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1076),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1061),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1134),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1094),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1134),
.B(n_0),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1301),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1112),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1178),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1381),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_994),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1048),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_994),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1331),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1331),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1112),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_978),
.B(n_1),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1402),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1402),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1082),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1477),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1115),
.B(n_1),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1049),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1187),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1212),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1377),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_974),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_977),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1341),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1375),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_983),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1477),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1209),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_980),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_988),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_997),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_978),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1026),
.B(n_1),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1016),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1022),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_1064),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1174),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1038),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_999),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1267),
.B(n_2),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1057),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1008),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1062),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1063),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1018),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1164),
.Y(n_1550)
);

INVxp33_ASAP7_75t_SL g1551 ( 
.A(n_1369),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1478),
.B(n_2),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1024),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1070),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1075),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1165),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1226),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1028),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1256),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1053),
.B(n_3),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1411),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1424),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1030),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1347),
.B(n_2),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1110),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1116),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1317),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1033),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1466),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1130),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1001),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1496),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1035),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1143),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1350),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1171),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1197),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1116),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1221),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1235),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1039),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1125),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1040),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1350),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1211),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1343),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_SL g1587 ( 
.A(n_1001),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1042),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1259),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1243),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1050),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1054),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1575),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1536),
.B(n_1351),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1001),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1510),
.A2(n_1315),
.B1(n_1311),
.B2(n_1019),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1532),
.A2(n_1069),
.B(n_992),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1065),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1511),
.B(n_1398),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1575),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1501),
.B(n_1120),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1526),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1566),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1504),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1584),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1508),
.Y(n_1606)
);

INVx6_ASAP7_75t_L g1607 ( 
.A(n_1516),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1541),
.Y(n_1608)
);

AND2x2_ASAP7_75t_SL g1609 ( 
.A(n_1560),
.B(n_1418),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1522),
.B(n_1400),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1586),
.B(n_1025),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1566),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1509),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1527),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1497),
.B(n_1066),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1587),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1564),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1538),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1539),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1566),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1542),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1545),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1547),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1548),
.A2(n_1069),
.B(n_992),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1512),
.A2(n_1315),
.B1(n_1311),
.B2(n_1105),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1499),
.B(n_1025),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1554),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1555),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1565),
.Y(n_1631)
);

BUFx8_ASAP7_75t_L g1632 ( 
.A(n_1523),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1570),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1574),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1566),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1578),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1578),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1578),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1576),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1577),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1579),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1580),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1505),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1589),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1578),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1537),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1528),
.B(n_982),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1529),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1503),
.B(n_982),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1544),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1500),
.A2(n_1146),
.B(n_1086),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1552),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1530),
.B(n_1037),
.Y(n_1653)
);

AND2x6_ASAP7_75t_L g1654 ( 
.A(n_1521),
.B(n_1372),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1507),
.B(n_1002),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1534),
.B(n_1080),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1535),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_1513),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1543),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1546),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1515),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1549),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1553),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1558),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1563),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1568),
.B(n_1037),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1592),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1572),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1573),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1581),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1517),
.B(n_1002),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1583),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1591),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1588),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1518),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1551),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1519),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1524),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1525),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1506),
.B(n_1037),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1533),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1582),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1585),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1590),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1498),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1502),
.Y(n_1686)
);

INVx5_ASAP7_75t_L g1687 ( 
.A(n_1550),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1556),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1557),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1514),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1520),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1559),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1531),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1561),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1562),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1569),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1532),
.Y(n_1697)
);

XNOR2xp5_ASAP7_75t_L g1698 ( 
.A(n_1510),
.B(n_1012),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1584),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1536),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1575),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1571),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1575),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1575),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1532),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1536),
.B(n_1003),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1536),
.B(n_1071),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1532),
.A2(n_1335),
.B(n_1151),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1575),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1532),
.A2(n_1335),
.B(n_1151),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1571),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1575),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1526),
.Y(n_1713)
);

AND2x2_ASAP7_75t_SL g1714 ( 
.A(n_1516),
.B(n_1004),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1587),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1532),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1575),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1532),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1575),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1575),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1575),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1587),
.B(n_1080),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1536),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1575),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1571),
.B(n_1148),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1571),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1536),
.B(n_1072),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1575),
.Y(n_1728)
);

NAND2x1_ASAP7_75t_L g1729 ( 
.A(n_1571),
.B(n_1353),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1536),
.B(n_1078),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1575),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1566),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1536),
.B(n_1079),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1536),
.B(n_1080),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1536),
.B(n_1081),
.Y(n_1735)
);

BUFx8_ASAP7_75t_L g1736 ( 
.A(n_1587),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1536),
.B(n_1091),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1575),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1575),
.Y(n_1739)
);

BUFx8_ASAP7_75t_L g1740 ( 
.A(n_1587),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1575),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1575),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1575),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1571),
.B(n_1148),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1536),
.B(n_1003),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1575),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1536),
.B(n_1085),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1536),
.B(n_1453),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1575),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1571),
.B(n_1148),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1575),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1587),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1536),
.B(n_1453),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1571),
.B(n_1148),
.Y(n_1754)
);

BUFx8_ASAP7_75t_L g1755 ( 
.A(n_1587),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1566),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_SL g1757 ( 
.A(n_1587),
.B(n_1453),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1575),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1575),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1575),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1575),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1532),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1587),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1618),
.B(n_1148),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1604),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1606),
.Y(n_1766)
);

INVx5_ASAP7_75t_L g1767 ( 
.A(n_1702),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1652),
.B(n_1087),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1736),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1650),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1650),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1626),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1614),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1713),
.B(n_990),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1711),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1631),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1700),
.B(n_1074),
.Y(n_1777)
);

INVx5_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_1699),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1615),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1633),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1595),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1700),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1688),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1597),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1723),
.B(n_1089),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1646),
.B(n_1463),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1646),
.Y(n_1788)
);

BUFx10_ASAP7_75t_L g1789 ( 
.A(n_1617),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_SL g1790 ( 
.A(n_1689),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1736),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1594),
.B(n_1230),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1734),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1740),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1620),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1611),
.B(n_1463),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_R g1797 ( 
.A(n_1715),
.B(n_1129),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1594),
.B(n_1090),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1737),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1740),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1707),
.B(n_1144),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1646),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1597),
.Y(n_1803)
);

INVx1_ASAP7_75t_SL g1804 ( 
.A(n_1748),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1753),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1708),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1727),
.B(n_1093),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1708),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1710),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1656),
.B(n_1463),
.Y(n_1810)
);

OR2x6_ASAP7_75t_SL g1811 ( 
.A(n_1752),
.B(n_1095),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1755),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1730),
.B(n_1733),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1735),
.B(n_1097),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1607),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1607),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1608),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1628),
.B(n_1643),
.Y(n_1818)
);

AND2x6_ASAP7_75t_L g1819 ( 
.A(n_1672),
.B(n_1372),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1602),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1755),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1613),
.A2(n_1600),
.B1(n_1701),
.B2(n_1593),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1660),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1747),
.B(n_1101),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1706),
.B(n_1107),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1643),
.B(n_1152),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1706),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1676),
.B(n_1173),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1710),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1722),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1669),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1658),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1745),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1745),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1619),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1598),
.B(n_1114),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1703),
.B(n_993),
.Y(n_1837)
);

OAI22xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1757),
.A2(n_1121),
.B1(n_1122),
.B2(n_1117),
.Y(n_1838)
);

AND2x6_ASAP7_75t_L g1839 ( 
.A(n_1667),
.B(n_1668),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1661),
.B(n_1141),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1662),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1698),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1651),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1625),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1616),
.B(n_1123),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_SL g1846 ( 
.A(n_1763),
.B(n_1126),
.Y(n_1846)
);

NAND2x1p5_ASAP7_75t_L g1847 ( 
.A(n_1661),
.B(n_1391),
.Y(n_1847)
);

INVx6_ASAP7_75t_L g1848 ( 
.A(n_1667),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1667),
.Y(n_1849)
);

AND2x6_ASAP7_75t_L g1850 ( 
.A(n_1668),
.B(n_1391),
.Y(n_1850)
);

NAND2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1668),
.B(n_1486),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_1698),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1675),
.B(n_1157),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1729),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1599),
.B(n_1128),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1714),
.A2(n_1132),
.B1(n_1133),
.B2(n_1131),
.Y(n_1856)
);

AND2x6_ASAP7_75t_L g1857 ( 
.A(n_1657),
.B(n_1486),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1729),
.Y(n_1858)
);

NAND2x1p5_ASAP7_75t_L g1859 ( 
.A(n_1677),
.B(n_1457),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1704),
.Y(n_1860)
);

INVx4_ASAP7_75t_SL g1861 ( 
.A(n_1654),
.Y(n_1861)
);

NAND3x1_ASAP7_75t_L g1862 ( 
.A(n_1696),
.B(n_1215),
.C(n_1206),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1621),
.B(n_1138),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1654),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1647),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1709),
.A2(n_1305),
.B1(n_1310),
.B2(n_1277),
.Y(n_1866)
);

INVx4_ASAP7_75t_L g1867 ( 
.A(n_1654),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1679),
.B(n_1228),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1664),
.B(n_1232),
.Y(n_1869)
);

OR2x6_ASAP7_75t_L g1870 ( 
.A(n_1689),
.B(n_1289),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1623),
.B(n_1488),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1599),
.B(n_1140),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1632),
.Y(n_1873)
);

INVx4_ASAP7_75t_L g1874 ( 
.A(n_1687),
.Y(n_1874)
);

NOR2x1p5_ASAP7_75t_L g1875 ( 
.A(n_1682),
.B(n_1147),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1712),
.B(n_993),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1624),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1687),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1717),
.B(n_993),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1648),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1610),
.B(n_1150),
.Y(n_1881)
);

NAND2xp33_ASAP7_75t_L g1882 ( 
.A(n_1629),
.B(n_1630),
.Y(n_1882)
);

INVx5_ASAP7_75t_L g1883 ( 
.A(n_1647),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1649),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1719),
.A2(n_1318),
.B1(n_1319),
.B2(n_1314),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1720),
.B(n_1200),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1670),
.B(n_1346),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1649),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1673),
.B(n_1379),
.Y(n_1889)
);

OR2x6_ASAP7_75t_L g1890 ( 
.A(n_1681),
.B(n_1004),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1674),
.B(n_1721),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1634),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1639),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1724),
.B(n_1156),
.Y(n_1894)
);

AND2x6_ASAP7_75t_L g1895 ( 
.A(n_1659),
.B(n_1663),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1640),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1692),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1728),
.B(n_1015),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1641),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1642),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1655),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1731),
.B(n_1161),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1644),
.B(n_1175),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1687),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1738),
.B(n_1176),
.Y(n_1905)
);

NOR2x1p5_ASAP7_75t_L g1906 ( 
.A(n_1684),
.B(n_1177),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1739),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1632),
.Y(n_1908)
);

NAND2x1p5_ASAP7_75t_L g1909 ( 
.A(n_1678),
.B(n_1355),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1741),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1596),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1627),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_1686),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1655),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1742),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1743),
.B(n_1015),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1665),
.B(n_1386),
.Y(n_1917)
);

INVx4_ASAP7_75t_L g1918 ( 
.A(n_1671),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1746),
.B(n_1182),
.Y(n_1919)
);

AND2x6_ASAP7_75t_L g1920 ( 
.A(n_1749),
.B(n_1410),
.Y(n_1920)
);

INVx4_ASAP7_75t_L g1921 ( 
.A(n_1671),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1751),
.B(n_1184),
.Y(n_1922)
);

BUFx3_ASAP7_75t_L g1923 ( 
.A(n_1758),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1759),
.Y(n_1924)
);

OR2x6_ASAP7_75t_L g1925 ( 
.A(n_1686),
.B(n_1098),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1760),
.Y(n_1926)
);

INVx4_ASAP7_75t_L g1927 ( 
.A(n_1686),
.Y(n_1927)
);

AND2x6_ASAP7_75t_L g1928 ( 
.A(n_1761),
.B(n_1116),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1697),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1605),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1601),
.B(n_1190),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1725),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1653),
.B(n_1191),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1683),
.B(n_1422),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1744),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_SL g1936 ( 
.A(n_1609),
.B(n_1192),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1705),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1666),
.B(n_1202),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1694),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1685),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1716),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1750),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1695),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1754),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1690),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1718),
.A2(n_1334),
.B1(n_1337),
.B2(n_1332),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1762),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1680),
.B(n_1205),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1691),
.B(n_1207),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1693),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1622),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1645),
.B(n_1438),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1635),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1603),
.Y(n_1954)
);

NAND3xp33_ASAP7_75t_L g1955 ( 
.A(n_1635),
.B(n_1223),
.C(n_1213),
.Y(n_1955)
);

INVx4_ASAP7_75t_L g1956 ( 
.A(n_1636),
.Y(n_1956)
);

NAND3x1_ASAP7_75t_L g1957 ( 
.A(n_1612),
.B(n_1469),
.C(n_1423),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1612),
.B(n_1083),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1612),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1638),
.B(n_1224),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1637),
.B(n_1068),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1638),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1732),
.B(n_1225),
.Y(n_1963)
);

INVx8_ASAP7_75t_L g1964 ( 
.A(n_1732),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1732),
.B(n_1229),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1756),
.B(n_1083),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1756),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1650),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1595),
.B(n_1083),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1604),
.Y(n_1970)
);

NAND2xp33_ASAP7_75t_L g1971 ( 
.A(n_1617),
.B(n_1209),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1723),
.B(n_1237),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1723),
.B(n_1242),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1618),
.B(n_1245),
.Y(n_1974)
);

INVx4_ASAP7_75t_L g1975 ( 
.A(n_1617),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1723),
.B(n_1246),
.Y(n_1976)
);

INVx4_ASAP7_75t_L g1977 ( 
.A(n_1617),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1604),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1615),
.B(n_1068),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1604),
.Y(n_1980)
);

INVx4_ASAP7_75t_L g1981 ( 
.A(n_1617),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1626),
.Y(n_1982)
);

INVx6_ASAP7_75t_L g1983 ( 
.A(n_1736),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1595),
.B(n_1103),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1736),
.Y(n_1985)
);

AND2x6_ASAP7_75t_L g1986 ( 
.A(n_1618),
.B(n_1116),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1595),
.B(n_1103),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1615),
.B(n_1092),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1652),
.B(n_1249),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1626),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1604),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1652),
.B(n_1473),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1626),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1604),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1626),
.Y(n_1995)
);

NOR2x1p5_ASAP7_75t_L g1996 ( 
.A(n_1617),
.B(n_1252),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1736),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1604),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1791),
.B(n_1470),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1813),
.B(n_1253),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1774),
.Y(n_2001)
);

NAND2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1780),
.B(n_1006),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1992),
.B(n_1244),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1794),
.B(n_1111),
.Y(n_2004)
);

OR2x6_ASAP7_75t_L g2005 ( 
.A(n_1983),
.B(n_1098),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1801),
.B(n_1257),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1817),
.Y(n_2007)
);

AO22x2_ASAP7_75t_L g2008 ( 
.A1(n_1784),
.A2(n_1266),
.B1(n_1382),
.B2(n_1248),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1804),
.A2(n_1269),
.B1(n_1270),
.B2(n_1258),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1800),
.B(n_1812),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1936),
.A2(n_1276),
.B1(n_1280),
.B2(n_1275),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1774),
.B(n_1282),
.Y(n_2012)
);

CKINVDCx20_ASAP7_75t_R g2013 ( 
.A(n_1769),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1820),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1777),
.B(n_1244),
.Y(n_2015)
);

AO22x2_ASAP7_75t_L g2016 ( 
.A1(n_1777),
.A2(n_1429),
.B1(n_989),
.B2(n_995),
.Y(n_2016)
);

OAI221xp5_ASAP7_75t_L g2017 ( 
.A1(n_1822),
.A2(n_1292),
.B1(n_1293),
.B2(n_1290),
.C(n_1285),
.Y(n_2017)
);

AO22x2_ASAP7_75t_L g2018 ( 
.A1(n_1869),
.A2(n_996),
.B1(n_1000),
.B2(n_981),
.Y(n_2018)
);

NAND2x1p5_ASAP7_75t_L g2019 ( 
.A(n_1831),
.B(n_1092),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1818),
.A2(n_1796),
.B1(n_1984),
.B2(n_1969),
.Y(n_2020)
);

OAI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_1828),
.A2(n_1308),
.B1(n_1316),
.B2(n_1300),
.C(n_1296),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1821),
.B(n_1007),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1877),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1892),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1893),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1985),
.Y(n_2026)
);

NAND2x1p5_ASAP7_75t_L g2027 ( 
.A(n_1997),
.B(n_1841),
.Y(n_2027)
);

NAND2x1p5_ASAP7_75t_L g2028 ( 
.A(n_1795),
.B(n_1127),
.Y(n_2028)
);

AO22x2_ASAP7_75t_L g2029 ( 
.A1(n_1887),
.A2(n_1014),
.B1(n_1029),
.B2(n_1013),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1896),
.Y(n_2030)
);

BUFx8_ASAP7_75t_L g2031 ( 
.A(n_1790),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1899),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1801),
.B(n_1768),
.Y(n_2033)
);

AO22x2_ASAP7_75t_L g2034 ( 
.A1(n_1889),
.A2(n_1051),
.B1(n_1058),
.B2(n_1032),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1900),
.Y(n_2035)
);

AO22x2_ASAP7_75t_L g2036 ( 
.A1(n_1868),
.A2(n_1077),
.B1(n_1104),
.B2(n_1073),
.Y(n_2036)
);

BUFx8_ASAP7_75t_L g2037 ( 
.A(n_1939),
.Y(n_2037)
);

NAND2x1p5_ASAP7_75t_L g2038 ( 
.A(n_1975),
.B(n_1183),
.Y(n_2038)
);

AO22x2_ASAP7_75t_L g2039 ( 
.A1(n_1826),
.A2(n_1108),
.B1(n_1119),
.B2(n_1113),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1764),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1765),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1766),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1772),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1974),
.B(n_1320),
.Y(n_2044)
);

NAND2x1p5_ASAP7_75t_L g2045 ( 
.A(n_1977),
.B(n_1183),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1773),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1970),
.Y(n_2047)
);

AO22x2_ASAP7_75t_L g2048 ( 
.A1(n_1826),
.A2(n_1142),
.B1(n_1145),
.B2(n_1136),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_1859),
.Y(n_2049)
);

NAND2x1p5_ASAP7_75t_L g2050 ( 
.A(n_1981),
.B(n_1250),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1772),
.Y(n_2051)
);

NAND2x1p5_ASAP7_75t_L g2052 ( 
.A(n_1878),
.B(n_1874),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1870),
.B(n_1149),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1982),
.Y(n_2054)
);

INVxp33_ASAP7_75t_SL g2055 ( 
.A(n_1797),
.Y(n_2055)
);

BUFx24_ASAP7_75t_SL g2056 ( 
.A(n_1856),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1847),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1982),
.Y(n_2058)
);

OAI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_1828),
.A2(n_1325),
.B1(n_1326),
.B2(n_1324),
.C(n_1322),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_L g2060 ( 
.A(n_1845),
.B(n_1340),
.C(n_1328),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1978),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1980),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1990),
.Y(n_2063)
);

AO22x2_ASAP7_75t_L g2064 ( 
.A1(n_1843),
.A2(n_1154),
.B1(n_1163),
.B2(n_1153),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1823),
.B(n_1366),
.Y(n_2065)
);

NAND2x1p5_ASAP7_75t_L g2066 ( 
.A(n_1904),
.B(n_1250),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1987),
.A2(n_1360),
.B1(n_1361),
.B2(n_1359),
.Y(n_2067)
);

AO22x2_ASAP7_75t_L g2068 ( 
.A1(n_1886),
.A2(n_1168),
.B1(n_1169),
.B2(n_1166),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1991),
.Y(n_2069)
);

AO22x2_ASAP7_75t_L g2070 ( 
.A1(n_1886),
.A2(n_1179),
.B1(n_1189),
.B2(n_1170),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1860),
.A2(n_1370),
.B1(n_1374),
.B2(n_1364),
.Y(n_2071)
);

NAND2x1p5_ASAP7_75t_L g2072 ( 
.A(n_1849),
.B(n_1278),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1994),
.Y(n_2073)
);

AO22x2_ASAP7_75t_L g2074 ( 
.A1(n_1917),
.A2(n_1853),
.B1(n_1830),
.B2(n_1785),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1909),
.B(n_1406),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1998),
.Y(n_2076)
);

NAND2xp33_ASAP7_75t_L g2077 ( 
.A(n_1819),
.B(n_1416),
.Y(n_2077)
);

AO22x2_ASAP7_75t_L g2078 ( 
.A1(n_1806),
.A2(n_1198),
.B1(n_1199),
.B2(n_1196),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_1873),
.Y(n_2079)
);

AO22x2_ASAP7_75t_L g2080 ( 
.A1(n_1808),
.A2(n_1217),
.B1(n_1218),
.B2(n_1203),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1833),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_1782),
.A2(n_1395),
.B1(n_1396),
.B2(n_1394),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1834),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1835),
.Y(n_2084)
);

INVxp67_ASAP7_75t_L g2085 ( 
.A(n_1908),
.Y(n_2085)
);

OR2x6_ASAP7_75t_L g2086 ( 
.A(n_1983),
.B(n_1102),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1990),
.Y(n_2087)
);

NAND2x1p5_ASAP7_75t_L g2088 ( 
.A(n_1849),
.B(n_1278),
.Y(n_2088)
);

NAND2xp33_ASAP7_75t_L g2089 ( 
.A(n_1819),
.B(n_1421),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1894),
.A2(n_1342),
.B(n_1389),
.C(n_1352),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1844),
.Y(n_2091)
);

NAND2x1p5_ASAP7_75t_L g2092 ( 
.A(n_1770),
.B(n_1342),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1993),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1918),
.B(n_1405),
.Y(n_2094)
);

AO22x2_ASAP7_75t_L g2095 ( 
.A1(n_1809),
.A2(n_1238),
.B1(n_1251),
.B2(n_1220),
.Y(n_2095)
);

AO22x2_ASAP7_75t_L g2096 ( 
.A1(n_1934),
.A2(n_1262),
.B1(n_1268),
.B2(n_1261),
.Y(n_2096)
);

NAND2x1p5_ASAP7_75t_L g2097 ( 
.A(n_1771),
.B(n_1389),
.Y(n_2097)
);

NAND2x1p5_ASAP7_75t_L g2098 ( 
.A(n_1968),
.B(n_1339),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1880),
.B(n_1923),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_1798),
.A2(n_1432),
.B1(n_1439),
.B2(n_1427),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_1920),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_1925),
.Y(n_2102)
);

AO22x2_ASAP7_75t_L g2103 ( 
.A1(n_1957),
.A2(n_1273),
.B1(n_1283),
.B2(n_1272),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1993),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1995),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1875),
.B(n_1284),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1907),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1910),
.Y(n_2108)
);

AO22x2_ASAP7_75t_L g2109 ( 
.A1(n_1779),
.A2(n_1307),
.B1(n_1309),
.B2(n_1298),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1915),
.Y(n_2110)
);

OAI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_1793),
.A2(n_1471),
.B1(n_1474),
.B2(n_1461),
.C(n_1449),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_1927),
.B(n_1376),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_SL g2113 ( 
.A(n_1789),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1924),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1926),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1930),
.B(n_1264),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1906),
.B(n_1327),
.Y(n_2117)
);

AO22x2_ASAP7_75t_L g2118 ( 
.A1(n_1783),
.A2(n_1861),
.B1(n_1827),
.B2(n_1788),
.Y(n_2118)
);

AO22x2_ASAP7_75t_L g2119 ( 
.A1(n_1861),
.A2(n_1356),
.B1(n_1363),
.B2(n_1354),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_1925),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1807),
.B(n_1476),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1882),
.Y(n_2122)
);

AOI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_1799),
.A2(n_976),
.B1(n_979),
.B2(n_975),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1814),
.B(n_1491),
.Y(n_2124)
);

BUFx10_ASAP7_75t_L g2125 ( 
.A(n_1996),
.Y(n_2125)
);

AO22x2_ASAP7_75t_L g2126 ( 
.A1(n_1897),
.A2(n_1373),
.B1(n_1378),
.B2(n_1368),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_SL g2127 ( 
.A(n_1950),
.B(n_1264),
.Y(n_2127)
);

AO22x2_ASAP7_75t_L g2128 ( 
.A1(n_1805),
.A2(n_1383),
.B1(n_1407),
.B2(n_1380),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1824),
.B(n_1479),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1832),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1865),
.Y(n_2131)
);

CKINVDCx16_ASAP7_75t_R g2132 ( 
.A(n_1811),
.Y(n_2132)
);

BUFx8_ASAP7_75t_L g2133 ( 
.A(n_1945),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1972),
.B(n_1487),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1930),
.B(n_1264),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1952),
.Y(n_2136)
);

BUFx8_ASAP7_75t_L g2137 ( 
.A(n_1888),
.Y(n_2137)
);

NAND3xp33_ASAP7_75t_SL g2138 ( 
.A(n_1940),
.B(n_1943),
.C(n_1913),
.Y(n_2138)
);

AO22x2_ASAP7_75t_L g2139 ( 
.A1(n_1815),
.A2(n_1412),
.B1(n_1440),
.B2(n_1408),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1952),
.Y(n_2140)
);

AO22x2_ASAP7_75t_L g2141 ( 
.A1(n_1816),
.A2(n_1446),
.B1(n_1450),
.B2(n_1441),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_SL g2142 ( 
.A1(n_1842),
.A2(n_985),
.B1(n_986),
.B2(n_984),
.Y(n_2142)
);

AO22x2_ASAP7_75t_L g2143 ( 
.A1(n_1854),
.A2(n_1483),
.B1(n_1492),
.B2(n_1454),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1837),
.B(n_1274),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1836),
.B(n_1867),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1876),
.B(n_1017),
.Y(n_2146)
);

INVxp67_ASAP7_75t_SL g2147 ( 
.A(n_1995),
.Y(n_2147)
);

NAND2x1p5_ASAP7_75t_L g2148 ( 
.A(n_1921),
.B(n_1385),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1958),
.Y(n_2149)
);

CKINVDCx11_ASAP7_75t_R g2150 ( 
.A(n_1852),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1890),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_1920),
.A2(n_1388),
.B1(n_1390),
.B2(n_1387),
.Y(n_2152)
);

AO22x2_ASAP7_75t_L g2153 ( 
.A1(n_1858),
.A2(n_1399),
.B1(n_1403),
.B2(n_1392),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1966),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1863),
.B(n_987),
.Y(n_2155)
);

NAND2x1p5_ASAP7_75t_L g2156 ( 
.A(n_1883),
.B(n_1404),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1973),
.B(n_1494),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1976),
.B(n_1495),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1776),
.Y(n_2159)
);

NAND2x1p5_ASAP7_75t_L g2160 ( 
.A(n_1883),
.B(n_1409),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1848),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_1839),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1781),
.Y(n_2163)
);

BUFx2_ASAP7_75t_L g2164 ( 
.A(n_1920),
.Y(n_2164)
);

OAI221xp5_ASAP7_75t_L g2165 ( 
.A1(n_1866),
.A2(n_1005),
.B1(n_1009),
.B2(n_998),
.C(n_991),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1879),
.B(n_1274),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_1898),
.B(n_1036),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1916),
.B(n_1274),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1871),
.B(n_1903),
.Y(n_2169)
);

AO22x2_ASAP7_75t_L g2170 ( 
.A1(n_1979),
.A2(n_1420),
.B1(n_1426),
.B2(n_1417),
.Y(n_2170)
);

NAND2x1p5_ASAP7_75t_L g2171 ( 
.A(n_1888),
.B(n_1430),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1825),
.B(n_1431),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1802),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1786),
.B(n_1443),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1947),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_1885),
.A2(n_1459),
.B1(n_1475),
.B2(n_1447),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1902),
.B(n_1011),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1905),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1855),
.A2(n_1021),
.B1(n_1023),
.B2(n_1020),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_1988),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1919),
.Y(n_2181)
);

AO22x2_ASAP7_75t_L g2182 ( 
.A1(n_1884),
.A2(n_1109),
.B1(n_1162),
.B2(n_1102),
.Y(n_2182)
);

BUFx12f_ASAP7_75t_L g2183 ( 
.A(n_1890),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1922),
.B(n_1297),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1840),
.B(n_1297),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_1989),
.B(n_1046),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1846),
.Y(n_2187)
);

NOR2xp67_ASAP7_75t_L g2188 ( 
.A(n_1767),
.B(n_3),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1787),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1872),
.B(n_1297),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_1810),
.B(n_1084),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1960),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1891),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1851),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1881),
.B(n_1321),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1901),
.B(n_1031),
.Y(n_2196)
);

AOI22xp5_ASAP7_75t_SL g2197 ( 
.A1(n_1911),
.A2(n_1041),
.B1(n_1043),
.B2(n_1034),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1775),
.Y(n_2198)
);

OAI221xp5_ASAP7_75t_L g2199 ( 
.A1(n_1792),
.A2(n_1047),
.B1(n_1055),
.B2(n_1045),
.C(n_1044),
.Y(n_2199)
);

INVxp67_ASAP7_75t_SL g2200 ( 
.A(n_1803),
.Y(n_2200)
);

AO22x2_ASAP7_75t_L g2201 ( 
.A1(n_1862),
.A2(n_1162),
.B1(n_1167),
.B2(n_1109),
.Y(n_2201)
);

NAND2x1p5_ASAP7_75t_L g2202 ( 
.A(n_1901),
.B(n_1914),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1803),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1929),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_1838),
.B(n_1056),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1937),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1949),
.A2(n_1059),
.B1(n_1067),
.B2(n_1060),
.Y(n_2207)
);

NAND3xp33_ASAP7_75t_SL g2208 ( 
.A(n_1912),
.B(n_1931),
.C(n_1946),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_SL g2209 ( 
.A(n_1839),
.B(n_1321),
.Y(n_2209)
);

AO22x2_ASAP7_75t_L g2210 ( 
.A1(n_1864),
.A2(n_1397),
.B1(n_1442),
.B2(n_1219),
.Y(n_2210)
);

AO22x2_ASAP7_75t_L g2211 ( 
.A1(n_1948),
.A2(n_1442),
.B1(n_1444),
.B2(n_1321),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1941),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_1914),
.B(n_1455),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_1767),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1829),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1778),
.B(n_1096),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1963),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1965),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1961),
.Y(n_2219)
);

INVx2_ASAP7_75t_SL g2220 ( 
.A(n_1778),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1850),
.Y(n_2221)
);

AO22x2_ASAP7_75t_L g2222 ( 
.A1(n_1857),
.A2(n_1444),
.B1(n_1455),
.B2(n_6),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_1857),
.B(n_1455),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_1895),
.B(n_1118),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1895),
.B(n_1124),
.Y(n_2225)
);

AO22x2_ASAP7_75t_L g2226 ( 
.A1(n_1839),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1933),
.Y(n_2227)
);

NAND2x1p5_ASAP7_75t_L g2228 ( 
.A(n_1956),
.B(n_1155),
.Y(n_2228)
);

AO22x2_ASAP7_75t_L g2229 ( 
.A1(n_1850),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_1986),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1932),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1935),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1942),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_1955),
.B(n_1088),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_1938),
.B(n_1099),
.Y(n_2235)
);

INVx2_ASAP7_75t_SL g2236 ( 
.A(n_1986),
.Y(n_2236)
);

CKINVDCx14_ASAP7_75t_R g2237 ( 
.A(n_1928),
.Y(n_2237)
);

AO22x2_ASAP7_75t_L g2238 ( 
.A1(n_1944),
.A2(n_8),
.B1(n_4),
.B2(n_7),
.Y(n_2238)
);

INVxp67_ASAP7_75t_L g2239 ( 
.A(n_1928),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_1967),
.Y(n_2240)
);

AO22x2_ASAP7_75t_L g2241 ( 
.A1(n_1971),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_1964),
.B(n_1106),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1954),
.Y(n_2243)
);

AO22x2_ASAP7_75t_L g2244 ( 
.A1(n_1959),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_1951),
.B(n_1135),
.Y(n_2245)
);

AO22x2_ASAP7_75t_L g2246 ( 
.A1(n_1962),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_1951),
.B(n_1137),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_1953),
.B(n_1158),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1992),
.Y(n_2249)
);

AO22x2_ASAP7_75t_L g2250 ( 
.A1(n_1992),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1992),
.Y(n_2251)
);

NAND2x1p5_ASAP7_75t_L g2252 ( 
.A(n_1780),
.B(n_1155),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1769),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1992),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1992),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_1791),
.B(n_1180),
.Y(n_2256)
);

AO22x2_ASAP7_75t_L g2257 ( 
.A1(n_1992),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1992),
.Y(n_2258)
);

AO22x2_ASAP7_75t_L g2259 ( 
.A1(n_1992),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1992),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_SL g2261 ( 
.A1(n_1842),
.A2(n_1159),
.B1(n_1172),
.B2(n_1160),
.Y(n_2261)
);

OAI21xp33_ASAP7_75t_L g2262 ( 
.A1(n_1992),
.A2(n_1467),
.B(n_1465),
.Y(n_2262)
);

AO22x2_ASAP7_75t_L g2263 ( 
.A1(n_1992),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1992),
.B(n_1181),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1992),
.Y(n_2265)
);

INVx4_ASAP7_75t_L g2266 ( 
.A(n_1983),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1992),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1992),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1992),
.Y(n_2269)
);

NAND3xp33_ASAP7_75t_SL g2270 ( 
.A(n_1784),
.B(n_1480),
.C(n_1472),
.Y(n_2270)
);

HB1xp67_ASAP7_75t_L g2271 ( 
.A(n_1774),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1849),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1992),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1992),
.B(n_1185),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2011),
.B(n_1482),
.Y(n_2275)
);

NAND2xp33_ASAP7_75t_SL g2276 ( 
.A(n_2101),
.B(n_1260),
.Y(n_2276)
);

NAND2xp33_ASAP7_75t_SL g2277 ( 
.A(n_2164),
.B(n_2272),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2014),
.B(n_1484),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2127),
.B(n_1485),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2208),
.B(n_1186),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2001),
.B(n_1490),
.Y(n_2281)
);

NAND2xp33_ASAP7_75t_SL g2282 ( 
.A(n_2272),
.B(n_1260),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2033),
.B(n_1188),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2178),
.B(n_15),
.Y(n_2284)
);

NAND2xp33_ASAP7_75t_SL g2285 ( 
.A(n_2221),
.B(n_1260),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2249),
.B(n_1193),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2049),
.B(n_1445),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2264),
.B(n_1448),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2274),
.B(n_1481),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2251),
.B(n_1489),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2254),
.B(n_1195),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2255),
.B(n_1452),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2258),
.B(n_1201),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2260),
.B(n_1458),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2271),
.B(n_1204),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2265),
.B(n_1208),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2267),
.B(n_1210),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_2268),
.B(n_1468),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2181),
.B(n_16),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2269),
.B(n_1493),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_2273),
.B(n_1216),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2002),
.B(n_1414),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2209),
.B(n_1415),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2224),
.B(n_1419),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2225),
.B(n_1425),
.Y(n_2305)
);

AND2x2_ASAP7_75t_SL g2306 ( 
.A(n_2077),
.B(n_1299),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2012),
.B(n_1428),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2009),
.B(n_1433),
.Y(n_2308)
);

NAND2xp33_ASAP7_75t_SL g2309 ( 
.A(n_2152),
.B(n_1299),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2120),
.B(n_1435),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2148),
.B(n_1222),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2136),
.B(n_1227),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2140),
.B(n_1231),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2003),
.B(n_1233),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2082),
.B(n_1460),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2098),
.B(n_1462),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2071),
.B(n_1234),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2000),
.B(n_1236),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2006),
.B(n_1365),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2112),
.B(n_1367),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2116),
.B(n_1371),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2135),
.B(n_1384),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2015),
.B(n_1393),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2156),
.B(n_1401),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2160),
.B(n_1239),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_SL g2326 ( 
.A(n_2040),
.B(n_1306),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2094),
.B(n_1413),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_2223),
.B(n_1434),
.Y(n_2328)
);

NAND2xp33_ASAP7_75t_SL g2329 ( 
.A(n_2122),
.B(n_1306),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2107),
.B(n_2108),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2248),
.B(n_1240),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_2262),
.B(n_2169),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2110),
.B(n_1241),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2019),
.B(n_1247),
.Y(n_2334)
);

NAND2xp33_ASAP7_75t_SL g2335 ( 
.A(n_2187),
.B(n_1254),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2055),
.B(n_1255),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2067),
.B(n_1263),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_SL g2338 ( 
.A(n_2037),
.B(n_1344),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2016),
.B(n_2068),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2133),
.B(n_1345),
.Y(n_2340)
);

NAND2xp33_ASAP7_75t_SL g2341 ( 
.A(n_2113),
.B(n_1265),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2151),
.B(n_2020),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_2146),
.B(n_1349),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2114),
.B(n_2115),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2167),
.B(n_1357),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2186),
.B(n_1358),
.Y(n_2346)
);

NAND2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2057),
.B(n_1271),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2234),
.B(n_2252),
.Y(n_2348)
);

NAND2xp33_ASAP7_75t_SL g2349 ( 
.A(n_2075),
.B(n_1279),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2162),
.B(n_1281),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_SL g2351 ( 
.A(n_2102),
.B(n_1286),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2007),
.B(n_1287),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2016),
.B(n_1288),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_SL g2354 ( 
.A(n_2266),
.B(n_2121),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_2079),
.B(n_1291),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2085),
.B(n_1294),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2261),
.B(n_1323),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2171),
.B(n_1302),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2004),
.B(n_1330),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2240),
.B(n_1333),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2242),
.B(n_1336),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2028),
.B(n_1303),
.Y(n_2362)
);

NAND2xp33_ASAP7_75t_SL g2363 ( 
.A(n_2044),
.B(n_1304),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2038),
.B(n_1312),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_2045),
.B(n_1313),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2050),
.B(n_1348),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2100),
.B(n_1437),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2068),
.B(n_1209),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2216),
.B(n_1306),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2245),
.B(n_1338),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2247),
.B(n_1338),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2197),
.B(n_2123),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2144),
.B(n_1436),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2166),
.B(n_1436),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2168),
.B(n_1436),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2053),
.B(n_1464),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2124),
.B(n_1295),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2129),
.B(n_1295),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_2132),
.B(n_1295),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2065),
.B(n_2183),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_2227),
.B(n_16),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_2256),
.B(n_2191),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2060),
.B(n_1451),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2184),
.B(n_1451),
.Y(n_2384)
);

NAND2xp33_ASAP7_75t_SL g2385 ( 
.A(n_2230),
.B(n_1052),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2142),
.B(n_1451),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2134),
.B(n_2157),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2207),
.B(n_1451),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2190),
.B(n_2195),
.Y(n_2389)
);

NAND2xp33_ASAP7_75t_SL g2390 ( 
.A(n_2023),
.B(n_1052),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2158),
.B(n_1451),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_SL g2392 ( 
.A(n_2024),
.B(n_1052),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2179),
.B(n_1194),
.Y(n_2393)
);

NAND2xp33_ASAP7_75t_SL g2394 ( 
.A(n_2025),
.B(n_1214),
.Y(n_2394)
);

NAND2xp33_ASAP7_75t_SL g2395 ( 
.A(n_2030),
.B(n_1214),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2070),
.B(n_17),
.Y(n_2396)
);

NAND2xp33_ASAP7_75t_SL g2397 ( 
.A(n_2032),
.B(n_1214),
.Y(n_2397)
);

NAND2xp33_ASAP7_75t_SL g2398 ( 
.A(n_2035),
.B(n_1329),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2192),
.B(n_17),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2052),
.B(n_2106),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2117),
.B(n_1362),
.Y(n_2401)
);

NAND2xp33_ASAP7_75t_SL g2402 ( 
.A(n_2236),
.B(n_1362),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2070),
.B(n_18),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2137),
.B(n_1456),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2159),
.B(n_19),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2125),
.B(n_2235),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_1999),
.B(n_20),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_2185),
.B(n_20),
.Y(n_2408)
);

NAND2xp33_ASAP7_75t_SL g2409 ( 
.A(n_2043),
.B(n_19),
.Y(n_2409)
);

NAND2xp33_ASAP7_75t_SL g2410 ( 
.A(n_2051),
.B(n_20),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2056),
.B(n_2172),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2196),
.B(n_22),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2188),
.B(n_22),
.Y(n_2413)
);

NAND2xp33_ASAP7_75t_SL g2414 ( 
.A(n_2054),
.B(n_21),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_SL g2415 ( 
.A(n_2149),
.B(n_22),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2154),
.B(n_2099),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2220),
.B(n_23),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_SL g2418 ( 
.A(n_2194),
.B(n_23),
.Y(n_2418)
);

NAND2xp33_ASAP7_75t_SL g2419 ( 
.A(n_2058),
.B(n_21),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2174),
.B(n_21),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2022),
.B(n_25),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2177),
.B(n_26),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2163),
.B(n_24),
.Y(n_2423)
);

NAND2xp33_ASAP7_75t_SL g2424 ( 
.A(n_2063),
.B(n_24),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_SL g2425 ( 
.A(n_2041),
.B(n_27),
.Y(n_2425)
);

NAND2xp33_ASAP7_75t_SL g2426 ( 
.A(n_2087),
.B(n_24),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_2042),
.B(n_29),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2046),
.B(n_29),
.Y(n_2428)
);

NAND2xp33_ASAP7_75t_L g2429 ( 
.A(n_2093),
.B(n_29),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_SL g2430 ( 
.A(n_2047),
.B(n_30),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2126),
.B(n_28),
.Y(n_2431)
);

NAND2xp33_ASAP7_75t_SL g2432 ( 
.A(n_2104),
.B(n_28),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_SL g2433 ( 
.A(n_2061),
.B(n_30),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_2062),
.B(n_31),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2126),
.B(n_28),
.Y(n_2435)
);

NAND2xp33_ASAP7_75t_SL g2436 ( 
.A(n_2069),
.B(n_32),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2039),
.B(n_32),
.Y(n_2437)
);

NAND2xp33_ASAP7_75t_SL g2438 ( 
.A(n_2073),
.B(n_32),
.Y(n_2438)
);

NAND2xp33_ASAP7_75t_SL g2439 ( 
.A(n_2076),
.B(n_2084),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2091),
.B(n_34),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2039),
.B(n_33),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2048),
.B(n_33),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2048),
.B(n_35),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2170),
.B(n_35),
.Y(n_2444)
);

NAND2xp33_ASAP7_75t_SL g2445 ( 
.A(n_2175),
.B(n_35),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2092),
.B(n_38),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2097),
.B(n_38),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2180),
.B(n_39),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2239),
.B(n_39),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2072),
.B(n_39),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2088),
.B(n_40),
.Y(n_2451)
);

NAND2xp33_ASAP7_75t_SL g2452 ( 
.A(n_2204),
.B(n_37),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2170),
.B(n_40),
.Y(n_2453)
);

NAND2xp33_ASAP7_75t_SL g2454 ( 
.A(n_2206),
.B(n_40),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2018),
.B(n_41),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2066),
.B(n_42),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_2212),
.B(n_42),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2026),
.B(n_42),
.Y(n_2458)
);

NAND2xp33_ASAP7_75t_SL g2459 ( 
.A(n_2237),
.B(n_41),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2253),
.B(n_44),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2176),
.B(n_44),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2228),
.B(n_45),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2214),
.B(n_45),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2189),
.B(n_45),
.Y(n_2464)
);

NAND2xp33_ASAP7_75t_SL g2465 ( 
.A(n_2013),
.B(n_43),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2010),
.B(n_46),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2202),
.B(n_46),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2213),
.B(n_46),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_2027),
.B(n_47),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2130),
.B(n_47),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2193),
.B(n_48),
.Y(n_2471)
);

NAND2xp33_ASAP7_75t_SL g2472 ( 
.A(n_2089),
.B(n_48),
.Y(n_2472)
);

NAND2xp33_ASAP7_75t_SL g2473 ( 
.A(n_2205),
.B(n_49),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2198),
.B(n_52),
.Y(n_2474)
);

NAND2xp33_ASAP7_75t_SL g2475 ( 
.A(n_2155),
.B(n_50),
.Y(n_2475)
);

NAND2xp33_ASAP7_75t_SL g2476 ( 
.A(n_2145),
.B(n_50),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_2217),
.B(n_50),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2161),
.B(n_55),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2081),
.B(n_54),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2083),
.B(n_55),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2218),
.B(n_56),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2219),
.B(n_56),
.Y(n_2482)
);

NAND2xp33_ASAP7_75t_SL g2483 ( 
.A(n_2105),
.B(n_55),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2018),
.B(n_56),
.Y(n_2484)
);

NAND2xp33_ASAP7_75t_SL g2485 ( 
.A(n_2203),
.B(n_57),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2029),
.B(n_57),
.Y(n_2486)
);

NAND2xp33_ASAP7_75t_SL g2487 ( 
.A(n_2215),
.B(n_58),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2131),
.B(n_59),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2182),
.B(n_58),
.Y(n_2489)
);

NAND2xp33_ASAP7_75t_SL g2490 ( 
.A(n_2173),
.B(n_58),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2182),
.B(n_60),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2243),
.B(n_62),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2109),
.B(n_61),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2090),
.B(n_62),
.Y(n_2494)
);

NAND2xp33_ASAP7_75t_SL g2495 ( 
.A(n_2222),
.B(n_61),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_2231),
.B(n_64),
.Y(n_2496)
);

NAND2xp33_ASAP7_75t_SL g2497 ( 
.A(n_2222),
.B(n_61),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2232),
.B(n_65),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2109),
.B(n_2153),
.Y(n_2499)
);

NAND2xp33_ASAP7_75t_SL g2500 ( 
.A(n_2233),
.B(n_64),
.Y(n_2500)
);

XNOR2x2_ASAP7_75t_L g2501 ( 
.A(n_2008),
.B(n_65),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2153),
.B(n_65),
.Y(n_2502)
);

NAND2xp33_ASAP7_75t_SL g2503 ( 
.A(n_2119),
.B(n_67),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2064),
.B(n_2078),
.Y(n_2504)
);

NAND2xp33_ASAP7_75t_SL g2505 ( 
.A(n_2119),
.B(n_67),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2064),
.B(n_67),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2147),
.B(n_69),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2029),
.B(n_68),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2080),
.B(n_69),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2080),
.B(n_2095),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2031),
.B(n_2200),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2034),
.B(n_70),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2095),
.B(n_70),
.Y(n_2513)
);

NAND2xp33_ASAP7_75t_SL g2514 ( 
.A(n_2226),
.B(n_71),
.Y(n_2514)
);

NAND2xp33_ASAP7_75t_SL g2515 ( 
.A(n_2226),
.B(n_71),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_2021),
.B(n_71),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2270),
.B(n_74),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2138),
.B(n_74),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2059),
.B(n_75),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2074),
.B(n_76),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_2005),
.B(n_76),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2005),
.B(n_77),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2086),
.B(n_77),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_2086),
.B(n_77),
.Y(n_2524)
);

NAND2xp33_ASAP7_75t_SL g2525 ( 
.A(n_2229),
.B(n_73),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2034),
.B(n_78),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2036),
.B(n_2008),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_2036),
.B(n_78),
.Y(n_2528)
);

AND2x4_ASAP7_75t_L g2529 ( 
.A(n_2118),
.B(n_73),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2210),
.B(n_78),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2128),
.B(n_73),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2210),
.B(n_80),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2017),
.B(n_80),
.Y(n_2533)
);

NAND2xp33_ASAP7_75t_SL g2534 ( 
.A(n_2229),
.B(n_79),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2128),
.B(n_79),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2118),
.B(n_81),
.Y(n_2536)
);

NAND2xp33_ASAP7_75t_SL g2537 ( 
.A(n_2250),
.B(n_79),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2111),
.B(n_83),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2139),
.B(n_83),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2139),
.B(n_83),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2141),
.B(n_84),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2141),
.B(n_84),
.Y(n_2542)
);

NAND2xp33_ASAP7_75t_SL g2543 ( 
.A(n_2250),
.B(n_82),
.Y(n_2543)
);

AND2x4_ASAP7_75t_L g2544 ( 
.A(n_2257),
.B(n_84),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2096),
.B(n_85),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2096),
.B(n_85),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_2103),
.B(n_87),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_SL g2548 ( 
.A(n_2257),
.B(n_86),
.Y(n_2548)
);

NAND2xp33_ASAP7_75t_SL g2549 ( 
.A(n_2259),
.B(n_87),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2259),
.B(n_88),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2143),
.B(n_89),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2103),
.B(n_90),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2143),
.B(n_89),
.Y(n_2553)
);

NAND2xp33_ASAP7_75t_SL g2554 ( 
.A(n_2263),
.B(n_90),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2211),
.B(n_90),
.Y(n_2555)
);

NAND2xp33_ASAP7_75t_L g2556 ( 
.A(n_2211),
.B(n_92),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2165),
.B(n_92),
.Y(n_2557)
);

NAND2xp33_ASAP7_75t_SL g2558 ( 
.A(n_2263),
.B(n_91),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2199),
.B(n_92),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2201),
.B(n_91),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2241),
.B(n_94),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2241),
.B(n_94),
.Y(n_2562)
);

NAND2xp33_ASAP7_75t_SL g2563 ( 
.A(n_2238),
.B(n_2246),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2244),
.B(n_94),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2244),
.B(n_95),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_SL g2566 ( 
.A(n_2150),
.B(n_93),
.Y(n_2566)
);

NAND2xp33_ASAP7_75t_SL g2567 ( 
.A(n_2101),
.B(n_93),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2033),
.B(n_95),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2208),
.B(n_95),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2011),
.B(n_97),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2011),
.B(n_97),
.Y(n_2571)
);

NAND2xp33_ASAP7_75t_SL g2572 ( 
.A(n_2101),
.B(n_96),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2011),
.B(n_97),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2011),
.B(n_98),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2011),
.B(n_99),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2011),
.B(n_99),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_2011),
.B(n_99),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2011),
.B(n_100),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2011),
.B(n_100),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_SL g2580 ( 
.A(n_2011),
.B(n_101),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2011),
.B(n_102),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2011),
.B(n_102),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2033),
.B(n_96),
.Y(n_2583)
);

NAND2xp33_ASAP7_75t_SL g2584 ( 
.A(n_2101),
.B(n_102),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2033),
.B(n_103),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2011),
.B(n_104),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2033),
.B(n_104),
.Y(n_2587)
);

NAND2xp33_ASAP7_75t_SL g2588 ( 
.A(n_2101),
.B(n_104),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_2011),
.B(n_106),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2011),
.B(n_106),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_2011),
.B(n_106),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2033),
.B(n_105),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_SL g2593 ( 
.A(n_2011),
.B(n_107),
.Y(n_2593)
);

NAND2xp33_ASAP7_75t_SL g2594 ( 
.A(n_2101),
.B(n_105),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2033),
.B(n_107),
.Y(n_2595)
);

NAND2xp33_ASAP7_75t_SL g2596 ( 
.A(n_2101),
.B(n_107),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_SL g2597 ( 
.A(n_2011),
.B(n_109),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2011),
.B(n_109),
.Y(n_2598)
);

NAND2xp33_ASAP7_75t_SL g2599 ( 
.A(n_2101),
.B(n_108),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_2011),
.B(n_110),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2033),
.B(n_108),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2178),
.B(n_111),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_2011),
.B(n_112),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_SL g2604 ( 
.A(n_2011),
.B(n_113),
.Y(n_2604)
);

NAND2xp33_ASAP7_75t_SL g2605 ( 
.A(n_2101),
.B(n_111),
.Y(n_2605)
);

NAND2xp33_ASAP7_75t_SL g2606 ( 
.A(n_2101),
.B(n_114),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_SL g2607 ( 
.A(n_2011),
.B(n_115),
.Y(n_2607)
);

NAND2xp33_ASAP7_75t_SL g2608 ( 
.A(n_2101),
.B(n_114),
.Y(n_2608)
);

NAND2xp33_ASAP7_75t_SL g2609 ( 
.A(n_2101),
.B(n_114),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_SL g2610 ( 
.A(n_2011),
.B(n_117),
.Y(n_2610)
);

NAND2xp33_ASAP7_75t_SL g2611 ( 
.A(n_2101),
.B(n_116),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_SL g2612 ( 
.A(n_2011),
.B(n_117),
.Y(n_2612)
);

NAND2xp33_ASAP7_75t_SL g2613 ( 
.A(n_2101),
.B(n_116),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2001),
.B(n_117),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2033),
.B(n_119),
.Y(n_2615)
);

NAND2xp33_ASAP7_75t_SL g2616 ( 
.A(n_2101),
.B(n_119),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2011),
.B(n_121),
.Y(n_2617)
);

NAND2xp33_ASAP7_75t_SL g2618 ( 
.A(n_2101),
.B(n_120),
.Y(n_2618)
);

NAND2xp33_ASAP7_75t_SL g2619 ( 
.A(n_2101),
.B(n_120),
.Y(n_2619)
);

AND2x4_ASAP7_75t_L g2620 ( 
.A(n_2178),
.B(n_120),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2264),
.B(n_122),
.Y(n_2621)
);

NAND2xp33_ASAP7_75t_SL g2622 ( 
.A(n_2101),
.B(n_122),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_2011),
.B(n_125),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2011),
.B(n_125),
.Y(n_2624)
);

NAND2xp33_ASAP7_75t_SL g2625 ( 
.A(n_2101),
.B(n_123),
.Y(n_2625)
);

NAND2xp33_ASAP7_75t_SL g2626 ( 
.A(n_2101),
.B(n_123),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_SL g2627 ( 
.A(n_2011),
.B(n_126),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2011),
.B(n_127),
.Y(n_2628)
);

NAND2xp33_ASAP7_75t_SL g2629 ( 
.A(n_2101),
.B(n_123),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2011),
.B(n_129),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2011),
.B(n_129),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2011),
.B(n_130),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2011),
.B(n_130),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2011),
.B(n_131),
.Y(n_2634)
);

NAND2xp33_ASAP7_75t_SL g2635 ( 
.A(n_2101),
.B(n_128),
.Y(n_2635)
);

NAND2xp33_ASAP7_75t_SL g2636 ( 
.A(n_2101),
.B(n_128),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2011),
.B(n_132),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2011),
.B(n_133),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2011),
.B(n_134),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2264),
.B(n_131),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2011),
.B(n_135),
.Y(n_2641)
);

NAND2xp33_ASAP7_75t_SL g2642 ( 
.A(n_2101),
.B(n_131),
.Y(n_2642)
);

NAND2xp33_ASAP7_75t_SL g2643 ( 
.A(n_2101),
.B(n_135),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2011),
.B(n_136),
.Y(n_2644)
);

NAND3xp33_ASAP7_75t_L g2645 ( 
.A(n_2235),
.B(n_135),
.C(n_136),
.Y(n_2645)
);

NAND2xp33_ASAP7_75t_SL g2646 ( 
.A(n_2101),
.B(n_138),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2011),
.B(n_139),
.Y(n_2647)
);

NAND2xp33_ASAP7_75t_SL g2648 ( 
.A(n_2101),
.B(n_138),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_2011),
.B(n_139),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_SL g2650 ( 
.A(n_2011),
.B(n_140),
.Y(n_2650)
);

NAND2xp33_ASAP7_75t_SL g2651 ( 
.A(n_2101),
.B(n_138),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_L g2652 ( 
.A(n_2208),
.B(n_140),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_SL g2653 ( 
.A(n_2132),
.B(n_141),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2011),
.B(n_142),
.Y(n_2654)
);

NAND2xp33_ASAP7_75t_SL g2655 ( 
.A(n_2101),
.B(n_141),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2011),
.B(n_144),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2033),
.B(n_143),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2033),
.B(n_143),
.Y(n_2658)
);

NAND2xp33_ASAP7_75t_SL g2659 ( 
.A(n_2101),
.B(n_143),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2264),
.B(n_146),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2264),
.B(n_148),
.Y(n_2661)
);

AND2x2_ASAP7_75t_SL g2662 ( 
.A(n_2101),
.B(n_148),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2264),
.B(n_149),
.Y(n_2663)
);

NAND2xp33_ASAP7_75t_SL g2664 ( 
.A(n_2101),
.B(n_150),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2011),
.B(n_151),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_SL g2666 ( 
.A(n_2011),
.B(n_151),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2033),
.B(n_150),
.Y(n_2667)
);

NAND2xp33_ASAP7_75t_SL g2668 ( 
.A(n_2101),
.B(n_152),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2011),
.B(n_153),
.Y(n_2669)
);

NAND2xp33_ASAP7_75t_SL g2670 ( 
.A(n_2101),
.B(n_152),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2011),
.B(n_155),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2011),
.B(n_155),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2011),
.B(n_156),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2011),
.B(n_156),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2011),
.B(n_156),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_2011),
.B(n_157),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2011),
.B(n_157),
.Y(n_2677)
);

NAND2xp33_ASAP7_75t_SL g2678 ( 
.A(n_2101),
.B(n_154),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2033),
.B(n_154),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2011),
.B(n_158),
.Y(n_2680)
);

AND2x4_ASAP7_75t_L g2681 ( 
.A(n_2178),
.B(n_157),
.Y(n_2681)
);

NAND2xp33_ASAP7_75t_SL g2682 ( 
.A(n_2101),
.B(n_159),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2011),
.B(n_161),
.Y(n_2683)
);

NAND2xp33_ASAP7_75t_SL g2684 ( 
.A(n_2101),
.B(n_160),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2033),
.B(n_162),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2011),
.B(n_163),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2011),
.B(n_163),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2033),
.B(n_162),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2011),
.B(n_165),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2033),
.B(n_164),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2011),
.B(n_166),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2011),
.B(n_166),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_2011),
.B(n_166),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2011),
.B(n_167),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_L g2695 ( 
.A(n_2208),
.B(n_164),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2011),
.B(n_167),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2011),
.B(n_168),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2011),
.B(n_168),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_2011),
.B(n_168),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_SL g2700 ( 
.A(n_2011),
.B(n_169),
.Y(n_2700)
);

NAND2xp33_ASAP7_75t_SL g2701 ( 
.A(n_2101),
.B(n_164),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2011),
.B(n_171),
.Y(n_2702)
);

NAND2xp33_ASAP7_75t_SL g2703 ( 
.A(n_2101),
.B(n_170),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2033),
.B(n_170),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_2011),
.B(n_172),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2011),
.B(n_173),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2011),
.B(n_174),
.Y(n_2707)
);

NAND2xp33_ASAP7_75t_SL g2708 ( 
.A(n_2101),
.B(n_172),
.Y(n_2708)
);

NAND2xp33_ASAP7_75t_SL g2709 ( 
.A(n_2101),
.B(n_175),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2208),
.B(n_176),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2011),
.B(n_177),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2011),
.B(n_178),
.Y(n_2712)
);

NAND2xp33_ASAP7_75t_SL g2713 ( 
.A(n_2101),
.B(n_176),
.Y(n_2713)
);

NAND2xp33_ASAP7_75t_SL g2714 ( 
.A(n_2101),
.B(n_178),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2011),
.B(n_179),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2011),
.B(n_179),
.Y(n_2716)
);

NAND2xp33_ASAP7_75t_SL g2717 ( 
.A(n_2101),
.B(n_178),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2264),
.B(n_179),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2011),
.B(n_182),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2264),
.B(n_180),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2264),
.B(n_183),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2011),
.B(n_185),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2264),
.B(n_183),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2387),
.B(n_186),
.Y(n_2724)
);

OAI21x1_ASAP7_75t_L g2725 ( 
.A1(n_2536),
.A2(n_186),
.B(n_187),
.Y(n_2725)
);

A2O1A1Ixp33_ASAP7_75t_L g2726 ( 
.A1(n_2326),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2529),
.Y(n_2727)
);

OR2x2_ASAP7_75t_L g2728 ( 
.A(n_2614),
.B(n_187),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2284),
.B(n_2299),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2306),
.B(n_540),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2339),
.B(n_188),
.Y(n_2731)
);

AOI21xp5_ASAP7_75t_SL g2732 ( 
.A1(n_2529),
.A2(n_189),
.B(n_190),
.Y(n_2732)
);

CKINVDCx8_ASAP7_75t_R g2733 ( 
.A(n_2544),
.Y(n_2733)
);

O2A1O1Ixp33_ASAP7_75t_SL g2734 ( 
.A1(n_2504),
.A2(n_2510),
.B(n_2562),
.C(n_2561),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2405),
.Y(n_2735)
);

INVx4_ASAP7_75t_L g2736 ( 
.A(n_2529),
.Y(n_2736)
);

AO31x2_ASAP7_75t_L g2737 ( 
.A1(n_2489),
.A2(n_192),
.A3(n_190),
.B(n_191),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2329),
.A2(n_191),
.B(n_192),
.Y(n_2738)
);

OA21x2_ASAP7_75t_L g2739 ( 
.A1(n_2530),
.A2(n_191),
.B(n_192),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2329),
.A2(n_193),
.B(n_194),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2411),
.B(n_193),
.Y(n_2741)
);

NAND3xp33_ASAP7_75t_SL g2742 ( 
.A(n_2566),
.B(n_193),
.C(n_194),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_2306),
.B(n_541),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2405),
.Y(n_2744)
);

O2A1O1Ixp33_ASAP7_75t_SL g2745 ( 
.A1(n_2532),
.A2(n_2565),
.B(n_2564),
.C(n_2413),
.Y(n_2745)
);

A2O1A1Ixp33_ASAP7_75t_L g2746 ( 
.A1(n_2390),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2372),
.B(n_195),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2621),
.B(n_197),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2640),
.B(n_2660),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2661),
.B(n_197),
.Y(n_2750)
);

NAND2xp33_ASAP7_75t_R g2751 ( 
.A(n_2544),
.B(n_197),
.Y(n_2751)
);

OAI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2653),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2405),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2351),
.Y(n_2754)
);

AO31x2_ASAP7_75t_L g2755 ( 
.A1(n_2491),
.A2(n_2555),
.A3(n_2499),
.B(n_2569),
.Y(n_2755)
);

BUFx12f_ASAP7_75t_L g2756 ( 
.A(n_2544),
.Y(n_2756)
);

OAI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2332),
.A2(n_198),
.B(n_199),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2663),
.B(n_199),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2382),
.B(n_200),
.Y(n_2759)
);

OAI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2284),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2760)
);

AO31x2_ASAP7_75t_L g2761 ( 
.A1(n_2652),
.A2(n_203),
.A3(n_201),
.B(n_202),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2718),
.B(n_201),
.Y(n_2762)
);

A2O1A1Ixp33_ASAP7_75t_L g2763 ( 
.A1(n_2392),
.A2(n_2394),
.B(n_2397),
.C(n_2395),
.Y(n_2763)
);

CKINVDCx20_ASAP7_75t_R g2764 ( 
.A(n_2341),
.Y(n_2764)
);

AO31x2_ASAP7_75t_L g2765 ( 
.A1(n_2695),
.A2(n_206),
.A3(n_204),
.B(n_205),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2395),
.A2(n_205),
.B(n_207),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2397),
.A2(n_208),
.B(n_209),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2284),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2720),
.B(n_210),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_SL g2770 ( 
.A1(n_2501),
.A2(n_211),
.B(n_212),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2721),
.B(n_211),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2330),
.Y(n_2772)
);

NOR2xp67_ASAP7_75t_L g2773 ( 
.A(n_2302),
.B(n_212),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2342),
.B(n_212),
.Y(n_2774)
);

O2A1O1Ixp33_ASAP7_75t_SL g2775 ( 
.A1(n_2494),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_2775)
);

OAI22x1_ASAP7_75t_L g2776 ( 
.A1(n_2527),
.A2(n_216),
.B1(n_213),
.B2(n_215),
.Y(n_2776)
);

NOR2xp67_ASAP7_75t_L g2777 ( 
.A(n_2380),
.B(n_215),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2437),
.B(n_216),
.Y(n_2778)
);

OAI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2568),
.A2(n_216),
.B(n_217),
.Y(n_2779)
);

OAI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2583),
.A2(n_217),
.B(n_218),
.Y(n_2780)
);

OAI21xp33_ASAP7_75t_L g2781 ( 
.A1(n_2353),
.A2(n_218),
.B(n_219),
.Y(n_2781)
);

AO31x2_ASAP7_75t_L g2782 ( 
.A1(n_2710),
.A2(n_221),
.A3(n_219),
.B(n_220),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2723),
.B(n_219),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2398),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_2784)
);

AOI21xp5_ASAP7_75t_SL g2785 ( 
.A1(n_2299),
.A2(n_221),
.B(n_222),
.Y(n_2785)
);

NAND2x1p5_ASAP7_75t_L g2786 ( 
.A(n_2662),
.B(n_223),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2442),
.B(n_224),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_2299),
.Y(n_2788)
);

NAND3x1_ASAP7_75t_L g2789 ( 
.A(n_2550),
.B(n_224),
.C(n_226),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2344),
.B(n_226),
.Y(n_2790)
);

BUFx3_ASAP7_75t_L g2791 ( 
.A(n_2602),
.Y(n_2791)
);

BUFx2_ASAP7_75t_L g2792 ( 
.A(n_2602),
.Y(n_2792)
);

AND2x4_ASAP7_75t_L g2793 ( 
.A(n_2602),
.B(n_226),
.Y(n_2793)
);

NAND2xp33_ASAP7_75t_SL g2794 ( 
.A(n_2620),
.B(n_227),
.Y(n_2794)
);

AND2x2_ASAP7_75t_SL g2795 ( 
.A(n_2662),
.B(n_227),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2423),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2398),
.A2(n_227),
.B(n_228),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2585),
.B(n_228),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2587),
.B(n_228),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2592),
.B(n_229),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2595),
.B(n_229),
.Y(n_2801)
);

A2O1A1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2563),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_2802)
);

OAI21x1_ASAP7_75t_SL g2803 ( 
.A1(n_2506),
.A2(n_230),
.B(n_231),
.Y(n_2803)
);

NAND2x1p5_ASAP7_75t_L g2804 ( 
.A(n_2423),
.B(n_231),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_SL g2805 ( 
.A1(n_2620),
.A2(n_232),
.B(n_233),
.Y(n_2805)
);

NAND3x1_ASAP7_75t_L g2806 ( 
.A(n_2455),
.B(n_232),
.C(n_233),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2601),
.B(n_233),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2423),
.Y(n_2808)
);

OAI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2615),
.A2(n_234),
.B(n_235),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2620),
.Y(n_2810)
);

INVx8_ASAP7_75t_L g2811 ( 
.A(n_2681),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_SL g2812 ( 
.A(n_2276),
.B(n_543),
.Y(n_2812)
);

BUFx2_ASAP7_75t_L g2813 ( 
.A(n_2681),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2681),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2537),
.A2(n_2548),
.B1(n_2549),
.B2(n_2543),
.Y(n_2815)
);

AND2x4_ASAP7_75t_L g2816 ( 
.A(n_2381),
.B(n_236),
.Y(n_2816)
);

A2O1A1Ixp33_ASAP7_75t_L g2817 ( 
.A1(n_2563),
.A2(n_2309),
.B(n_2497),
.C(n_2495),
.Y(n_2817)
);

AOI31xp67_ASAP7_75t_L g2818 ( 
.A1(n_2520),
.A2(n_238),
.A3(n_236),
.B(n_237),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_SL g2819 ( 
.A1(n_2399),
.A2(n_236),
.B(n_237),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2657),
.B(n_237),
.Y(n_2820)
);

AO22x2_ASAP7_75t_L g2821 ( 
.A1(n_2539),
.A2(n_2541),
.B1(n_2542),
.B2(n_2540),
.Y(n_2821)
);

A2O1A1Ixp33_ASAP7_75t_L g2822 ( 
.A1(n_2309),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2822)
);

INVxp67_ASAP7_75t_L g2823 ( 
.A(n_2295),
.Y(n_2823)
);

BUFx6f_ASAP7_75t_L g2824 ( 
.A(n_2399),
.Y(n_2824)
);

A2O1A1Ixp33_ASAP7_75t_L g2825 ( 
.A1(n_2525),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_2825)
);

NAND2x1p5_ASAP7_75t_L g2826 ( 
.A(n_2404),
.B(n_240),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_2399),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2381),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2828)
);

CKINVDCx20_ASAP7_75t_R g2829 ( 
.A(n_2465),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2658),
.B(n_2667),
.Y(n_2830)
);

AOI21x1_ASAP7_75t_L g2831 ( 
.A1(n_2393),
.A2(n_2507),
.B(n_2391),
.Y(n_2831)
);

AO32x2_ASAP7_75t_L g2832 ( 
.A1(n_2554),
.A2(n_245),
.A3(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_2832)
);

BUFx2_ASAP7_75t_L g2833 ( 
.A(n_2381),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2679),
.B(n_245),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2685),
.B(n_247),
.Y(n_2835)
);

O2A1O1Ixp33_ASAP7_75t_L g2836 ( 
.A1(n_2389),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2688),
.B(n_249),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2377),
.A2(n_250),
.B(n_251),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2378),
.A2(n_251),
.B(n_252),
.Y(n_2839)
);

CKINVDCx8_ASAP7_75t_R g2840 ( 
.A(n_2471),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2479),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2484),
.B(n_252),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_2276),
.B(n_546),
.Y(n_2843)
);

AOI211x1_ASAP7_75t_L g2844 ( 
.A1(n_2547),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2285),
.B(n_547),
.Y(n_2845)
);

AO22x1_ASAP7_75t_L g2846 ( 
.A1(n_2531),
.A2(n_2535),
.B1(n_2453),
.B2(n_2444),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2480),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2690),
.B(n_253),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2439),
.A2(n_253),
.B(n_254),
.Y(n_2849)
);

OAI22xp5_ASAP7_75t_L g2850 ( 
.A1(n_2704),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_2850)
);

AND2x4_ASAP7_75t_L g2851 ( 
.A(n_2348),
.B(n_255),
.Y(n_2851)
);

AO21x1_ASAP7_75t_L g2852 ( 
.A1(n_2514),
.A2(n_2515),
.B(n_2534),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2324),
.B(n_257),
.Y(n_2853)
);

NAND3x1_ASAP7_75t_L g2854 ( 
.A(n_2486),
.B(n_257),
.C(n_258),
.Y(n_2854)
);

INVx1_ASAP7_75t_SL g2855 ( 
.A(n_2400),
.Y(n_2855)
);

BUFx12f_ASAP7_75t_L g2856 ( 
.A(n_2477),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2558),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_2338),
.Y(n_2858)
);

OAI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2420),
.A2(n_262),
.B(n_263),
.Y(n_2859)
);

AND2x6_ASAP7_75t_L g2860 ( 
.A(n_2477),
.B(n_263),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2516),
.B(n_264),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2285),
.B(n_548),
.Y(n_2862)
);

OAI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_2533),
.A2(n_2557),
.B(n_2318),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2509),
.Y(n_2864)
);

OAI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2477),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2513),
.Y(n_2866)
);

A2O1A1Ixp33_ASAP7_75t_L g2867 ( 
.A1(n_2452),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2422),
.A2(n_267),
.B(n_268),
.Y(n_2868)
);

OAI22x1_ASAP7_75t_L g2869 ( 
.A1(n_2508),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_2869)
);

NAND3xp33_ASAP7_75t_L g2870 ( 
.A(n_2556),
.B(n_270),
.C(n_271),
.Y(n_2870)
);

OAI22x1_ASAP7_75t_L g2871 ( 
.A1(n_2512),
.A2(n_273),
.B1(n_270),
.B2(n_272),
.Y(n_2871)
);

OAI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2538),
.A2(n_272),
.B(n_273),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2283),
.B(n_272),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2280),
.B(n_274),
.Y(n_2874)
);

NOR2x1_ASAP7_75t_L g2875 ( 
.A(n_2340),
.B(n_275),
.Y(n_2875)
);

OAI22xp5_ASAP7_75t_L g2876 ( 
.A1(n_2431),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2606),
.B(n_2608),
.Y(n_2877)
);

OAI21x1_ASAP7_75t_L g2878 ( 
.A1(n_2370),
.A2(n_2371),
.B(n_2383),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2296),
.B(n_277),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2346),
.B(n_278),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2286),
.B(n_278),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2347),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2291),
.B(n_279),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2293),
.B(n_279),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2312),
.B(n_280),
.Y(n_2885)
);

OAI22x1_ASAP7_75t_L g2886 ( 
.A1(n_2552),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_2886)
);

AOI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2388),
.A2(n_2384),
.B(n_2429),
.Y(n_2887)
);

BUFx3_ASAP7_75t_L g2888 ( 
.A(n_2368),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2334),
.Y(n_2889)
);

BUFx10_ASAP7_75t_L g2890 ( 
.A(n_2354),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2313),
.B(n_285),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2435),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2425),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2468),
.B(n_285),
.Y(n_2894)
);

OAI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2645),
.A2(n_2519),
.B(n_2559),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2408),
.B(n_286),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_SL g2897 ( 
.A(n_2606),
.B(n_550),
.Y(n_2897)
);

OAI21x1_ASAP7_75t_L g2898 ( 
.A1(n_2457),
.A2(n_286),
.B(n_287),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2359),
.B(n_287),
.Y(n_2899)
);

AOI211x1_ASAP7_75t_L g2900 ( 
.A1(n_2526),
.A2(n_2528),
.B(n_2493),
.C(n_2443),
.Y(n_2900)
);

CKINVDCx20_ASAP7_75t_R g2901 ( 
.A(n_2335),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2314),
.B(n_288),
.Y(n_2902)
);

AO31x2_ASAP7_75t_L g2903 ( 
.A1(n_2502),
.A2(n_292),
.A3(n_290),
.B(n_291),
.Y(n_2903)
);

OR2x6_ASAP7_75t_L g2904 ( 
.A(n_2521),
.B(n_291),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2461),
.B(n_293),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2560),
.B(n_293),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2333),
.B(n_295),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_SL g2908 ( 
.A1(n_2570),
.A2(n_295),
.B(n_296),
.Y(n_2908)
);

AND2x4_ASAP7_75t_L g2909 ( 
.A(n_2325),
.B(n_2316),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2427),
.Y(n_2910)
);

AOI211x1_ASAP7_75t_L g2911 ( 
.A1(n_2441),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2545),
.B(n_298),
.Y(n_2912)
);

NAND3xp33_ASAP7_75t_L g2913 ( 
.A(n_2503),
.B(n_299),
.C(n_300),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2373),
.A2(n_299),
.B(n_300),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2374),
.A2(n_2375),
.B(n_2385),
.Y(n_2915)
);

AOI211x1_ASAP7_75t_L g2916 ( 
.A1(n_2396),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_2511),
.Y(n_2917)
);

O2A1O1Ixp5_ASAP7_75t_L g2918 ( 
.A1(n_2402),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2608),
.B(n_551),
.Y(n_2919)
);

CKINVDCx5p33_ASAP7_75t_R g2920 ( 
.A(n_2459),
.Y(n_2920)
);

OAI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2415),
.A2(n_303),
.B(n_304),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2352),
.B(n_303),
.Y(n_2922)
);

INVxp67_ASAP7_75t_L g2923 ( 
.A(n_2522),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2428),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2403),
.B(n_304),
.Y(n_2925)
);

OAI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2430),
.A2(n_305),
.B(n_306),
.Y(n_2926)
);

HB1xp67_ASAP7_75t_L g2927 ( 
.A(n_2523),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2546),
.B(n_305),
.Y(n_2928)
);

AOI221x1_ASAP7_75t_L g2929 ( 
.A1(n_2505),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.C(n_308),
.Y(n_2929)
);

AO31x2_ASAP7_75t_L g2930 ( 
.A1(n_2551),
.A2(n_309),
.A3(n_307),
.B(n_308),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2290),
.B(n_308),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2553),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2482),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2292),
.B(n_309),
.Y(n_2934)
);

AO31x2_ASAP7_75t_L g2935 ( 
.A1(n_2409),
.A2(n_2414),
.A3(n_2419),
.B(n_2410),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2294),
.B(n_310),
.Y(n_2936)
);

OAI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2450),
.A2(n_310),
.B(n_311),
.Y(n_2937)
);

OAI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_2571),
.A2(n_314),
.B1(n_311),
.B2(n_313),
.Y(n_2938)
);

A2O1A1Ixp33_ASAP7_75t_L g2939 ( 
.A1(n_2454),
.A2(n_315),
.B(n_311),
.C(n_314),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2436),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2940)
);

CKINVDCx5p33_ASAP7_75t_R g2941 ( 
.A(n_2343),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2448),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2297),
.B(n_316),
.Y(n_2943)
);

BUFx2_ASAP7_75t_L g2944 ( 
.A(n_2609),
.Y(n_2944)
);

AOI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2476),
.A2(n_316),
.B(n_317),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2418),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2433),
.Y(n_2947)
);

CKINVDCx5p33_ASAP7_75t_R g2948 ( 
.A(n_2345),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2524),
.B(n_317),
.Y(n_2949)
);

OAI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2434),
.A2(n_318),
.B(n_319),
.Y(n_2950)
);

NAND3x1_ASAP7_75t_L g2951 ( 
.A(n_2609),
.B(n_318),
.C(n_319),
.Y(n_2951)
);

BUFx2_ASAP7_75t_L g2952 ( 
.A(n_2611),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2298),
.B(n_2300),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2301),
.B(n_320),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_L g2955 ( 
.A(n_2462),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2337),
.B(n_320),
.Y(n_2956)
);

AO31x2_ASAP7_75t_L g2957 ( 
.A1(n_2409),
.A2(n_323),
.A3(n_321),
.B(n_322),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2277),
.Y(n_2958)
);

BUFx4f_ASAP7_75t_L g2959 ( 
.A(n_2458),
.Y(n_2959)
);

OAI21x1_ASAP7_75t_L g2960 ( 
.A1(n_2451),
.A2(n_321),
.B(n_322),
.Y(n_2960)
);

BUFx2_ASAP7_75t_L g2961 ( 
.A(n_2611),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_SL g2962 ( 
.A1(n_2573),
.A2(n_324),
.B(n_325),
.Y(n_2962)
);

OR2x2_ASAP7_75t_L g2963 ( 
.A(n_2311),
.B(n_327),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2440),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2307),
.B(n_2323),
.Y(n_2965)
);

AOI21x1_ASAP7_75t_SL g2966 ( 
.A1(n_2282),
.A2(n_328),
.B(n_329),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2319),
.B(n_330),
.Y(n_2967)
);

CKINVDCx5p33_ASAP7_75t_R g2968 ( 
.A(n_2349),
.Y(n_2968)
);

NOR2xp67_ASAP7_75t_L g2969 ( 
.A(n_2406),
.B(n_331),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2288),
.B(n_331),
.Y(n_2970)
);

OAI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2496),
.A2(n_332),
.B(n_333),
.Y(n_2971)
);

INVx4_ASAP7_75t_L g2972 ( 
.A(n_2613),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2289),
.B(n_332),
.Y(n_2973)
);

AOI21x1_ASAP7_75t_SL g2974 ( 
.A1(n_2282),
.A2(n_332),
.B(n_333),
.Y(n_2974)
);

AOI211x1_ASAP7_75t_L g2975 ( 
.A1(n_2518),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2417),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2367),
.B(n_334),
.Y(n_2977)
);

OAI21x1_ASAP7_75t_L g2978 ( 
.A1(n_2498),
.A2(n_335),
.B(n_336),
.Y(n_2978)
);

INVx5_ASAP7_75t_L g2979 ( 
.A(n_2613),
.Y(n_2979)
);

OAI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2464),
.A2(n_336),
.B(n_337),
.Y(n_2980)
);

BUFx3_ASAP7_75t_L g2981 ( 
.A(n_2277),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2321),
.B(n_337),
.Y(n_2982)
);

BUFx10_ASAP7_75t_L g2983 ( 
.A(n_2362),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_2616),
.Y(n_2984)
);

AOI21xp33_ASAP7_75t_L g2985 ( 
.A1(n_2369),
.A2(n_339),
.B(n_340),
.Y(n_2985)
);

OAI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2574),
.A2(n_339),
.B(n_341),
.Y(n_2986)
);

OAI21x1_ASAP7_75t_SL g2987 ( 
.A1(n_2616),
.A2(n_341),
.B(n_342),
.Y(n_2987)
);

OAI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2575),
.A2(n_341),
.B(n_342),
.Y(n_2988)
);

BUFx6f_ASAP7_75t_L g2989 ( 
.A(n_2467),
.Y(n_2989)
);

BUFx2_ASAP7_75t_L g2990 ( 
.A(n_2618),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2322),
.B(n_342),
.Y(n_2991)
);

O2A1O1Ixp5_ASAP7_75t_L g2992 ( 
.A1(n_2412),
.A2(n_2303),
.B(n_2577),
.C(n_2576),
.Y(n_2992)
);

BUFx3_ASAP7_75t_L g2993 ( 
.A(n_2331),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2315),
.B(n_2317),
.Y(n_2994)
);

AO31x2_ASAP7_75t_L g2995 ( 
.A1(n_2410),
.A2(n_345),
.A3(n_343),
.B(n_344),
.Y(n_2995)
);

NOR2x1_ASAP7_75t_SL g2996 ( 
.A(n_2456),
.B(n_2446),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2308),
.B(n_343),
.Y(n_2997)
);

OR2x2_ASAP7_75t_L g2998 ( 
.A(n_2320),
.B(n_343),
.Y(n_2998)
);

OAI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2578),
.A2(n_345),
.B(n_346),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_L g3000 ( 
.A1(n_2472),
.A2(n_346),
.B(n_347),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2438),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2463),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2481),
.A2(n_348),
.B(n_349),
.Y(n_3003)
);

AO21x1_ASAP7_75t_L g3004 ( 
.A1(n_2618),
.A2(n_552),
.B(n_551),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2619),
.B(n_552),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2447),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2364),
.B(n_348),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2365),
.B(n_349),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2287),
.Y(n_3009)
);

OAI21xp33_ASAP7_75t_L g3010 ( 
.A1(n_2579),
.A2(n_349),
.B(n_350),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2580),
.A2(n_2716),
.B(n_2715),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2366),
.B(n_350),
.Y(n_3012)
);

O2A1O1Ixp33_ASAP7_75t_SL g3013 ( 
.A1(n_2581),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2492),
.Y(n_3014)
);

AO31x2_ASAP7_75t_L g3015 ( 
.A1(n_2414),
.A2(n_2419),
.A3(n_2426),
.B(n_2424),
.Y(n_3015)
);

AOI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2416),
.A2(n_351),
.B(n_352),
.Y(n_3016)
);

O2A1O1Ixp5_ASAP7_75t_L g3017 ( 
.A1(n_2582),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2470),
.B(n_353),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2488),
.A2(n_354),
.B(n_355),
.Y(n_3019)
);

OAI21x1_ASAP7_75t_L g3020 ( 
.A1(n_2474),
.A2(n_355),
.B(n_356),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2421),
.B(n_357),
.Y(n_3021)
);

AO31x2_ASAP7_75t_L g3022 ( 
.A1(n_2424),
.A2(n_360),
.A3(n_357),
.B(n_359),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2327),
.B(n_357),
.Y(n_3023)
);

AOI221xp5_ASAP7_75t_L g3024 ( 
.A1(n_2407),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.C(n_362),
.Y(n_3024)
);

OR2x2_ASAP7_75t_L g3025 ( 
.A(n_2281),
.B(n_360),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_L g3026 ( 
.A(n_2469),
.Y(n_3026)
);

AOI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2586),
.A2(n_362),
.B(n_363),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2478),
.Y(n_3028)
);

OAI21x1_ASAP7_75t_L g3029 ( 
.A1(n_2589),
.A2(n_363),
.B(n_364),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2304),
.B(n_364),
.Y(n_3030)
);

NAND3xp33_ASAP7_75t_L g3031 ( 
.A(n_2473),
.B(n_2500),
.C(n_2445),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2590),
.A2(n_2591),
.B1(n_2597),
.B2(n_2593),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2598),
.A2(n_365),
.B(n_366),
.Y(n_3033)
);

OAI21x1_ASAP7_75t_L g3034 ( 
.A1(n_2722),
.A2(n_365),
.B(n_366),
.Y(n_3034)
);

INVx2_ASAP7_75t_SL g3035 ( 
.A(n_2466),
.Y(n_3035)
);

OR2x2_ASAP7_75t_L g3036 ( 
.A(n_2357),
.B(n_367),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2619),
.B(n_553),
.Y(n_3037)
);

OR2x6_ASAP7_75t_L g3038 ( 
.A(n_2279),
.B(n_367),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_SL g3039 ( 
.A(n_2460),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2278),
.B(n_368),
.Y(n_3040)
);

AO31x2_ASAP7_75t_L g3041 ( 
.A1(n_2426),
.A2(n_371),
.A3(n_369),
.B(n_370),
.Y(n_3041)
);

INVxp67_ASAP7_75t_SL g3042 ( 
.A(n_2600),
.Y(n_3042)
);

AOI221x1_ASAP7_75t_L g3043 ( 
.A1(n_2622),
.A2(n_2626),
.B1(n_2635),
.B2(n_2629),
.C(n_2625),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2355),
.B(n_371),
.Y(n_3044)
);

AOI221x1_ASAP7_75t_L g3045 ( 
.A1(n_2622),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.C(n_376),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2490),
.Y(n_3046)
);

OAI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2603),
.A2(n_373),
.B(n_374),
.Y(n_3047)
);

OAI21x1_ASAP7_75t_L g3048 ( 
.A1(n_2604),
.A2(n_375),
.B(n_376),
.Y(n_3048)
);

AOI221x1_ASAP7_75t_L g3049 ( 
.A1(n_2625),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.C(n_381),
.Y(n_3049)
);

INVxp67_ASAP7_75t_SL g3050 ( 
.A(n_2607),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2610),
.A2(n_381),
.B(n_382),
.Y(n_3051)
);

OAI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2612),
.A2(n_382),
.B(n_383),
.Y(n_3052)
);

BUFx6f_ASAP7_75t_L g3053 ( 
.A(n_2376),
.Y(n_3053)
);

AO31x2_ASAP7_75t_L g3054 ( 
.A1(n_2432),
.A2(n_384),
.A3(n_382),
.B(n_383),
.Y(n_3054)
);

AO21x1_ASAP7_75t_L g3055 ( 
.A1(n_2626),
.A2(n_554),
.B(n_553),
.Y(n_3055)
);

OR2x6_ASAP7_75t_L g3056 ( 
.A(n_2358),
.B(n_385),
.Y(n_3056)
);

INVx2_ASAP7_75t_SL g3057 ( 
.A(n_2350),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_R g3058 ( 
.A(n_2629),
.B(n_385),
.Y(n_3058)
);

AOI221x1_ASAP7_75t_L g3059 ( 
.A1(n_2635),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.C(n_389),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2328),
.B(n_386),
.Y(n_3060)
);

OAI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2617),
.A2(n_386),
.B(n_387),
.Y(n_3061)
);

AOI221xp5_ASAP7_75t_L g3062 ( 
.A1(n_2363),
.A2(n_390),
.B1(n_387),
.B2(n_388),
.C(n_391),
.Y(n_3062)
);

CKINVDCx5p33_ASAP7_75t_R g3063 ( 
.A(n_2336),
.Y(n_3063)
);

AO31x2_ASAP7_75t_L g3064 ( 
.A1(n_2432),
.A2(n_391),
.A3(n_388),
.B(n_390),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2356),
.B(n_2305),
.Y(n_3065)
);

NAND2x1p5_ASAP7_75t_L g3066 ( 
.A(n_2360),
.B(n_2401),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2623),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2275),
.B(n_2517),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2624),
.B(n_392),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2475),
.Y(n_3070)
);

A2O1A1Ixp33_ASAP7_75t_L g3071 ( 
.A1(n_2636),
.A2(n_395),
.B(n_393),
.C(n_394),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2627),
.B(n_395),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2628),
.B(n_397),
.Y(n_3073)
);

NOR2x1_ASAP7_75t_L g3074 ( 
.A(n_2310),
.B(n_398),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2630),
.B(n_398),
.Y(n_3075)
);

OAI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2631),
.A2(n_399),
.B(n_400),
.Y(n_3076)
);

AOI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_2636),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_3077)
);

BUFx3_ASAP7_75t_L g3078 ( 
.A(n_2379),
.Y(n_3078)
);

NOR2x1_ASAP7_75t_R g3079 ( 
.A(n_2386),
.B(n_400),
.Y(n_3079)
);

OAI21xp33_ASAP7_75t_L g3080 ( 
.A1(n_2632),
.A2(n_401),
.B(n_402),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_2633),
.A2(n_401),
.B(n_402),
.Y(n_3081)
);

OAI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2634),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2637),
.A2(n_403),
.B(n_405),
.Y(n_3083)
);

OAI22x1_ASAP7_75t_L g3084 ( 
.A1(n_2638),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2639),
.A2(n_406),
.B(n_407),
.Y(n_3085)
);

BUFx2_ASAP7_75t_L g3086 ( 
.A(n_2642),
.Y(n_3086)
);

AO22x2_ASAP7_75t_L g3087 ( 
.A1(n_2641),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2644),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2647),
.B(n_410),
.Y(n_3089)
);

A2O1A1Ixp33_ASAP7_75t_L g3090 ( 
.A1(n_2642),
.A2(n_414),
.B(n_411),
.C(n_413),
.Y(n_3090)
);

OR2x6_ASAP7_75t_L g3091 ( 
.A(n_2449),
.B(n_413),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2649),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2650),
.Y(n_3093)
);

BUFx4_ASAP7_75t_SL g3094 ( 
.A(n_2643),
.Y(n_3094)
);

NAND2x1p5_ASAP7_75t_L g3095 ( 
.A(n_2654),
.B(n_413),
.Y(n_3095)
);

AOI221xp5_ASAP7_75t_L g3096 ( 
.A1(n_2361),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_3096)
);

NAND3x1_ASAP7_75t_L g3097 ( 
.A(n_2643),
.B(n_414),
.C(n_415),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2656),
.A2(n_416),
.B(n_417),
.Y(n_3098)
);

AOI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2646),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_3099)
);

OAI21x1_ASAP7_75t_SL g3100 ( 
.A1(n_2646),
.A2(n_419),
.B(n_420),
.Y(n_3100)
);

O2A1O1Ixp5_ASAP7_75t_L g3101 ( 
.A1(n_2665),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2666),
.Y(n_3102)
);

OAI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2669),
.A2(n_422),
.B(n_423),
.Y(n_3103)
);

BUFx3_ASAP7_75t_L g3104 ( 
.A(n_2648),
.Y(n_3104)
);

OAI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2671),
.A2(n_422),
.B(n_423),
.Y(n_3105)
);

AO31x2_ASAP7_75t_L g3106 ( 
.A1(n_2648),
.A2(n_2655),
.A3(n_2659),
.B(n_2651),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2672),
.A2(n_422),
.B(n_423),
.Y(n_3107)
);

AO31x2_ASAP7_75t_L g3108 ( 
.A1(n_2651),
.A2(n_426),
.A3(n_424),
.B(n_425),
.Y(n_3108)
);

INVx3_ASAP7_75t_L g3109 ( 
.A(n_2655),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2673),
.A2(n_424),
.B(n_425),
.Y(n_3110)
);

AOI211x1_ASAP7_75t_L g3111 ( 
.A1(n_2674),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_3111)
);

O2A1O1Ixp5_ASAP7_75t_L g3112 ( 
.A1(n_2675),
.A2(n_2677),
.B(n_2680),
.C(n_2676),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2659),
.B(n_555),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2683),
.Y(n_3114)
);

A2O1A1Ixp33_ASAP7_75t_L g3115 ( 
.A1(n_2664),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_3115)
);

BUFx3_ASAP7_75t_L g3116 ( 
.A(n_2664),
.Y(n_3116)
);

AND2x4_ASAP7_75t_L g3117 ( 
.A(n_2686),
.B(n_432),
.Y(n_3117)
);

BUFx10_ASAP7_75t_L g3118 ( 
.A(n_2668),
.Y(n_3118)
);

CKINVDCx16_ASAP7_75t_R g3119 ( 
.A(n_2668),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_SL g3120 ( 
.A1(n_2687),
.A2(n_432),
.B(n_433),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2689),
.B(n_433),
.Y(n_3121)
);

BUFx3_ASAP7_75t_L g3122 ( 
.A(n_2670),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2691),
.B(n_434),
.Y(n_3123)
);

INVxp67_ASAP7_75t_SL g3124 ( 
.A(n_2692),
.Y(n_3124)
);

O2A1O1Ixp33_ASAP7_75t_SL g3125 ( 
.A1(n_2693),
.A2(n_436),
.B(n_434),
.C(n_435),
.Y(n_3125)
);

BUFx2_ASAP7_75t_L g3126 ( 
.A(n_2670),
.Y(n_3126)
);

NOR2x1_ASAP7_75t_R g3127 ( 
.A(n_2694),
.B(n_435),
.Y(n_3127)
);

HB1xp67_ASAP7_75t_L g3128 ( 
.A(n_2696),
.Y(n_3128)
);

O2A1O1Ixp5_ASAP7_75t_L g3129 ( 
.A1(n_2697),
.A2(n_2699),
.B(n_2700),
.C(n_2698),
.Y(n_3129)
);

OAI21x1_ASAP7_75t_SL g3130 ( 
.A1(n_2972),
.A2(n_2682),
.B(n_2678),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2737),
.Y(n_3131)
);

INVxp67_ASAP7_75t_SL g3132 ( 
.A(n_2729),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2737),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2737),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_SL g3135 ( 
.A(n_2733),
.B(n_2678),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2795),
.A2(n_2714),
.B1(n_2717),
.B2(n_2713),
.Y(n_3136)
);

AOI221xp5_ASAP7_75t_L g3137 ( 
.A1(n_2861),
.A2(n_2701),
.B1(n_2703),
.B2(n_2684),
.C(n_2682),
.Y(n_3137)
);

AO221x2_ASAP7_75t_L g3138 ( 
.A1(n_2846),
.A2(n_2703),
.B1(n_2708),
.B2(n_2701),
.C(n_2684),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_SL g3139 ( 
.A(n_2840),
.B(n_2708),
.Y(n_3139)
);

AO21x2_ASAP7_75t_L g3140 ( 
.A1(n_2763),
.A2(n_2705),
.B(n_2702),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2772),
.Y(n_3141)
);

AOI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2877),
.A2(n_2707),
.B(n_2706),
.Y(n_3142)
);

OAI21x1_ASAP7_75t_SL g3143 ( 
.A1(n_2972),
.A2(n_2713),
.B(n_2709),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_SL g3144 ( 
.A(n_2764),
.B(n_2709),
.Y(n_3144)
);

AOI22xp33_ASAP7_75t_L g3145 ( 
.A1(n_2756),
.A2(n_2717),
.B1(n_2714),
.B2(n_2572),
.Y(n_3145)
);

OA21x2_ASAP7_75t_L g3146 ( 
.A1(n_2817),
.A2(n_2712),
.B(n_2711),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2727),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2957),
.Y(n_3148)
);

BUFx2_ASAP7_75t_L g3149 ( 
.A(n_2856),
.Y(n_3149)
);

AO21x2_ASAP7_75t_L g3150 ( 
.A1(n_3031),
.A2(n_2719),
.B(n_2485),
.Y(n_3150)
);

BUFx6f_ASAP7_75t_L g3151 ( 
.A(n_2811),
.Y(n_3151)
);

CKINVDCx16_ASAP7_75t_R g3152 ( 
.A(n_2751),
.Y(n_3152)
);

AO21x1_ASAP7_75t_L g3153 ( 
.A1(n_2794),
.A2(n_2786),
.B(n_2743),
.Y(n_3153)
);

OA21x2_ASAP7_75t_L g3154 ( 
.A1(n_3043),
.A2(n_2487),
.B(n_2483),
.Y(n_3154)
);

OAI21x1_ASAP7_75t_L g3155 ( 
.A1(n_2958),
.A2(n_2584),
.B(n_2567),
.Y(n_3155)
);

OAI21x1_ASAP7_75t_L g3156 ( 
.A1(n_2966),
.A2(n_2974),
.B(n_2831),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2957),
.Y(n_3157)
);

AOI221xp5_ASAP7_75t_L g3158 ( 
.A1(n_2759),
.A2(n_2596),
.B1(n_2599),
.B2(n_2594),
.C(n_2588),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2957),
.Y(n_3159)
);

OAI21x1_ASAP7_75t_L g3160 ( 
.A1(n_2878),
.A2(n_2605),
.B(n_438),
.Y(n_3160)
);

OAI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_3119),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2932),
.B(n_436),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2995),
.Y(n_3163)
);

AOI21x1_ASAP7_75t_L g3164 ( 
.A1(n_2944),
.A2(n_557),
.B(n_556),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2995),
.Y(n_3165)
);

OA21x2_ASAP7_75t_L g3166 ( 
.A1(n_2852),
.A2(n_437),
.B(n_438),
.Y(n_3166)
);

INVx4_ASAP7_75t_L g3167 ( 
.A(n_2811),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2978),
.Y(n_3168)
);

OAI21x1_ASAP7_75t_L g3169 ( 
.A1(n_3109),
.A2(n_440),
.B(n_439),
.Y(n_3169)
);

HB1xp67_ASAP7_75t_L g3170 ( 
.A(n_2793),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2793),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2816),
.Y(n_3172)
);

OAI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2729),
.A2(n_440),
.B1(n_437),
.B2(n_439),
.Y(n_3173)
);

OR2x6_ASAP7_75t_L g3174 ( 
.A(n_2732),
.B(n_440),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2892),
.B(n_441),
.Y(n_3175)
);

INVx4_ASAP7_75t_L g3176 ( 
.A(n_2860),
.Y(n_3176)
);

AOI21xp33_ASAP7_75t_L g3177 ( 
.A1(n_3032),
.A2(n_441),
.B(n_442),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2823),
.B(n_2923),
.Y(n_3178)
);

AOI21xp5_ASAP7_75t_L g3179 ( 
.A1(n_2812),
.A2(n_442),
.B(n_443),
.Y(n_3179)
);

HB1xp67_ASAP7_75t_L g3180 ( 
.A(n_2816),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2842),
.B(n_442),
.Y(n_3181)
);

OAI22xp33_ASAP7_75t_L g3182 ( 
.A1(n_2904),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_3182)
);

BUFx12f_ASAP7_75t_L g3183 ( 
.A(n_2858),
.Y(n_3183)
);

AOI21xp33_ASAP7_75t_L g3184 ( 
.A1(n_2895),
.A2(n_443),
.B(n_444),
.Y(n_3184)
);

AOI22xp33_ASAP7_75t_L g3185 ( 
.A1(n_2860),
.A2(n_2904),
.B1(n_3058),
.B2(n_2961),
.Y(n_3185)
);

OAI21x1_ASAP7_75t_L g3186 ( 
.A1(n_3109),
.A2(n_447),
.B(n_446),
.Y(n_3186)
);

INVx1_ASAP7_75t_SL g3187 ( 
.A(n_3094),
.Y(n_3187)
);

OAI21x1_ASAP7_75t_L g3188 ( 
.A1(n_2887),
.A2(n_447),
.B(n_446),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3022),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2778),
.B(n_444),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3022),
.Y(n_3191)
);

A2O1A1Ixp33_ASAP7_75t_L g3192 ( 
.A1(n_2766),
.A2(n_448),
.B(n_446),
.C(n_447),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3022),
.Y(n_3193)
);

OAI21x1_ASAP7_75t_L g3194 ( 
.A1(n_2915),
.A2(n_450),
.B(n_449),
.Y(n_3194)
);

O2A1O1Ixp33_ASAP7_75t_L g3195 ( 
.A1(n_2874),
.A2(n_450),
.B(n_448),
.C(n_449),
.Y(n_3195)
);

INVxp67_ASAP7_75t_SL g3196 ( 
.A(n_2791),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2898),
.Y(n_3197)
);

AO32x2_ASAP7_75t_L g3198 ( 
.A1(n_2760),
.A2(n_453),
.A3(n_451),
.B1(n_452),
.B2(n_454),
.Y(n_3198)
);

OAI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_2804),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_3199)
);

AND2x6_ASAP7_75t_L g3200 ( 
.A(n_2768),
.B(n_454),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2843),
.A2(n_455),
.B(n_456),
.Y(n_3201)
);

NAND3xp33_ASAP7_75t_L g3202 ( 
.A(n_2911),
.B(n_455),
.C(n_457),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_2727),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.Y(n_3203)
);

BUFx4f_ASAP7_75t_SL g3204 ( 
.A(n_2901),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3041),
.Y(n_3205)
);

INVxp67_ASAP7_75t_L g3206 ( 
.A(n_3056),
.Y(n_3206)
);

BUFx2_ASAP7_75t_L g3207 ( 
.A(n_2736),
.Y(n_3207)
);

AOI221xp5_ASAP7_75t_L g3208 ( 
.A1(n_2864),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.C(n_460),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_2979),
.B(n_461),
.Y(n_3209)
);

NOR2x1p5_ASAP7_75t_L g3210 ( 
.A(n_2742),
.B(n_461),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2829),
.B(n_461),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_2787),
.B(n_462),
.Y(n_3212)
);

AOI21x1_ASAP7_75t_L g3213 ( 
.A1(n_2952),
.A2(n_559),
.B(n_558),
.Y(n_3213)
);

INVxp67_ASAP7_75t_L g3214 ( 
.A(n_3056),
.Y(n_3214)
);

INVx3_ASAP7_75t_L g3215 ( 
.A(n_2736),
.Y(n_3215)
);

AOI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_2860),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2830),
.A2(n_462),
.B(n_463),
.Y(n_3217)
);

BUFx4_ASAP7_75t_SL g3218 ( 
.A(n_3009),
.Y(n_3218)
);

OA21x2_ASAP7_75t_L g3219 ( 
.A1(n_2929),
.A2(n_463),
.B(n_466),
.Y(n_3219)
);

INVx3_ASAP7_75t_L g3220 ( 
.A(n_3118),
.Y(n_3220)
);

AO31x2_ASAP7_75t_L g3221 ( 
.A1(n_3004),
.A2(n_469),
.A3(n_466),
.B(n_468),
.Y(n_3221)
);

AO21x2_ASAP7_75t_L g3222 ( 
.A1(n_2734),
.A2(n_468),
.B(n_469),
.Y(n_3222)
);

AO21x2_ASAP7_75t_L g3223 ( 
.A1(n_2803),
.A2(n_469),
.B(n_470),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2741),
.B(n_470),
.Y(n_3224)
);

INVxp67_ASAP7_75t_L g3225 ( 
.A(n_2860),
.Y(n_3225)
);

OAI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_3112),
.A2(n_470),
.B(n_471),
.Y(n_3226)
);

INVx1_ASAP7_75t_SL g3227 ( 
.A(n_2754),
.Y(n_3227)
);

OA21x2_ASAP7_75t_L g3228 ( 
.A1(n_3045),
.A2(n_471),
.B(n_472),
.Y(n_3228)
);

O2A1O1Ixp33_ASAP7_75t_SL g3229 ( 
.A1(n_2726),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2866),
.B(n_474),
.Y(n_3230)
);

OAI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_3129),
.A2(n_474),
.B(n_475),
.Y(n_3231)
);

OA21x2_ASAP7_75t_L g3232 ( 
.A1(n_3049),
.A2(n_3059),
.B(n_2725),
.Y(n_3232)
);

CKINVDCx8_ASAP7_75t_R g3233 ( 
.A(n_2882),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2827),
.A2(n_475),
.B(n_476),
.Y(n_3234)
);

AO21x2_ASAP7_75t_L g3235 ( 
.A1(n_2987),
.A2(n_476),
.B(n_477),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2984),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_3236)
);

AO21x1_ASAP7_75t_L g3237 ( 
.A1(n_2730),
.A2(n_477),
.B(n_478),
.Y(n_3237)
);

CKINVDCx5p33_ASAP7_75t_R g3238 ( 
.A(n_3063),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2724),
.B(n_479),
.Y(n_3239)
);

OA21x2_ASAP7_75t_L g3240 ( 
.A1(n_2870),
.A2(n_481),
.B(n_483),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3054),
.Y(n_3241)
);

OAI221xp5_ASAP7_75t_L g3242 ( 
.A1(n_2747),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.C(n_486),
.Y(n_3242)
);

INVx1_ASAP7_75t_SL g3243 ( 
.A(n_2983),
.Y(n_3243)
);

HB1xp67_ASAP7_75t_L g3244 ( 
.A(n_2792),
.Y(n_3244)
);

OAI21x1_ASAP7_75t_SL g3245 ( 
.A1(n_3100),
.A2(n_484),
.B(n_485),
.Y(n_3245)
);

OAI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2992),
.A2(n_485),
.B(n_486),
.Y(n_3246)
);

INVx4_ASAP7_75t_L g3247 ( 
.A(n_2768),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2749),
.B(n_486),
.Y(n_3248)
);

OAI221xp5_ASAP7_75t_L g3249 ( 
.A1(n_2880),
.A2(n_3030),
.B1(n_2899),
.B2(n_2774),
.C(n_3035),
.Y(n_3249)
);

INVx2_ASAP7_75t_SL g3250 ( 
.A(n_2890),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2990),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_3251)
);

INVx5_ASAP7_75t_L g3252 ( 
.A(n_2768),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3019),
.Y(n_3253)
);

OR2x6_ASAP7_75t_L g3254 ( 
.A(n_2785),
.B(n_487),
.Y(n_3254)
);

AOI221xp5_ASAP7_75t_L g3255 ( 
.A1(n_2916),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.C(n_491),
.Y(n_3255)
);

AO21x2_ASAP7_75t_L g3256 ( 
.A1(n_2757),
.A2(n_490),
.B(n_491),
.Y(n_3256)
);

OR2x2_ASAP7_75t_L g3257 ( 
.A(n_2728),
.B(n_490),
.Y(n_3257)
);

AOI22xp33_ASAP7_75t_L g3258 ( 
.A1(n_3086),
.A2(n_3126),
.B1(n_2815),
.B2(n_3104),
.Y(n_3258)
);

AOI22x1_ASAP7_75t_L g3259 ( 
.A1(n_2767),
.A2(n_495),
.B1(n_492),
.B2(n_494),
.Y(n_3259)
);

BUFx10_ASAP7_75t_L g3260 ( 
.A(n_3039),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_2979),
.B(n_494),
.Y(n_3261)
);

OR2x6_ASAP7_75t_L g3262 ( 
.A(n_2805),
.B(n_495),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_2979),
.B(n_496),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3064),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_2731),
.B(n_496),
.Y(n_3265)
);

AO31x2_ASAP7_75t_L g3266 ( 
.A1(n_3055),
.A2(n_498),
.A3(n_496),
.B(n_497),
.Y(n_3266)
);

O2A1O1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_2879),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_3267)
);

NAND2x1p5_ASAP7_75t_L g3268 ( 
.A(n_2959),
.B(n_498),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2841),
.B(n_499),
.Y(n_3269)
);

AOI21xp33_ASAP7_75t_L g3270 ( 
.A1(n_2863),
.A2(n_499),
.B(n_500),
.Y(n_3270)
);

AO21x2_ASAP7_75t_L g3271 ( 
.A1(n_3011),
.A2(n_500),
.B(n_501),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3020),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3064),
.Y(n_3273)
);

OAI22xp5_ASAP7_75t_SL g3274 ( 
.A1(n_2920),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2847),
.B(n_502),
.Y(n_3275)
);

OA21x2_ASAP7_75t_L g3276 ( 
.A1(n_2738),
.A2(n_2740),
.B(n_2918),
.Y(n_3276)
);

HB1xp67_ASAP7_75t_L g3277 ( 
.A(n_2813),
.Y(n_3277)
);

CKINVDCx16_ASAP7_75t_R g3278 ( 
.A(n_3038),
.Y(n_3278)
);

AOI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_2788),
.A2(n_504),
.B(n_505),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3108),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3108),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3108),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2790),
.B(n_506),
.Y(n_3283)
);

OA21x2_ASAP7_75t_L g3284 ( 
.A1(n_2797),
.A2(n_506),
.B(n_507),
.Y(n_3284)
);

NAND2x1p5_ASAP7_75t_L g3285 ( 
.A(n_2824),
.B(n_507),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2903),
.Y(n_3286)
);

HB1xp67_ASAP7_75t_L g3287 ( 
.A(n_2833),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2993),
.B(n_509),
.Y(n_3288)
);

BUFx3_ASAP7_75t_L g3289 ( 
.A(n_2917),
.Y(n_3289)
);

A2O1A1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_3116),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_3290)
);

AO21x2_ASAP7_75t_L g3291 ( 
.A1(n_2897),
.A2(n_511),
.B(n_512),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_3118),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2903),
.Y(n_3293)
);

OA21x2_ASAP7_75t_L g3294 ( 
.A1(n_3046),
.A2(n_3034),
.B(n_3029),
.Y(n_3294)
);

OAI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3017),
.A2(n_512),
.B(n_513),
.Y(n_3295)
);

AO21x2_ASAP7_75t_L g3296 ( 
.A1(n_2919),
.A2(n_513),
.B(n_514),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2845),
.A2(n_516),
.B(n_517),
.Y(n_3297)
);

OAI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_3101),
.A2(n_518),
.B(n_519),
.Y(n_3298)
);

INVx3_ASAP7_75t_L g3299 ( 
.A(n_2824),
.Y(n_3299)
);

BUFx2_ASAP7_75t_SL g3300 ( 
.A(n_2969),
.Y(n_3300)
);

OAI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_2872),
.A2(n_518),
.B(n_520),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_SL g3302 ( 
.A(n_3122),
.B(n_518),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2739),
.Y(n_3303)
);

INVxp33_ASAP7_75t_L g3304 ( 
.A(n_2777),
.Y(n_3304)
);

OR2x6_ASAP7_75t_L g3305 ( 
.A(n_2819),
.B(n_521),
.Y(n_3305)
);

OR2x6_ASAP7_75t_L g3306 ( 
.A(n_3038),
.B(n_522),
.Y(n_3306)
);

OAI21x1_ASAP7_75t_L g3307 ( 
.A1(n_3048),
.A2(n_523),
.B(n_524),
.Y(n_3307)
);

AO32x2_ASAP7_75t_L g3308 ( 
.A1(n_2828),
.A2(n_525),
.A3(n_523),
.B1(n_524),
.B2(n_526),
.Y(n_3308)
);

INVxp67_ASAP7_75t_SL g3309 ( 
.A(n_2824),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_2941),
.B(n_523),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_SL g3311 ( 
.A1(n_2770),
.A2(n_524),
.B(n_525),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2945),
.A2(n_525),
.B(n_526),
.Y(n_3312)
);

OAI21x1_ASAP7_75t_SL g3313 ( 
.A1(n_2996),
.A2(n_526),
.B(n_527),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2903),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_2851),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3077),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_3316)
);

AND2x4_ASAP7_75t_L g3317 ( 
.A(n_3106),
.B(n_530),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2930),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_2930),
.Y(n_3319)
);

AND2x2_ASAP7_75t_L g3320 ( 
.A(n_2912),
.B(n_532),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_2862),
.A2(n_533),
.B(n_534),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3099),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_3322)
);

BUFx2_ASAP7_75t_L g3323 ( 
.A(n_2981),
.Y(n_3323)
);

A2O1A1Ixp33_ASAP7_75t_L g3324 ( 
.A1(n_3000),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_3324)
);

INVx3_ASAP7_75t_L g3325 ( 
.A(n_2890),
.Y(n_3325)
);

OAI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3091),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_3326)
);

NAND2xp33_ASAP7_75t_SL g3327 ( 
.A(n_3005),
.B(n_538),
.Y(n_3327)
);

OAI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_2951),
.A2(n_539),
.B1(n_560),
.B2(n_559),
.Y(n_3328)
);

AND2x4_ASAP7_75t_L g3329 ( 
.A(n_3106),
.B(n_561),
.Y(n_3329)
);

OAI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3091),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_3330)
);

AND2x4_ASAP7_75t_L g3331 ( 
.A(n_3106),
.B(n_565),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2739),
.Y(n_3332)
);

OAI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_3097),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_3333)
);

INVx2_ASAP7_75t_SL g3334 ( 
.A(n_2983),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3003),
.Y(n_3335)
);

OR3x4_ASAP7_75t_SL g3336 ( 
.A(n_2789),
.B(n_568),
.C(n_570),
.Y(n_3336)
);

AO21x2_ASAP7_75t_L g3337 ( 
.A1(n_3037),
.A2(n_570),
.B(n_571),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2927),
.B(n_571),
.Y(n_3338)
);

NAND2x1p5_ASAP7_75t_L g3339 ( 
.A(n_2851),
.B(n_2853),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_2821),
.A2(n_576),
.B1(n_572),
.B2(n_574),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_2821),
.A2(n_578),
.B1(n_574),
.B2(n_577),
.Y(n_3341)
);

NOR2x1_ASAP7_75t_SL g3342 ( 
.A(n_3113),
.B(n_579),
.Y(n_3342)
);

OAI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_2857),
.A2(n_582),
.B1(n_579),
.B2(n_581),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2900),
.B(n_973),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_2888),
.A2(n_584),
.B1(n_581),
.B2(n_583),
.Y(n_3345)
);

OAI21x1_ASAP7_75t_SL g3346 ( 
.A1(n_2859),
.A2(n_583),
.B(n_584),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_SL g3347 ( 
.A1(n_2853),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_3347)
);

AND2x4_ASAP7_75t_L g3348 ( 
.A(n_2810),
.B(n_2814),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2925),
.B(n_2906),
.Y(n_3349)
);

AO31x2_ASAP7_75t_L g3350 ( 
.A1(n_3084),
.A2(n_590),
.A3(n_588),
.B(n_589),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_3053),
.Y(n_3351)
);

NAND2x1p5_ASAP7_75t_L g3352 ( 
.A(n_2773),
.B(n_590),
.Y(n_3352)
);

OAI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_3001),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.Y(n_3353)
);

OAI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3071),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_L g3355 ( 
.A1(n_3128),
.A2(n_602),
.B1(n_598),
.B2(n_599),
.Y(n_3355)
);

OAI21x1_ASAP7_75t_L g3356 ( 
.A1(n_2937),
.A2(n_2960),
.B(n_2744),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3042),
.A2(n_3124),
.B(n_3050),
.Y(n_3357)
);

BUFx3_ASAP7_75t_L g3358 ( 
.A(n_2948),
.Y(n_3358)
);

AOI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_2949),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2818),
.Y(n_3360)
);

NOR3xp33_ASAP7_75t_L g3361 ( 
.A(n_2752),
.B(n_603),
.C(n_604),
.Y(n_3361)
);

OR2x6_ASAP7_75t_L g3362 ( 
.A(n_2826),
.B(n_605),
.Y(n_3362)
);

INVx3_ASAP7_75t_L g3363 ( 
.A(n_2935),
.Y(n_3363)
);

OR2x6_ASAP7_75t_L g3364 ( 
.A(n_2844),
.B(n_606),
.Y(n_3364)
);

INVx4_ASAP7_75t_L g3365 ( 
.A(n_2968),
.Y(n_3365)
);

OAI21x1_ASAP7_75t_L g3366 ( 
.A1(n_2735),
.A2(n_2796),
.B(n_2753),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_2808),
.B(n_606),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_2755),
.Y(n_3368)
);

OA21x2_ASAP7_75t_L g3369 ( 
.A1(n_2913),
.A2(n_3080),
.B(n_3010),
.Y(n_3369)
);

BUFx2_ASAP7_75t_L g3370 ( 
.A(n_2909),
.Y(n_3370)
);

NAND2xp33_ASAP7_75t_L g3371 ( 
.A(n_2822),
.B(n_607),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_3070),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_3372)
);

OR2x6_ASAP7_75t_L g3373 ( 
.A(n_2975),
.B(n_609),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2755),
.Y(n_3374)
);

OAI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_2873),
.A2(n_610),
.B(n_611),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2963),
.Y(n_3376)
);

O2A1O1Ixp33_ASAP7_75t_SL g3377 ( 
.A1(n_2746),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2755),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_2928),
.B(n_972),
.Y(n_3379)
);

O2A1O1Ixp33_ASAP7_75t_L g3380 ( 
.A1(n_2802),
.A2(n_616),
.B(n_614),
.C(n_615),
.Y(n_3380)
);

OA21x2_ASAP7_75t_L g3381 ( 
.A1(n_2779),
.A2(n_618),
.B(n_619),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2832),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2832),
.Y(n_3383)
);

NOR2x1_ASAP7_75t_R g3384 ( 
.A(n_3007),
.B(n_619),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2832),
.Y(n_3385)
);

NOR2xp67_ASAP7_75t_L g3386 ( 
.A(n_3057),
.B(n_620),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2881),
.B(n_2883),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2884),
.B(n_972),
.Y(n_3388)
);

OA21x2_ASAP7_75t_L g3389 ( 
.A1(n_2780),
.A2(n_622),
.B(n_623),
.Y(n_3389)
);

A2O1A1Ixp33_ASAP7_75t_L g3390 ( 
.A1(n_2781),
.A2(n_626),
.B(n_624),
.C(n_625),
.Y(n_3390)
);

NOR2x1_ASAP7_75t_R g3391 ( 
.A(n_3007),
.B(n_628),
.Y(n_3391)
);

AO21x2_ASAP7_75t_L g3392 ( 
.A1(n_2745),
.A2(n_2809),
.B(n_3103),
.Y(n_3392)
);

A2O1A1Ixp33_ASAP7_75t_L g3393 ( 
.A1(n_3090),
.A2(n_631),
.B(n_629),
.C(n_630),
.Y(n_3393)
);

BUFx2_ASAP7_75t_L g3394 ( 
.A(n_2909),
.Y(n_3394)
);

OAI21x1_ASAP7_75t_L g3395 ( 
.A1(n_3088),
.A2(n_629),
.B(n_630),
.Y(n_3395)
);

BUFx4f_ASAP7_75t_L g3396 ( 
.A(n_3008),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2885),
.B(n_632),
.Y(n_3397)
);

OR2x2_ASAP7_75t_L g3398 ( 
.A(n_2748),
.B(n_633),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3092),
.A2(n_633),
.B(n_635),
.Y(n_3399)
);

OAI21x1_ASAP7_75t_L g3400 ( 
.A1(n_3093),
.A2(n_635),
.B(n_636),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_2869),
.B(n_638),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3102),
.A2(n_638),
.B(n_639),
.Y(n_3402)
);

INVx2_ASAP7_75t_SL g3403 ( 
.A(n_3008),
.Y(n_3403)
);

AOI21x1_ASAP7_75t_L g3404 ( 
.A1(n_3114),
.A2(n_639),
.B(n_640),
.Y(n_3404)
);

NAND2x1p5_ASAP7_75t_L g3405 ( 
.A(n_3012),
.B(n_971),
.Y(n_3405)
);

O2A1O1Ixp33_ASAP7_75t_SL g3406 ( 
.A1(n_2784),
.A2(n_643),
.B(n_641),
.C(n_642),
.Y(n_3406)
);

AOI221xp5_ASAP7_75t_L g3407 ( 
.A1(n_2876),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.C(n_647),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2761),
.Y(n_3408)
);

AO31x2_ASAP7_75t_L g3409 ( 
.A1(n_2886),
.A2(n_650),
.A3(n_648),
.B(n_649),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2761),
.Y(n_3410)
);

OA21x2_ASAP7_75t_L g3411 ( 
.A1(n_2849),
.A2(n_648),
.B(n_649),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2893),
.Y(n_3412)
);

AND2x4_ASAP7_75t_L g3413 ( 
.A(n_2935),
.B(n_3015),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2910),
.Y(n_3414)
);

INVx3_ASAP7_75t_SL g3415 ( 
.A(n_3012),
.Y(n_3415)
);

OR2x6_ASAP7_75t_L g3416 ( 
.A(n_2806),
.B(n_650),
.Y(n_3416)
);

OR2x2_ASAP7_75t_L g3417 ( 
.A(n_2750),
.B(n_651),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_2924),
.Y(n_3418)
);

AOI222xp33_ASAP7_75t_L g3419 ( 
.A1(n_2871),
.A2(n_654),
.B1(n_656),
.B2(n_651),
.C1(n_652),
.C2(n_655),
.Y(n_3419)
);

CKINVDCx5p33_ASAP7_75t_R g3420 ( 
.A(n_3065),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_2889),
.B(n_659),
.Y(n_3421)
);

OAI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_2914),
.A2(n_659),
.B(n_660),
.Y(n_3422)
);

INVx3_ASAP7_75t_L g3423 ( 
.A(n_2935),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3015),
.B(n_660),
.Y(n_3424)
);

BUFx2_ASAP7_75t_L g3425 ( 
.A(n_3066),
.Y(n_3425)
);

AOI22x1_ASAP7_75t_L g3426 ( 
.A1(n_3087),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_3426)
);

BUFx2_ASAP7_75t_L g3427 ( 
.A(n_3015),
.Y(n_3427)
);

OA21x2_ASAP7_75t_L g3428 ( 
.A1(n_2825),
.A2(n_666),
.B(n_667),
.Y(n_3428)
);

AOI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_2947),
.A2(n_669),
.B(n_671),
.Y(n_3429)
);

OAI21x1_ASAP7_75t_SL g3430 ( 
.A1(n_2986),
.A2(n_2999),
.B(n_2988),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2765),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3040),
.B(n_669),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3053),
.Y(n_3433)
);

AND2x4_ASAP7_75t_L g3434 ( 
.A(n_2964),
.B(n_672),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3044),
.B(n_2758),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3115),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_3436)
);

NAND2x1p5_ASAP7_75t_L g3437 ( 
.A(n_2875),
.B(n_970),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_SL g3438 ( 
.A1(n_2867),
.A2(n_673),
.B(n_674),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2891),
.B(n_970),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_2905),
.Y(n_3440)
);

AO21x2_ASAP7_75t_L g3441 ( 
.A1(n_3047),
.A2(n_675),
.B(n_676),
.Y(n_3441)
);

AOI22xp33_ASAP7_75t_L g3442 ( 
.A1(n_3117),
.A2(n_677),
.B1(n_675),
.B2(n_676),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2765),
.Y(n_3443)
);

OAI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_2838),
.A2(n_677),
.B(n_678),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_2782),
.Y(n_3445)
);

AO31x2_ASAP7_75t_L g3446 ( 
.A1(n_2939),
.A2(n_682),
.A3(n_679),
.B(n_681),
.Y(n_3446)
);

OAI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_2839),
.A2(n_3033),
.B(n_3027),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3117),
.A2(n_685),
.B1(n_682),
.B2(n_684),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_2902),
.B(n_685),
.Y(n_3449)
);

INVx6_ASAP7_75t_L g3450 ( 
.A(n_3026),
.Y(n_3450)
);

NAND2x1p5_ASAP7_75t_L g3451 ( 
.A(n_3074),
.B(n_969),
.Y(n_3451)
);

NAND3xp33_ASAP7_75t_L g3452 ( 
.A(n_3111),
.B(n_686),
.C(n_687),
.Y(n_3452)
);

INVx1_ASAP7_75t_SL g3453 ( 
.A(n_2998),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_2782),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_2762),
.B(n_688),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_2782),
.Y(n_3456)
);

OAI21x1_ASAP7_75t_L g3457 ( 
.A1(n_3014),
.A2(n_689),
.B(n_691),
.Y(n_3457)
);

O2A1O1Ixp33_ASAP7_75t_L g3458 ( 
.A1(n_2907),
.A2(n_693),
.B(n_691),
.C(n_692),
.Y(n_3458)
);

INVx2_ASAP7_75t_SL g3459 ( 
.A(n_3036),
.Y(n_3459)
);

OAI21x1_ASAP7_75t_L g3460 ( 
.A1(n_3051),
.A2(n_692),
.B(n_694),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_2946),
.B(n_3002),
.Y(n_3461)
);

AND2x2_ASAP7_75t_SL g3462 ( 
.A(n_2940),
.B(n_695),
.Y(n_3462)
);

AND2x4_ASAP7_75t_L g3463 ( 
.A(n_3028),
.B(n_695),
.Y(n_3463)
);

OAI21x1_ASAP7_75t_L g3464 ( 
.A1(n_3081),
.A2(n_696),
.B(n_697),
.Y(n_3464)
);

HB1xp67_ASAP7_75t_L g3465 ( 
.A(n_3025),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3069),
.Y(n_3466)
);

BUFx3_ASAP7_75t_L g3467 ( 
.A(n_2965),
.Y(n_3467)
);

AOI21x1_ASAP7_75t_L g3468 ( 
.A1(n_2798),
.A2(n_696),
.B(n_697),
.Y(n_3468)
);

INVx1_ASAP7_75t_SL g3469 ( 
.A(n_2855),
.Y(n_3469)
);

INVx4_ASAP7_75t_L g3470 ( 
.A(n_3026),
.Y(n_3470)
);

OAI21x1_ASAP7_75t_L g3471 ( 
.A1(n_3083),
.A2(n_698),
.B(n_699),
.Y(n_3471)
);

AND2x4_ASAP7_75t_L g3472 ( 
.A(n_2933),
.B(n_700),
.Y(n_3472)
);

OAI22xp5_ASAP7_75t_L g3473 ( 
.A1(n_3095),
.A2(n_2854),
.B1(n_2865),
.B2(n_2771),
.Y(n_3473)
);

CKINVDCx5p33_ASAP7_75t_R g3474 ( 
.A(n_2776),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_2769),
.B(n_700),
.Y(n_3475)
);

OR2x2_ASAP7_75t_L g3476 ( 
.A(n_2783),
.B(n_702),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3087),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3072),
.Y(n_3478)
);

AOI21x1_ASAP7_75t_L g3479 ( 
.A1(n_2799),
.A2(n_702),
.B(n_703),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3024),
.B(n_704),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2775),
.Y(n_3481)
);

AND2x4_ASAP7_75t_L g3482 ( 
.A(n_2976),
.B(n_704),
.Y(n_3482)
);

AOI21x1_ASAP7_75t_L g3483 ( 
.A1(n_2800),
.A2(n_705),
.B(n_706),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3021),
.B(n_705),
.Y(n_3484)
);

OAI21x1_ASAP7_75t_L g3485 ( 
.A1(n_3085),
.A2(n_706),
.B(n_707),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_3026),
.B(n_707),
.Y(n_3486)
);

AND2x4_ASAP7_75t_L g3487 ( 
.A(n_2942),
.B(n_709),
.Y(n_3487)
);

OAI21x1_ASAP7_75t_L g3488 ( 
.A1(n_3098),
.A2(n_3110),
.B(n_3107),
.Y(n_3488)
);

OR2x6_ASAP7_75t_L g3489 ( 
.A(n_2908),
.B(n_711),
.Y(n_3489)
);

AOI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3121),
.A2(n_3068),
.B1(n_3062),
.B2(n_3018),
.Y(n_3490)
);

OA21x2_ASAP7_75t_L g3491 ( 
.A1(n_3052),
.A2(n_714),
.B(n_716),
.Y(n_3491)
);

CKINVDCx12_ASAP7_75t_R g3492 ( 
.A(n_3127),
.Y(n_3492)
);

OAI21x1_ASAP7_75t_L g3493 ( 
.A1(n_2801),
.A2(n_717),
.B(n_718),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3073),
.Y(n_3494)
);

OAI21x1_ASAP7_75t_L g3495 ( 
.A1(n_2807),
.A2(n_719),
.B(n_720),
.Y(n_3495)
);

AND2x4_ASAP7_75t_L g3496 ( 
.A(n_3006),
.B(n_719),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2922),
.B(n_721),
.Y(n_3497)
);

CKINVDCx8_ASAP7_75t_R g3498 ( 
.A(n_3006),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3013),
.Y(n_3499)
);

INVx3_ASAP7_75t_L g3500 ( 
.A(n_3053),
.Y(n_3500)
);

INVx2_ASAP7_75t_SL g3501 ( 
.A(n_3078),
.Y(n_3501)
);

NOR2xp67_ASAP7_75t_L g3502 ( 
.A(n_2970),
.B(n_721),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3125),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3006),
.B(n_722),
.Y(n_3504)
);

INVxp67_ASAP7_75t_L g3505 ( 
.A(n_3079),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_2953),
.B(n_723),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_2982),
.B(n_723),
.Y(n_3507)
);

INVx3_ASAP7_75t_SL g3508 ( 
.A(n_2955),
.Y(n_3508)
);

INVx3_ASAP7_75t_L g3509 ( 
.A(n_2955),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2991),
.Y(n_3510)
);

BUFx6f_ASAP7_75t_L g3511 ( 
.A(n_2955),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_2973),
.B(n_724),
.Y(n_3512)
);

NAND3xp33_ASAP7_75t_L g3513 ( 
.A(n_3096),
.B(n_2850),
.C(n_3016),
.Y(n_3513)
);

AOI22x1_ASAP7_75t_L g3514 ( 
.A1(n_3061),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2820),
.B(n_725),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3123),
.Y(n_3516)
);

OAI21x1_ASAP7_75t_L g3517 ( 
.A1(n_2834),
.A2(n_726),
.B(n_727),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_2896),
.B(n_2931),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_2994),
.B(n_3060),
.Y(n_3519)
);

INVx3_ASAP7_75t_L g3520 ( 
.A(n_2989),
.Y(n_3520)
);

OAI21x1_ASAP7_75t_L g3521 ( 
.A1(n_2835),
.A2(n_728),
.B(n_729),
.Y(n_3521)
);

OA21x2_ASAP7_75t_L g3522 ( 
.A1(n_3076),
.A2(n_728),
.B(n_730),
.Y(n_3522)
);

BUFx6f_ASAP7_75t_L g3523 ( 
.A(n_3151),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3148),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3148),
.Y(n_3525)
);

OR2x2_ASAP7_75t_L g3526 ( 
.A(n_3152),
.B(n_2837),
.Y(n_3526)
);

AND2x4_ASAP7_75t_L g3527 ( 
.A(n_3176),
.B(n_2989),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3141),
.Y(n_3528)
);

BUFx6f_ASAP7_75t_L g3529 ( 
.A(n_3151),
.Y(n_3529)
);

INVxp67_ASAP7_75t_SL g3530 ( 
.A(n_3176),
.Y(n_3530)
);

OR2x2_ASAP7_75t_L g3531 ( 
.A(n_3278),
.B(n_2848),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3157),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_3151),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3149),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3157),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3412),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3181),
.B(n_730),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3414),
.Y(n_3538)
);

INVx3_ASAP7_75t_L g3539 ( 
.A(n_3167),
.Y(n_3539)
);

INVx1_ASAP7_75t_SL g3540 ( 
.A(n_3218),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3505),
.B(n_2934),
.Y(n_3541)
);

OR2x2_ASAP7_75t_L g3542 ( 
.A(n_3257),
.B(n_2894),
.Y(n_3542)
);

CKINVDCx20_ASAP7_75t_R g3543 ( 
.A(n_3204),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3159),
.Y(n_3544)
);

AO21x2_ASAP7_75t_L g3545 ( 
.A1(n_3360),
.A2(n_3105),
.B(n_2980),
.Y(n_3545)
);

HB1xp67_ASAP7_75t_L g3546 ( 
.A(n_3170),
.Y(n_3546)
);

CKINVDCx5p33_ASAP7_75t_R g3547 ( 
.A(n_3183),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3159),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3163),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3163),
.Y(n_3550)
);

HB1xp67_ASAP7_75t_L g3551 ( 
.A(n_3180),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3165),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3418),
.Y(n_3553)
);

OR2x2_ASAP7_75t_L g3554 ( 
.A(n_3190),
.B(n_3075),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3466),
.Y(n_3555)
);

OA21x2_ASAP7_75t_L g3556 ( 
.A1(n_3156),
.A2(n_2950),
.B(n_2926),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3165),
.Y(n_3557)
);

BUFx2_ASAP7_75t_L g3558 ( 
.A(n_3207),
.Y(n_3558)
);

INVxp33_ASAP7_75t_L g3559 ( 
.A(n_3384),
.Y(n_3559)
);

HB1xp67_ASAP7_75t_L g3560 ( 
.A(n_3244),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3212),
.B(n_732),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3478),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_3277),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3494),
.Y(n_3564)
);

OR2x6_ASAP7_75t_L g3565 ( 
.A(n_3306),
.B(n_2962),
.Y(n_3565)
);

HB1xp67_ASAP7_75t_L g3566 ( 
.A(n_3287),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3376),
.Y(n_3567)
);

AND2x4_ASAP7_75t_L g3568 ( 
.A(n_3225),
.B(n_2989),
.Y(n_3568)
);

AND2x4_ASAP7_75t_L g3569 ( 
.A(n_3477),
.B(n_3067),
.Y(n_3569)
);

AO21x2_ASAP7_75t_L g3570 ( 
.A1(n_3357),
.A2(n_2971),
.B(n_2921),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3477),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3440),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3516),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3169),
.Y(n_3574)
);

OA21x2_ASAP7_75t_L g3575 ( 
.A1(n_3189),
.A2(n_2868),
.B(n_3089),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3265),
.B(n_732),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3465),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3344),
.Y(n_3578)
);

INVx3_ASAP7_75t_L g3579 ( 
.A(n_3167),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3186),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3261),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3261),
.Y(n_3582)
);

INVx2_ASAP7_75t_SL g3583 ( 
.A(n_3260),
.Y(n_3583)
);

INVx2_ASAP7_75t_SL g3584 ( 
.A(n_3260),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3263),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3263),
.Y(n_3586)
);

BUFx2_ASAP7_75t_L g3587 ( 
.A(n_3323),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3367),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3367),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3435),
.B(n_733),
.Y(n_3590)
);

O2A1O1Ixp5_ASAP7_75t_L g3591 ( 
.A1(n_3396),
.A2(n_3082),
.B(n_2938),
.C(n_2985),
.Y(n_3591)
);

NOR2xp67_ASAP7_75t_R g3592 ( 
.A(n_3220),
.B(n_3067),
.Y(n_3592)
);

INVx6_ASAP7_75t_L g3593 ( 
.A(n_3306),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3303),
.Y(n_3594)
);

INVxp67_ASAP7_75t_L g3595 ( 
.A(n_3391),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3320),
.B(n_733),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3138),
.A2(n_3462),
.B1(n_3254),
.B2(n_3305),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3432),
.B(n_734),
.Y(n_3598)
);

OR2x2_ASAP7_75t_L g3599 ( 
.A(n_3469),
.B(n_3453),
.Y(n_3599)
);

AO21x2_ASAP7_75t_L g3600 ( 
.A1(n_3246),
.A2(n_3120),
.B(n_2997),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3221),
.Y(n_3601)
);

OR2x6_ASAP7_75t_L g3602 ( 
.A(n_3300),
.B(n_2836),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3303),
.Y(n_3603)
);

INVx1_ASAP7_75t_SL g3604 ( 
.A(n_3243),
.Y(n_3604)
);

BUFx4f_ASAP7_75t_SL g3605 ( 
.A(n_3187),
.Y(n_3605)
);

INVx3_ASAP7_75t_L g3606 ( 
.A(n_3147),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_3332),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3221),
.Y(n_3608)
);

BUFx2_ASAP7_75t_L g3609 ( 
.A(n_3415),
.Y(n_3609)
);

INVxp67_ASAP7_75t_SL g3610 ( 
.A(n_3339),
.Y(n_3610)
);

INVx3_ASAP7_75t_L g3611 ( 
.A(n_3147),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3221),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3266),
.Y(n_3613)
);

AO21x2_ASAP7_75t_L g3614 ( 
.A1(n_3226),
.A2(n_3231),
.B(n_3191),
.Y(n_3614)
);

HB1xp67_ASAP7_75t_L g3615 ( 
.A(n_3403),
.Y(n_3615)
);

INVxp67_ASAP7_75t_SL g3616 ( 
.A(n_3396),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3266),
.Y(n_3617)
);

AO21x2_ASAP7_75t_L g3618 ( 
.A1(n_3189),
.A2(n_2956),
.B(n_2977),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3459),
.B(n_734),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3266),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3332),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3434),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3434),
.Y(n_3623)
);

CKINVDCx16_ASAP7_75t_R g3624 ( 
.A(n_3358),
.Y(n_3624)
);

OA21x2_ASAP7_75t_L g3625 ( 
.A1(n_3191),
.A2(n_2967),
.B(n_2943),
.Y(n_3625)
);

CKINVDCx6p67_ASAP7_75t_R g3626 ( 
.A(n_3492),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3472),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3472),
.Y(n_3628)
);

OR2x2_ASAP7_75t_L g3629 ( 
.A(n_3227),
.B(n_2936),
.Y(n_3629)
);

BUFx2_ASAP7_75t_L g3630 ( 
.A(n_3220),
.Y(n_3630)
);

INVx3_ASAP7_75t_L g3631 ( 
.A(n_3215),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3370),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3394),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3269),
.Y(n_3634)
);

OAI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3513),
.A2(n_2954),
.B(n_3023),
.Y(n_3635)
);

AND2x4_ASAP7_75t_L g3636 ( 
.A(n_3215),
.B(n_3067),
.Y(n_3636)
);

INVx2_ASAP7_75t_SL g3637 ( 
.A(n_3289),
.Y(n_3637)
);

INVx3_ASAP7_75t_SL g3638 ( 
.A(n_3238),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3275),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3463),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3463),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3467),
.B(n_969),
.Y(n_3642)
);

AND2x4_ASAP7_75t_L g3643 ( 
.A(n_3424),
.B(n_736),
.Y(n_3643)
);

AND2x2_ASAP7_75t_L g3644 ( 
.A(n_3401),
.B(n_736),
.Y(n_3644)
);

AO21x2_ASAP7_75t_L g3645 ( 
.A1(n_3193),
.A2(n_737),
.B(n_738),
.Y(n_3645)
);

OA21x2_ASAP7_75t_L g3646 ( 
.A1(n_3193),
.A2(n_737),
.B(n_739),
.Y(n_3646)
);

INVx3_ASAP7_75t_L g3647 ( 
.A(n_3292),
.Y(n_3647)
);

OAI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3390),
.A2(n_3393),
.B(n_3298),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_3252),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3162),
.Y(n_3650)
);

INVx3_ASAP7_75t_L g3651 ( 
.A(n_3292),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3205),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3205),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_3130),
.A2(n_740),
.B(n_741),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3241),
.Y(n_3655)
);

INVx1_ASAP7_75t_SL g3656 ( 
.A(n_3334),
.Y(n_3656)
);

HB1xp67_ASAP7_75t_L g3657 ( 
.A(n_3233),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3264),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3420),
.B(n_742),
.Y(n_3659)
);

INVx4_ASAP7_75t_L g3660 ( 
.A(n_3200),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3264),
.Y(n_3661)
);

INVx3_ASAP7_75t_L g3662 ( 
.A(n_3325),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3273),
.Y(n_3663)
);

INVx3_ASAP7_75t_L g3664 ( 
.A(n_3325),
.Y(n_3664)
);

BUFx2_ASAP7_75t_SL g3665 ( 
.A(n_3200),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3349),
.B(n_744),
.Y(n_3666)
);

OAI22xp5_ASAP7_75t_L g3667 ( 
.A1(n_3136),
.A2(n_747),
.B1(n_745),
.B2(n_746),
.Y(n_3667)
);

INVx3_ASAP7_75t_L g3668 ( 
.A(n_3498),
.Y(n_3668)
);

OR2x6_ASAP7_75t_L g3669 ( 
.A(n_3362),
.B(n_745),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3175),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3230),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3482),
.Y(n_3672)
);

INVx3_ASAP7_75t_L g3673 ( 
.A(n_3138),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3482),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3487),
.Y(n_3675)
);

OA21x2_ASAP7_75t_L g3676 ( 
.A1(n_3280),
.A2(n_748),
.B(n_749),
.Y(n_3676)
);

OR2x2_ASAP7_75t_L g3677 ( 
.A(n_3132),
.B(n_748),
.Y(n_3677)
);

AND2x4_ASAP7_75t_L g3678 ( 
.A(n_3424),
.B(n_750),
.Y(n_3678)
);

BUFx3_ASAP7_75t_L g3679 ( 
.A(n_3508),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3487),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3501),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3171),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3172),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3510),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3350),
.Y(n_3685)
);

BUFx3_ASAP7_75t_L g3686 ( 
.A(n_3365),
.Y(n_3686)
);

OAI22xp5_ASAP7_75t_L g3687 ( 
.A1(n_3185),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3281),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3206),
.B(n_751),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3282),
.Y(n_3690)
);

HB1xp67_ASAP7_75t_L g3691 ( 
.A(n_3196),
.Y(n_3691)
);

BUFx6f_ASAP7_75t_L g3692 ( 
.A(n_3252),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3131),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3131),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3475),
.B(n_752),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3382),
.Y(n_3696)
);

INVx2_ASAP7_75t_SL g3697 ( 
.A(n_3365),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3295),
.A2(n_968),
.B(n_754),
.Y(n_3698)
);

INVxp67_ASAP7_75t_L g3699 ( 
.A(n_3178),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3133),
.Y(n_3700)
);

BUFx6f_ASAP7_75t_L g3701 ( 
.A(n_3252),
.Y(n_3701)
);

NAND2x1p5_ASAP7_75t_L g3702 ( 
.A(n_3250),
.B(n_755),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3518),
.B(n_756),
.Y(n_3703)
);

AOI21x1_ASAP7_75t_L g3704 ( 
.A1(n_3164),
.A2(n_756),
.B(n_757),
.Y(n_3704)
);

HB1xp67_ASAP7_75t_L g3705 ( 
.A(n_3214),
.Y(n_3705)
);

BUFx8_ASAP7_75t_L g3706 ( 
.A(n_3200),
.Y(n_3706)
);

OAI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3145),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3382),
.Y(n_3708)
);

INVx4_ASAP7_75t_L g3709 ( 
.A(n_3200),
.Y(n_3709)
);

AND2x4_ASAP7_75t_L g3710 ( 
.A(n_3329),
.B(n_761),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3383),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3133),
.Y(n_3712)
);

INVx3_ASAP7_75t_L g3713 ( 
.A(n_3247),
.Y(n_3713)
);

BUFx8_ASAP7_75t_L g3714 ( 
.A(n_3425),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3254),
.B(n_3262),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3134),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3350),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3262),
.B(n_968),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3350),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3383),
.Y(n_3720)
);

HB1xp67_ASAP7_75t_L g3721 ( 
.A(n_3317),
.Y(n_3721)
);

INVx3_ASAP7_75t_L g3722 ( 
.A(n_3247),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3409),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3409),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3385),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3385),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3409),
.Y(n_3727)
);

O2A1O1Ixp5_ASAP7_75t_L g3728 ( 
.A1(n_3153),
.A2(n_765),
.B(n_762),
.C(n_764),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3305),
.B(n_967),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3452),
.Y(n_3730)
);

INVx2_ASAP7_75t_SL g3731 ( 
.A(n_3268),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3202),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3329),
.B(n_764),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3519),
.B(n_3490),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3457),
.Y(n_3735)
);

AOI22xp33_ASAP7_75t_L g3736 ( 
.A1(n_3174),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.Y(n_3736)
);

BUFx3_ASAP7_75t_L g3737 ( 
.A(n_3450),
.Y(n_3737)
);

INVx4_ASAP7_75t_L g3738 ( 
.A(n_3362),
.Y(n_3738)
);

INVx3_ASAP7_75t_L g3739 ( 
.A(n_3470),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3507),
.B(n_766),
.Y(n_3740)
);

HB1xp67_ASAP7_75t_L g3741 ( 
.A(n_3317),
.Y(n_3741)
);

INVx3_ASAP7_75t_L g3742 ( 
.A(n_3470),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3387),
.B(n_769),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_3304),
.B(n_3474),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3373),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3484),
.B(n_770),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3373),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_3211),
.Y(n_3748)
);

BUFx6f_ASAP7_75t_L g3749 ( 
.A(n_3351),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3450),
.Y(n_3750)
);

INVx2_ASAP7_75t_SL g3751 ( 
.A(n_3405),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3174),
.B(n_770),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3364),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3364),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3446),
.Y(n_3755)
);

OAI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3444),
.A2(n_967),
.B(n_771),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3228),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3446),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3446),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3228),
.Y(n_3760)
);

INVx2_ASAP7_75t_SL g3761 ( 
.A(n_3352),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3288),
.B(n_964),
.Y(n_3762)
);

HB1xp67_ASAP7_75t_L g3763 ( 
.A(n_3309),
.Y(n_3763)
);

AOI22xp33_ASAP7_75t_L g3764 ( 
.A1(n_3210),
.A2(n_775),
.B1(n_772),
.B2(n_774),
.Y(n_3764)
);

HB1xp67_ASAP7_75t_L g3765 ( 
.A(n_3299),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3307),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3143),
.A2(n_776),
.B(n_777),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3284),
.Y(n_3768)
);

BUFx2_ASAP7_75t_SL g3769 ( 
.A(n_3386),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3416),
.B(n_778),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3284),
.Y(n_3771)
);

AND2x4_ASAP7_75t_L g3772 ( 
.A(n_3331),
.B(n_779),
.Y(n_3772)
);

AOI22xp33_ASAP7_75t_L g3773 ( 
.A1(n_3137),
.A2(n_782),
.B1(n_779),
.B2(n_780),
.Y(n_3773)
);

AO21x2_ASAP7_75t_L g3774 ( 
.A1(n_3346),
.A2(n_780),
.B(n_782),
.Y(n_3774)
);

AOI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3489),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3416),
.B(n_963),
.Y(n_3776)
);

AND2x4_ASAP7_75t_L g3777 ( 
.A(n_3331),
.B(n_783),
.Y(n_3777)
);

BUFx2_ASAP7_75t_L g3778 ( 
.A(n_3511),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_SL g3779 ( 
.A(n_3144),
.B(n_785),
.Y(n_3779)
);

INVx2_ASAP7_75t_SL g3780 ( 
.A(n_3299),
.Y(n_3780)
);

INVx3_ASAP7_75t_L g3781 ( 
.A(n_3511),
.Y(n_3781)
);

OR2x6_ASAP7_75t_L g3782 ( 
.A(n_3489),
.B(n_788),
.Y(n_3782)
);

AOI22xp33_ASAP7_75t_L g3783 ( 
.A1(n_3249),
.A2(n_790),
.B1(n_788),
.B2(n_789),
.Y(n_3783)
);

INVx3_ASAP7_75t_L g3784 ( 
.A(n_3511),
.Y(n_3784)
);

AND2x4_ASAP7_75t_SL g3785 ( 
.A(n_3216),
.B(n_790),
.Y(n_3785)
);

BUFx2_ASAP7_75t_L g3786 ( 
.A(n_3509),
.Y(n_3786)
);

INVx2_ASAP7_75t_SL g3787 ( 
.A(n_3509),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3310),
.B(n_791),
.Y(n_3788)
);

OAI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_3324),
.A2(n_791),
.B(n_792),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3408),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3408),
.Y(n_3791)
);

OR2x2_ASAP7_75t_L g3792 ( 
.A(n_3248),
.B(n_793),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3410),
.Y(n_3793)
);

OAI222xp33_ASAP7_75t_L g3794 ( 
.A1(n_3426),
.A2(n_793),
.B1(n_794),
.B2(n_795),
.C1(n_796),
.C2(n_797),
.Y(n_3794)
);

AND2x4_ASAP7_75t_SL g3795 ( 
.A(n_3486),
.B(n_794),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3410),
.Y(n_3796)
);

HB1xp67_ASAP7_75t_L g3797 ( 
.A(n_3486),
.Y(n_3797)
);

HB1xp67_ASAP7_75t_L g3798 ( 
.A(n_3496),
.Y(n_3798)
);

HB1xp67_ASAP7_75t_L g3799 ( 
.A(n_3496),
.Y(n_3799)
);

OR2x2_ASAP7_75t_L g3800 ( 
.A(n_3398),
.B(n_795),
.Y(n_3800)
);

BUFx3_ASAP7_75t_L g3801 ( 
.A(n_3520),
.Y(n_3801)
);

BUFx2_ASAP7_75t_L g3802 ( 
.A(n_3520),
.Y(n_3802)
);

NOR2x1_ASAP7_75t_SL g3803 ( 
.A(n_3209),
.B(n_796),
.Y(n_3803)
);

INVx3_ASAP7_75t_L g3804 ( 
.A(n_3285),
.Y(n_3804)
);

BUFx3_ASAP7_75t_L g3805 ( 
.A(n_3433),
.Y(n_3805)
);

AOI21x1_ASAP7_75t_L g3806 ( 
.A1(n_3213),
.A2(n_798),
.B(n_799),
.Y(n_3806)
);

INVx3_ASAP7_75t_L g3807 ( 
.A(n_3155),
.Y(n_3807)
);

INVx3_ASAP7_75t_L g3808 ( 
.A(n_3351),
.Y(n_3808)
);

AND2x4_ASAP7_75t_L g3809 ( 
.A(n_3413),
.B(n_799),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3166),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3431),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3461),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3461),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3286),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3293),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3255),
.B(n_800),
.Y(n_3816)
);

INVxp67_ASAP7_75t_SL g3817 ( 
.A(n_3351),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3166),
.Y(n_3818)
);

AO31x2_ASAP7_75t_L g3819 ( 
.A1(n_3427),
.A2(n_3374),
.A3(n_3378),
.B(n_3368),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3219),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3443),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3219),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3419),
.B(n_963),
.Y(n_3823)
);

BUFx6f_ASAP7_75t_L g3824 ( 
.A(n_3433),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3314),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3224),
.B(n_800),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3421),
.B(n_801),
.Y(n_3827)
);

INVx3_ASAP7_75t_L g3828 ( 
.A(n_3504),
.Y(n_3828)
);

OR2x2_ASAP7_75t_L g3829 ( 
.A(n_3417),
.B(n_801),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3443),
.Y(n_3830)
);

OAI22xp5_ASAP7_75t_L g3831 ( 
.A1(n_3258),
.A2(n_804),
.B1(n_802),
.B2(n_803),
.Y(n_3831)
);

OAI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_3347),
.A2(n_805),
.B1(n_802),
.B2(n_803),
.Y(n_3832)
);

AND2x4_ASAP7_75t_L g3833 ( 
.A(n_3413),
.B(n_3348),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_L g3834 ( 
.A(n_3506),
.B(n_805),
.Y(n_3834)
);

BUFx6f_ASAP7_75t_L g3835 ( 
.A(n_3500),
.Y(n_3835)
);

OAI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3301),
.A2(n_808),
.B(n_809),
.Y(n_3836)
);

INVx2_ASAP7_75t_SL g3837 ( 
.A(n_3437),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3318),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3445),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3445),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3454),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3504),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3361),
.A2(n_811),
.B1(n_808),
.B2(n_810),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3319),
.Y(n_3844)
);

OR2x2_ASAP7_75t_L g3845 ( 
.A(n_3455),
.B(n_810),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3476),
.B(n_812),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3274),
.B(n_813),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_3512),
.B(n_814),
.Y(n_3848)
);

INVx2_ASAP7_75t_SL g3849 ( 
.A(n_3451),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3188),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3315),
.B(n_962),
.Y(n_3851)
);

INVx1_ASAP7_75t_SL g3852 ( 
.A(n_3135),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3359),
.B(n_962),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3468),
.Y(n_3854)
);

AO31x2_ASAP7_75t_L g3855 ( 
.A1(n_3368),
.A2(n_818),
.A3(n_816),
.B(n_817),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3479),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3483),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3338),
.B(n_816),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3502),
.B(n_961),
.Y(n_3859)
);

INVx2_ASAP7_75t_SL g3860 ( 
.A(n_3500),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3473),
.B(n_817),
.Y(n_3861)
);

BUFx2_ASAP7_75t_L g3862 ( 
.A(n_3381),
.Y(n_3862)
);

INVxp67_ASAP7_75t_L g3863 ( 
.A(n_3139),
.Y(n_3863)
);

BUFx2_ASAP7_75t_L g3864 ( 
.A(n_3381),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_L g3865 ( 
.A(n_3559),
.B(n_3242),
.Y(n_3865)
);

AND2x4_ASAP7_75t_L g3866 ( 
.A(n_3558),
.B(n_3348),
.Y(n_3866)
);

NAND2xp33_ASAP7_75t_R g3867 ( 
.A(n_3669),
.B(n_3389),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3567),
.B(n_3456),
.Y(n_3868)
);

INVxp67_ASAP7_75t_L g3869 ( 
.A(n_3691),
.Y(n_3869)
);

BUFx3_ASAP7_75t_L g3870 ( 
.A(n_3534),
.Y(n_3870)
);

NAND2xp33_ASAP7_75t_R g3871 ( 
.A(n_3669),
.B(n_3389),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3684),
.B(n_3456),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3572),
.B(n_3577),
.Y(n_3873)
);

CKINVDCx5p33_ASAP7_75t_R g3874 ( 
.A(n_3626),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3587),
.B(n_3374),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3528),
.Y(n_3876)
);

OR2x6_ASAP7_75t_L g3877 ( 
.A(n_3738),
.B(n_3313),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3555),
.Y(n_3878)
);

NAND2xp33_ASAP7_75t_R g3879 ( 
.A(n_3782),
.B(n_3491),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3590),
.B(n_3378),
.Y(n_3880)
);

INVx8_ASAP7_75t_L g3881 ( 
.A(n_3543),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3537),
.B(n_3363),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3562),
.B(n_3340),
.Y(n_3883)
);

BUFx3_ASAP7_75t_L g3884 ( 
.A(n_3679),
.Y(n_3884)
);

CKINVDCx5p33_ASAP7_75t_R g3885 ( 
.A(n_3547),
.Y(n_3885)
);

NAND2xp33_ASAP7_75t_R g3886 ( 
.A(n_3782),
.B(n_3491),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3564),
.B(n_3341),
.Y(n_3887)
);

OR2x2_ASAP7_75t_L g3888 ( 
.A(n_3560),
.B(n_3379),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_R g3889 ( 
.A(n_3540),
.B(n_3327),
.Y(n_3889)
);

INVxp67_ASAP7_75t_L g3890 ( 
.A(n_3609),
.Y(n_3890)
);

NAND2xp33_ASAP7_75t_R g3891 ( 
.A(n_3539),
.B(n_3522),
.Y(n_3891)
);

XNOR2xp5_ASAP7_75t_L g3892 ( 
.A(n_3748),
.B(n_3199),
.Y(n_3892)
);

XNOR2xp5_ASAP7_75t_L g3893 ( 
.A(n_3583),
.B(n_3584),
.Y(n_3893)
);

BUFx3_ASAP7_75t_L g3894 ( 
.A(n_3714),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3660),
.B(n_3366),
.Y(n_3895)
);

OR2x6_ASAP7_75t_L g3896 ( 
.A(n_3738),
.B(n_3245),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_R g3897 ( 
.A(n_3706),
.B(n_818),
.Y(n_3897)
);

NOR2xp33_ASAP7_75t_R g3898 ( 
.A(n_3706),
.B(n_820),
.Y(n_3898)
);

BUFx24_ASAP7_75t_SL g3899 ( 
.A(n_3597),
.Y(n_3899)
);

OR2x6_ASAP7_75t_L g3900 ( 
.A(n_3665),
.B(n_3593),
.Y(n_3900)
);

NAND2xp33_ASAP7_75t_R g3901 ( 
.A(n_3539),
.B(n_3522),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3563),
.Y(n_3902)
);

OR2x2_ASAP7_75t_L g3903 ( 
.A(n_3566),
.B(n_3363),
.Y(n_3903)
);

AND2x4_ASAP7_75t_L g3904 ( 
.A(n_3660),
.B(n_3423),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3573),
.B(n_3182),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_R g3906 ( 
.A(n_3624),
.B(n_821),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3536),
.Y(n_3907)
);

AND2x4_ASAP7_75t_L g3908 ( 
.A(n_3709),
.B(n_3423),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3634),
.B(n_3161),
.Y(n_3909)
);

OR2x2_ASAP7_75t_L g3910 ( 
.A(n_3599),
.B(n_3239),
.Y(n_3910)
);

HB1xp67_ASAP7_75t_L g3911 ( 
.A(n_3763),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3561),
.B(n_3223),
.Y(n_3912)
);

NOR2xp33_ASAP7_75t_R g3913 ( 
.A(n_3605),
.B(n_822),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3639),
.B(n_3650),
.Y(n_3914)
);

XNOR2xp5_ASAP7_75t_L g3915 ( 
.A(n_3659),
.B(n_3326),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3576),
.B(n_3235),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3682),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3596),
.B(n_3198),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3721),
.B(n_3198),
.Y(n_3919)
);

NAND2xp33_ASAP7_75t_SL g3920 ( 
.A(n_3709),
.B(n_3328),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3741),
.B(n_3198),
.Y(n_3921)
);

AND2x4_ASAP7_75t_L g3922 ( 
.A(n_3579),
.B(n_3342),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_R g3923 ( 
.A(n_3579),
.B(n_823),
.Y(n_3923)
);

NAND2xp33_ASAP7_75t_R g3924 ( 
.A(n_3715),
.B(n_3428),
.Y(n_3924)
);

OR2x4_ASAP7_75t_L g3925 ( 
.A(n_3744),
.B(n_3336),
.Y(n_3925)
);

BUFx10_ASAP7_75t_L g3926 ( 
.A(n_3593),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3809),
.B(n_3308),
.Y(n_3927)
);

NAND2xp33_ASAP7_75t_R g3928 ( 
.A(n_3770),
.B(n_3428),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3809),
.B(n_3308),
.Y(n_3929)
);

INVxp67_ASAP7_75t_L g3930 ( 
.A(n_3531),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_R g3931 ( 
.A(n_3638),
.B(n_826),
.Y(n_3931)
);

INVxp67_ASAP7_75t_L g3932 ( 
.A(n_3705),
.Y(n_3932)
);

XNOR2xp5_ASAP7_75t_L g3933 ( 
.A(n_3657),
.B(n_3426),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_SL g3934 ( 
.A(n_3643),
.B(n_3330),
.Y(n_3934)
);

CKINVDCx8_ASAP7_75t_R g3935 ( 
.A(n_3769),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3538),
.Y(n_3936)
);

CKINVDCx14_ASAP7_75t_R g3937 ( 
.A(n_3686),
.Y(n_3937)
);

AND2x4_ASAP7_75t_L g3938 ( 
.A(n_3530),
.B(n_3342),
.Y(n_3938)
);

INVxp67_ASAP7_75t_L g3939 ( 
.A(n_3526),
.Y(n_3939)
);

NAND2xp33_ASAP7_75t_R g3940 ( 
.A(n_3776),
.B(n_3240),
.Y(n_3940)
);

BUFx10_ASAP7_75t_L g3941 ( 
.A(n_3523),
.Y(n_3941)
);

NOR2xp33_ASAP7_75t_L g3942 ( 
.A(n_3595),
.B(n_3283),
.Y(n_3942)
);

XNOR2xp5_ASAP7_75t_L g3943 ( 
.A(n_3637),
.B(n_3173),
.Y(n_3943)
);

AND2x4_ASAP7_75t_L g3944 ( 
.A(n_3610),
.B(n_3302),
.Y(n_3944)
);

CKINVDCx20_ASAP7_75t_R g3945 ( 
.A(n_3714),
.Y(n_3945)
);

BUFx3_ASAP7_75t_L g3946 ( 
.A(n_3523),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3683),
.Y(n_3947)
);

NOR2xp33_ASAP7_75t_R g3948 ( 
.A(n_3673),
.B(n_826),
.Y(n_3948)
);

NAND2xp33_ASAP7_75t_R g3949 ( 
.A(n_3718),
.B(n_3240),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3546),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3553),
.Y(n_3951)
);

BUFx10_ASAP7_75t_L g3952 ( 
.A(n_3523),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3644),
.B(n_3615),
.Y(n_3953)
);

INVxp67_ASAP7_75t_L g3954 ( 
.A(n_3681),
.Y(n_3954)
);

NAND2xp33_ASAP7_75t_R g3955 ( 
.A(n_3729),
.B(n_3154),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3551),
.Y(n_3956)
);

NAND2xp33_ASAP7_75t_R g3957 ( 
.A(n_3752),
.B(n_3643),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3594),
.Y(n_3958)
);

XNOR2xp5_ASAP7_75t_L g3959 ( 
.A(n_3604),
.B(n_3333),
.Y(n_3959)
);

XNOR2xp5_ASAP7_75t_L g3960 ( 
.A(n_3656),
.B(n_3203),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3603),
.Y(n_3961)
);

CKINVDCx5p33_ASAP7_75t_R g3962 ( 
.A(n_3697),
.Y(n_3962)
);

INVx8_ASAP7_75t_L g3963 ( 
.A(n_3529),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3670),
.B(n_3208),
.Y(n_3964)
);

XOR2xp5_ASAP7_75t_L g3965 ( 
.A(n_3734),
.B(n_3316),
.Y(n_3965)
);

NOR2xp33_ASAP7_75t_R g3966 ( 
.A(n_3673),
.B(n_3731),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_R g3967 ( 
.A(n_3529),
.B(n_3533),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3571),
.Y(n_3968)
);

NOR2xp33_ASAP7_75t_R g3969 ( 
.A(n_3529),
.B(n_827),
.Y(n_3969)
);

NAND2xp33_ASAP7_75t_R g3970 ( 
.A(n_3678),
.B(n_3710),
.Y(n_3970)
);

NOR2xp33_ASAP7_75t_R g3971 ( 
.A(n_3533),
.B(n_3668),
.Y(n_3971)
);

NOR2xp33_ASAP7_75t_R g3972 ( 
.A(n_3533),
.B(n_827),
.Y(n_3972)
);

INVxp67_ASAP7_75t_L g3973 ( 
.A(n_3642),
.Y(n_3973)
);

NOR2xp33_ASAP7_75t_R g3974 ( 
.A(n_3668),
.B(n_3745),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3671),
.B(n_3236),
.Y(n_3975)
);

INVxp67_ASAP7_75t_L g3976 ( 
.A(n_3630),
.Y(n_3976)
);

NOR2xp33_ASAP7_75t_R g3977 ( 
.A(n_3747),
.B(n_828),
.Y(n_3977)
);

BUFx2_ASAP7_75t_L g3978 ( 
.A(n_3739),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_3678),
.B(n_3237),
.Y(n_3979)
);

BUFx3_ASAP7_75t_L g3980 ( 
.A(n_3649),
.Y(n_3980)
);

NOR2xp33_ASAP7_75t_R g3981 ( 
.A(n_3753),
.B(n_828),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3598),
.B(n_3308),
.Y(n_3982)
);

NOR2xp33_ASAP7_75t_R g3983 ( 
.A(n_3754),
.B(n_829),
.Y(n_3983)
);

NAND2xp33_ASAP7_75t_R g3984 ( 
.A(n_3710),
.B(n_3154),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3632),
.B(n_3251),
.Y(n_3985)
);

CKINVDCx5p33_ASAP7_75t_R g3986 ( 
.A(n_3699),
.Y(n_3986)
);

NAND2xp33_ASAP7_75t_R g3987 ( 
.A(n_3733),
.B(n_830),
.Y(n_3987)
);

AND2x4_ASAP7_75t_L g3988 ( 
.A(n_3713),
.B(n_3291),
.Y(n_3988)
);

NAND2xp33_ASAP7_75t_R g3989 ( 
.A(n_3733),
.B(n_832),
.Y(n_3989)
);

NAND2xp33_ASAP7_75t_R g3990 ( 
.A(n_3772),
.B(n_3777),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_R g3991 ( 
.A(n_3751),
.B(n_833),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3633),
.B(n_3480),
.Y(n_3992)
);

AND2x4_ASAP7_75t_L g3993 ( 
.A(n_3713),
.B(n_3296),
.Y(n_3993)
);

NAND2xp33_ASAP7_75t_R g3994 ( 
.A(n_3772),
.B(n_833),
.Y(n_3994)
);

BUFx10_ASAP7_75t_L g3995 ( 
.A(n_3649),
.Y(n_3995)
);

AND2x4_ASAP7_75t_L g3996 ( 
.A(n_3722),
.B(n_3271),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3722),
.B(n_3168),
.Y(n_3997)
);

AND2x4_ASAP7_75t_L g3998 ( 
.A(n_3833),
.B(n_3739),
.Y(n_3998)
);

OR2x6_ASAP7_75t_L g3999 ( 
.A(n_3565),
.B(n_3311),
.Y(n_3999)
);

OR2x6_ASAP7_75t_L g4000 ( 
.A(n_3565),
.B(n_3438),
.Y(n_4000)
);

BUFx3_ASAP7_75t_L g4001 ( 
.A(n_3649),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3833),
.B(n_3294),
.Y(n_4002)
);

INVx8_ASAP7_75t_L g4003 ( 
.A(n_3692),
.Y(n_4003)
);

INVxp67_ASAP7_75t_L g4004 ( 
.A(n_3541),
.Y(n_4004)
);

HB1xp67_ASAP7_75t_L g4005 ( 
.A(n_3742),
.Y(n_4005)
);

AND2x4_ASAP7_75t_L g4006 ( 
.A(n_3742),
.B(n_3197),
.Y(n_4006)
);

AND2x4_ASAP7_75t_L g4007 ( 
.A(n_3616),
.B(n_3253),
.Y(n_4007)
);

AND2x4_ASAP7_75t_L g4008 ( 
.A(n_3606),
.B(n_3272),
.Y(n_4008)
);

NOR2xp33_ASAP7_75t_R g4009 ( 
.A(n_3761),
.B(n_834),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3622),
.B(n_3442),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3693),
.Y(n_4011)
);

AND2x4_ASAP7_75t_L g4012 ( 
.A(n_3606),
.B(n_3335),
.Y(n_4012)
);

AND2x4_ASAP7_75t_L g4013 ( 
.A(n_3611),
.B(n_3337),
.Y(n_4013)
);

AND2x4_ASAP7_75t_L g4014 ( 
.A(n_3611),
.B(n_3499),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_R g4015 ( 
.A(n_3692),
.B(n_835),
.Y(n_4015)
);

NOR2xp33_ASAP7_75t_R g4016 ( 
.A(n_3692),
.B(n_836),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3812),
.B(n_3294),
.Y(n_4017)
);

INVx2_ASAP7_75t_SL g4018 ( 
.A(n_3701),
.Y(n_4018)
);

AND2x4_ASAP7_75t_L g4019 ( 
.A(n_3631),
.B(n_3499),
.Y(n_4019)
);

CKINVDCx20_ASAP7_75t_R g4020 ( 
.A(n_3737),
.Y(n_4020)
);

OR2x2_ASAP7_75t_L g4021 ( 
.A(n_3554),
.B(n_3515),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3623),
.B(n_3448),
.Y(n_4022)
);

CKINVDCx5p33_ASAP7_75t_R g4023 ( 
.A(n_3852),
.Y(n_4023)
);

NAND2xp33_ASAP7_75t_R g4024 ( 
.A(n_3777),
.B(n_836),
.Y(n_4024)
);

OR2x6_ASAP7_75t_L g4025 ( 
.A(n_3863),
.B(n_3430),
.Y(n_4025)
);

XOR2xp5_ASAP7_75t_L g4026 ( 
.A(n_3542),
.B(n_3322),
.Y(n_4026)
);

NOR2xp33_ASAP7_75t_R g4027 ( 
.A(n_3701),
.B(n_837),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3627),
.B(n_3392),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3693),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3628),
.B(n_3375),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_R g4031 ( 
.A(n_3701),
.B(n_838),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3694),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3640),
.B(n_3217),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3641),
.B(n_3449),
.Y(n_4034)
);

XNOR2xp5_ASAP7_75t_L g4035 ( 
.A(n_3695),
.B(n_3514),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3694),
.Y(n_4036)
);

NOR2xp33_ASAP7_75t_R g4037 ( 
.A(n_3631),
.B(n_839),
.Y(n_4037)
);

NAND2xp33_ASAP7_75t_R g4038 ( 
.A(n_3662),
.B(n_840),
.Y(n_4038)
);

BUFx10_ASAP7_75t_L g4039 ( 
.A(n_3795),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3672),
.B(n_3388),
.Y(n_4040)
);

AND2x4_ASAP7_75t_L g4041 ( 
.A(n_3647),
.B(n_3503),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3647),
.B(n_3503),
.Y(n_4042)
);

BUFx3_ASAP7_75t_L g4043 ( 
.A(n_3750),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_3813),
.B(n_3222),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_R g4045 ( 
.A(n_3837),
.B(n_840),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3700),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3674),
.B(n_3675),
.Y(n_4047)
);

BUFx6f_ASAP7_75t_L g4048 ( 
.A(n_3749),
.Y(n_4048)
);

XNOR2xp5_ASAP7_75t_L g4049 ( 
.A(n_3702),
.B(n_3762),
.Y(n_4049)
);

XOR2xp5_ASAP7_75t_L g4050 ( 
.A(n_3800),
.B(n_3353),
.Y(n_4050)
);

INVxp67_ASAP7_75t_L g4051 ( 
.A(n_3619),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3680),
.B(n_3397),
.Y(n_4052)
);

AND2x4_ASAP7_75t_L g4053 ( 
.A(n_3651),
.B(n_3481),
.Y(n_4053)
);

NAND2xp33_ASAP7_75t_R g4054 ( 
.A(n_3662),
.B(n_841),
.Y(n_4054)
);

AND2x4_ASAP7_75t_L g4055 ( 
.A(n_3651),
.B(n_3481),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_R g4056 ( 
.A(n_3849),
.B(n_842),
.Y(n_4056)
);

BUFx8_ASAP7_75t_SL g4057 ( 
.A(n_3602),
.Y(n_4057)
);

BUFx3_ASAP7_75t_L g4058 ( 
.A(n_3801),
.Y(n_4058)
);

NAND2xp33_ASAP7_75t_R g4059 ( 
.A(n_3664),
.B(n_843),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_R g4060 ( 
.A(n_3664),
.B(n_843),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3581),
.B(n_3146),
.Y(n_4061)
);

BUFx3_ASAP7_75t_L g4062 ( 
.A(n_3805),
.Y(n_4062)
);

NOR2xp33_ASAP7_75t_R g4063 ( 
.A(n_3804),
.B(n_845),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_R g4064 ( 
.A(n_3804),
.B(n_845),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3588),
.B(n_3439),
.Y(n_4065)
);

NAND2xp33_ASAP7_75t_SL g4066 ( 
.A(n_3861),
.B(n_3441),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_3582),
.B(n_3447),
.Y(n_4067)
);

INVxp67_ASAP7_75t_L g4068 ( 
.A(n_3689),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3585),
.B(n_3146),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3700),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3589),
.B(n_3497),
.Y(n_4071)
);

NAND2xp33_ASAP7_75t_R g4072 ( 
.A(n_3847),
.B(n_3823),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3712),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_3629),
.B(n_3256),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_3527),
.B(n_3158),
.Y(n_4075)
);

NAND2xp33_ASAP7_75t_R g4076 ( 
.A(n_3788),
.B(n_846),
.Y(n_4076)
);

AND2x4_ASAP7_75t_L g4077 ( 
.A(n_3586),
.B(n_3312),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3712),
.Y(n_4078)
);

BUFx3_ASAP7_75t_L g4079 ( 
.A(n_3778),
.Y(n_4079)
);

BUFx12f_ASAP7_75t_L g4080 ( 
.A(n_3602),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3578),
.B(n_3177),
.Y(n_4081)
);

HB1xp67_ASAP7_75t_L g4082 ( 
.A(n_3765),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3607),
.Y(n_4083)
);

NAND2xp33_ASAP7_75t_R g4084 ( 
.A(n_3527),
.B(n_846),
.Y(n_4084)
);

NOR2xp33_ASAP7_75t_R g4085 ( 
.A(n_3704),
.B(n_847),
.Y(n_4085)
);

CKINVDCx16_ASAP7_75t_R g4086 ( 
.A(n_3740),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_R g4087 ( 
.A(n_3806),
.B(n_848),
.Y(n_4087)
);

BUFx10_ASAP7_75t_L g4088 ( 
.A(n_3785),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3716),
.Y(n_4089)
);

NAND2xp33_ASAP7_75t_R g4090 ( 
.A(n_3646),
.B(n_849),
.Y(n_4090)
);

AND2x4_ASAP7_75t_L g4091 ( 
.A(n_3636),
.B(n_3356),
.Y(n_4091)
);

NOR2xp33_ASAP7_75t_R g4092 ( 
.A(n_3781),
.B(n_3784),
.Y(n_4092)
);

CKINVDCx12_ASAP7_75t_R g4093 ( 
.A(n_3829),
.Y(n_4093)
);

INVxp67_ASAP7_75t_L g4094 ( 
.A(n_3703),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_R g4095 ( 
.A(n_3781),
.B(n_849),
.Y(n_4095)
);

NAND2xp33_ASAP7_75t_R g4096 ( 
.A(n_3646),
.B(n_850),
.Y(n_4096)
);

NAND2xp33_ASAP7_75t_R g4097 ( 
.A(n_3676),
.B(n_850),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3846),
.B(n_3290),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3746),
.B(n_3267),
.Y(n_4099)
);

NAND2xp33_ASAP7_75t_R g4100 ( 
.A(n_3676),
.B(n_851),
.Y(n_4100)
);

OR2x6_ASAP7_75t_L g4101 ( 
.A(n_3779),
.B(n_3160),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_3797),
.B(n_3140),
.Y(n_4102)
);

NOR2xp33_ASAP7_75t_R g4103 ( 
.A(n_3784),
.B(n_851),
.Y(n_4103)
);

AND2x4_ASAP7_75t_L g4104 ( 
.A(n_3636),
.B(n_3521),
.Y(n_4104)
);

BUFx10_ASAP7_75t_L g4105 ( 
.A(n_3848),
.Y(n_4105)
);

NAND2xp33_ASAP7_75t_R g4106 ( 
.A(n_3827),
.B(n_852),
.Y(n_4106)
);

NOR2xp33_ASAP7_75t_L g4107 ( 
.A(n_3845),
.B(n_853),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3716),
.Y(n_4108)
);

NAND2xp33_ASAP7_75t_R g4109 ( 
.A(n_3834),
.B(n_855),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3792),
.B(n_3666),
.Y(n_4110)
);

CKINVDCx5p33_ASAP7_75t_R g4111 ( 
.A(n_3859),
.Y(n_4111)
);

NOR2xp33_ASAP7_75t_R g4112 ( 
.A(n_3808),
.B(n_855),
.Y(n_4112)
);

AND2x4_ASAP7_75t_L g4113 ( 
.A(n_3568),
.B(n_3517),
.Y(n_4113)
);

NAND2xp33_ASAP7_75t_R g4114 ( 
.A(n_3853),
.B(n_857),
.Y(n_4114)
);

OR2x6_ASAP7_75t_L g4115 ( 
.A(n_3654),
.B(n_3767),
.Y(n_4115)
);

OR2x6_ASAP7_75t_L g4116 ( 
.A(n_3677),
.B(n_3234),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_3743),
.B(n_3195),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_3621),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_3798),
.B(n_3232),
.Y(n_4119)
);

AND2x4_ASAP7_75t_L g4120 ( 
.A(n_3568),
.B(n_3493),
.Y(n_4120)
);

NAND2xp33_ASAP7_75t_R g4121 ( 
.A(n_3786),
.B(n_857),
.Y(n_4121)
);

BUFx3_ASAP7_75t_L g4122 ( 
.A(n_3802),
.Y(n_4122)
);

OR2x6_ASAP7_75t_L g4123 ( 
.A(n_3756),
.B(n_3422),
.Y(n_4123)
);

BUFx3_ASAP7_75t_L g4124 ( 
.A(n_3824),
.Y(n_4124)
);

NAND2xp33_ASAP7_75t_R g4125 ( 
.A(n_3858),
.B(n_858),
.Y(n_4125)
);

AND2x4_ASAP7_75t_L g4126 ( 
.A(n_3780),
.B(n_3495),
.Y(n_4126)
);

INVxp67_ASAP7_75t_L g4127 ( 
.A(n_3592),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3524),
.B(n_3355),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_3799),
.B(n_3232),
.Y(n_4129)
);

AND2x4_ASAP7_75t_L g4130 ( 
.A(n_3787),
.B(n_3395),
.Y(n_4130)
);

INVxp67_ASAP7_75t_L g4131 ( 
.A(n_3826),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_3860),
.B(n_3400),
.Y(n_4132)
);

INVxp67_ASAP7_75t_L g4133 ( 
.A(n_3803),
.Y(n_4133)
);

NAND2xp33_ASAP7_75t_R g4134 ( 
.A(n_3828),
.B(n_858),
.Y(n_4134)
);

AND2x4_ASAP7_75t_L g4135 ( 
.A(n_3817),
.B(n_3194),
.Y(n_4135)
);

NAND2xp33_ASAP7_75t_R g4136 ( 
.A(n_3828),
.B(n_859),
.Y(n_4136)
);

NOR2xp33_ASAP7_75t_R g4137 ( 
.A(n_3808),
.B(n_3736),
.Y(n_4137)
);

CKINVDCx11_ASAP7_75t_R g4138 ( 
.A(n_3945),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3911),
.Y(n_4139)
);

OAI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_4123),
.A2(n_3775),
.B1(n_3764),
.B2(n_3773),
.Y(n_4140)
);

INVxp67_ASAP7_75t_L g4141 ( 
.A(n_3870),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_3953),
.B(n_3569),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3978),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_3882),
.B(n_3569),
.Y(n_4144)
);

OAI22xp5_ASAP7_75t_L g4145 ( 
.A1(n_4123),
.A2(n_3836),
.B1(n_3783),
.B2(n_3732),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3918),
.B(n_3696),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3873),
.Y(n_4147)
);

OAI222xp33_ASAP7_75t_L g4148 ( 
.A1(n_3999),
.A2(n_3842),
.B1(n_3730),
.B2(n_3759),
.C1(n_3758),
.C2(n_3755),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3968),
.B(n_3601),
.Y(n_4149)
);

OR2x2_ASAP7_75t_L g4150 ( 
.A(n_3869),
.B(n_3524),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3917),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3947),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3880),
.B(n_3902),
.Y(n_4153)
);

AND2x2_ASAP7_75t_L g4154 ( 
.A(n_3875),
.B(n_3708),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3950),
.Y(n_4155)
);

INVxp67_ASAP7_75t_SL g4156 ( 
.A(n_4005),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3956),
.Y(n_4157)
);

INVxp67_ASAP7_75t_SL g4158 ( 
.A(n_4082),
.Y(n_4158)
);

BUFx2_ASAP7_75t_L g4159 ( 
.A(n_3966),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_3973),
.B(n_3711),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4122),
.B(n_3720),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4011),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3958),
.Y(n_4163)
);

INVxp67_ASAP7_75t_SL g4164 ( 
.A(n_3867),
.Y(n_4164)
);

BUFx3_ASAP7_75t_L g4165 ( 
.A(n_3884),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_SL g4166 ( 
.A(n_3948),
.B(n_3824),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3961),
.Y(n_4167)
);

INVx2_ASAP7_75t_SL g4168 ( 
.A(n_3894),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4029),
.Y(n_4169)
);

INVxp67_ASAP7_75t_SL g4170 ( 
.A(n_3871),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4032),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_3865),
.A2(n_3600),
.B1(n_3514),
.B2(n_3687),
.Y(n_4172)
);

HB1xp67_ASAP7_75t_L g4173 ( 
.A(n_3976),
.Y(n_4173)
);

NOR2xp33_ASAP7_75t_L g4174 ( 
.A(n_3937),
.B(n_3707),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4036),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_3998),
.B(n_3725),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4046),
.Y(n_4177)
);

NOR2x1_ASAP7_75t_SL g4178 ( 
.A(n_3900),
.B(n_3645),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_3866),
.B(n_3726),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3932),
.B(n_3525),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4070),
.Y(n_4181)
);

CKINVDCx20_ASAP7_75t_R g4182 ( 
.A(n_4020),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3982),
.B(n_3525),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4073),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_SL g4185 ( 
.A(n_4057),
.B(n_3794),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3919),
.B(n_3921),
.Y(n_4186)
);

HB1xp67_ASAP7_75t_L g4187 ( 
.A(n_4079),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3916),
.B(n_3532),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_3939),
.B(n_3532),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4078),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4089),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4108),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3914),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4083),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_4118),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3876),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4002),
.B(n_3535),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_3907),
.Y(n_4198)
);

AND2x2_ASAP7_75t_L g4199 ( 
.A(n_3910),
.B(n_3535),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4028),
.B(n_3608),
.Y(n_4200)
);

INVx1_ASAP7_75t_SL g4201 ( 
.A(n_4058),
.Y(n_4201)
);

INVx2_ASAP7_75t_SL g4202 ( 
.A(n_4003),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_4102),
.B(n_3544),
.Y(n_4203)
);

HB1xp67_ASAP7_75t_L g4204 ( 
.A(n_3878),
.Y(n_4204)
);

NAND3xp33_ASAP7_75t_L g4205 ( 
.A(n_3987),
.B(n_3728),
.C(n_3635),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_4000),
.A2(n_3648),
.B1(n_3259),
.B2(n_3570),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_3936),
.Y(n_4207)
);

BUFx2_ASAP7_75t_L g4208 ( 
.A(n_3971),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3912),
.B(n_3544),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_4000),
.A2(n_3259),
.B1(n_3667),
.B2(n_3789),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3930),
.B(n_3548),
.Y(n_4211)
);

BUFx2_ASAP7_75t_L g4212 ( 
.A(n_3967),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3868),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4051),
.B(n_3548),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_L g4215 ( 
.A(n_4086),
.B(n_860),
.Y(n_4215)
);

OR2x2_ASAP7_75t_L g4216 ( 
.A(n_3903),
.B(n_3549),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3927),
.B(n_3549),
.Y(n_4217)
);

INVx1_ASAP7_75t_SL g4218 ( 
.A(n_4062),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3872),
.Y(n_4219)
);

INVxp67_ASAP7_75t_SL g4220 ( 
.A(n_3879),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3951),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4047),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4017),
.Y(n_4223)
);

INVx1_ASAP7_75t_SL g4224 ( 
.A(n_4092),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3888),
.Y(n_4225)
);

OAI222xp33_ASAP7_75t_L g4226 ( 
.A1(n_3999),
.A2(n_3856),
.B1(n_3857),
.B2(n_3854),
.C1(n_3620),
.C2(n_3613),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4119),
.Y(n_4227)
);

AND2x2_ASAP7_75t_L g4228 ( 
.A(n_4129),
.B(n_3550),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3929),
.B(n_3550),
.Y(n_4229)
);

AOI22xp33_ASAP7_75t_L g4230 ( 
.A1(n_4080),
.A2(n_3774),
.B1(n_3851),
.B2(n_3371),
.Y(n_4230)
);

INVxp67_ASAP7_75t_SL g4231 ( 
.A(n_3886),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4074),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4067),
.B(n_3552),
.Y(n_4233)
);

OAI22xp5_ASAP7_75t_L g4234 ( 
.A1(n_3934),
.A2(n_3843),
.B1(n_3698),
.B2(n_3345),
.Y(n_4234)
);

INVx3_ASAP7_75t_L g4235 ( 
.A(n_3900),
.Y(n_4235)
);

OAI222xp33_ASAP7_75t_L g4236 ( 
.A1(n_3896),
.A2(n_3617),
.B1(n_3612),
.B2(n_3717),
.C1(n_3719),
.C2(n_3685),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_3904),
.B(n_3552),
.Y(n_4237)
);

AND2x4_ASAP7_75t_L g4238 ( 
.A(n_3908),
.B(n_3557),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_SL g4239 ( 
.A(n_3923),
.B(n_4037),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4061),
.B(n_3557),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3997),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4069),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4034),
.Y(n_4243)
);

OR2x2_ASAP7_75t_L g4244 ( 
.A(n_4021),
.B(n_3652),
.Y(n_4244)
);

OR2x2_ASAP7_75t_L g4245 ( 
.A(n_3890),
.B(n_3652),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_3954),
.B(n_3653),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4040),
.Y(n_4247)
);

CKINVDCx6p67_ASAP7_75t_R g4248 ( 
.A(n_3881),
.Y(n_4248)
);

AOI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_3989),
.A2(n_3831),
.B1(n_3832),
.B2(n_3343),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4052),
.Y(n_4250)
);

INVx1_ASAP7_75t_SL g4251 ( 
.A(n_3980),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4065),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4094),
.B(n_3653),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4071),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3992),
.Y(n_4255)
);

OAI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_3979),
.A2(n_3380),
.B(n_3192),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4033),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4025),
.B(n_3655),
.Y(n_4258)
);

INVxp67_ASAP7_75t_L g4259 ( 
.A(n_3970),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4006),
.Y(n_4260)
);

AND2x4_ASAP7_75t_L g4261 ( 
.A(n_4091),
.B(n_3655),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4025),
.B(n_3658),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_4001),
.Y(n_4263)
);

AOI22xp33_ASAP7_75t_L g4264 ( 
.A1(n_3920),
.A2(n_3614),
.B1(n_3545),
.B2(n_3436),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4077),
.B(n_3658),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4004),
.B(n_3661),
.Y(n_4266)
);

NOR2xp33_ASAP7_75t_L g4267 ( 
.A(n_3925),
.B(n_860),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4162),
.Y(n_4268)
);

INVxp67_ASAP7_75t_SL g4269 ( 
.A(n_4156),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4142),
.B(n_4023),
.Y(n_4270)
);

AND2x2_ASAP7_75t_L g4271 ( 
.A(n_4144),
.B(n_3895),
.Y(n_4271)
);

INVx4_ASAP7_75t_L g4272 ( 
.A(n_4165),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4151),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4152),
.Y(n_4274)
);

INVx5_ASAP7_75t_L g4275 ( 
.A(n_4159),
.Y(n_4275)
);

OR2x2_ASAP7_75t_L g4276 ( 
.A(n_4186),
.B(n_3819),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4153),
.B(n_3986),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_4224),
.B(n_3906),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4257),
.B(n_4044),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4266),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_4164),
.B(n_4111),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4150),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_4255),
.B(n_4243),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4170),
.B(n_4008),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4204),
.Y(n_4285)
);

OR2x2_ASAP7_75t_L g4286 ( 
.A(n_4232),
.B(n_3819),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4220),
.B(n_4012),
.Y(n_4287)
);

INVxp67_ASAP7_75t_L g4288 ( 
.A(n_4187),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_4231),
.B(n_4007),
.Y(n_4289)
);

NAND3xp33_ASAP7_75t_L g4290 ( 
.A(n_4264),
.B(n_3955),
.C(n_3924),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_4225),
.B(n_3819),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4161),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4196),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_4158),
.B(n_4173),
.Y(n_4294)
);

OAI211xp5_ASAP7_75t_SL g4295 ( 
.A1(n_4239),
.A2(n_4131),
.B(n_4068),
.C(n_3935),
.Y(n_4295)
);

NAND3xp33_ASAP7_75t_L g4296 ( 
.A(n_4206),
.B(n_4185),
.C(n_4205),
.Y(n_4296)
);

BUFx2_ASAP7_75t_L g4297 ( 
.A(n_4208),
.Y(n_4297)
);

AND2x4_ASAP7_75t_SL g4298 ( 
.A(n_4248),
.B(n_4039),
.Y(n_4298)
);

AOI221xp5_ASAP7_75t_L g4299 ( 
.A1(n_4145),
.A2(n_4110),
.B1(n_4107),
.B2(n_4026),
.C(n_3965),
.Y(n_4299)
);

AOI221xp5_ASAP7_75t_L g4300 ( 
.A1(n_4145),
.A2(n_3942),
.B1(n_4050),
.B2(n_3931),
.C(n_4066),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4169),
.Y(n_4301)
);

HB1xp67_ASAP7_75t_L g4302 ( 
.A(n_4201),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4179),
.B(n_4088),
.Y(n_4303)
);

NOR2xp33_ASAP7_75t_L g4304 ( 
.A(n_4168),
.B(n_3962),
.Y(n_4304)
);

NOR3xp33_ASAP7_75t_L g4305 ( 
.A(n_4205),
.B(n_4117),
.C(n_4133),
.Y(n_4305)
);

INVxp67_ASAP7_75t_L g4306 ( 
.A(n_4267),
.Y(n_4306)
);

AND2x4_ASAP7_75t_L g4307 ( 
.A(n_4258),
.B(n_4013),
.Y(n_4307)
);

INVx5_ASAP7_75t_SL g4308 ( 
.A(n_4138),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4197),
.B(n_3996),
.Y(n_4309)
);

AND2x2_ASAP7_75t_L g4310 ( 
.A(n_4253),
.B(n_4041),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4198),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4199),
.B(n_4042),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4171),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4245),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4160),
.B(n_4053),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_4207),
.Y(n_4316)
);

AND2x2_ASAP7_75t_L g4317 ( 
.A(n_4176),
.B(n_4055),
.Y(n_4317)
);

AND2x2_ASAP7_75t_L g4318 ( 
.A(n_4203),
.B(n_4014),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4139),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4221),
.Y(n_4320)
);

AOI221xp5_ASAP7_75t_L g4321 ( 
.A1(n_4234),
.A2(n_4099),
.B1(n_3913),
.B2(n_3933),
.C(n_4075),
.Y(n_4321)
);

INVx1_ASAP7_75t_SL g4322 ( 
.A(n_4201),
.Y(n_4322)
);

AOI33xp33_ASAP7_75t_L g4323 ( 
.A1(n_4247),
.A2(n_3899),
.A3(n_3372),
.B1(n_4072),
.B2(n_4125),
.B3(n_4114),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4180),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4155),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_4250),
.B(n_3661),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4157),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4244),
.Y(n_4328)
);

OAI211xp5_ASAP7_75t_L g4329 ( 
.A1(n_4259),
.A2(n_3897),
.B(n_3898),
.C(n_4045),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4163),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4154),
.B(n_4019),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_4224),
.A2(n_3896),
.B1(n_4218),
.B2(n_4166),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4167),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4175),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4177),
.Y(n_4335)
);

HB1xp67_ASAP7_75t_L g4336 ( 
.A(n_4218),
.Y(n_4336)
);

INVxp67_ASAP7_75t_SL g4337 ( 
.A(n_4143),
.Y(n_4337)
);

INVxp67_ASAP7_75t_L g4338 ( 
.A(n_4215),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_4252),
.B(n_3663),
.Y(n_4339)
);

NOR2xp33_ASAP7_75t_L g4340 ( 
.A(n_4141),
.B(n_3893),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4181),
.Y(n_4341)
);

BUFx2_ASAP7_75t_L g4342 ( 
.A(n_4212),
.Y(n_4342)
);

AND2x4_ASAP7_75t_L g4343 ( 
.A(n_4262),
.B(n_3988),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4189),
.B(n_3993),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_4254),
.B(n_4193),
.Y(n_4345)
);

NOR2xp33_ASAP7_75t_L g4346 ( 
.A(n_4182),
.B(n_3881),
.Y(n_4346)
);

OR2x2_ASAP7_75t_L g4347 ( 
.A(n_4188),
.B(n_3663),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4194),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4195),
.Y(n_4349)
);

OAI221xp5_ASAP7_75t_L g4350 ( 
.A1(n_4185),
.A2(n_4024),
.B1(n_3994),
.B2(n_4054),
.C(n_4038),
.Y(n_4350)
);

OAI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_4230),
.A2(n_3877),
.B1(n_4035),
.B2(n_4049),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4211),
.B(n_3974),
.Y(n_4352)
);

AOI33xp33_ASAP7_75t_L g4353 ( 
.A1(n_4214),
.A2(n_3458),
.A3(n_4121),
.B1(n_3407),
.B2(n_3944),
.B3(n_4109),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4184),
.Y(n_4354)
);

NAND2xp33_ASAP7_75t_SL g4355 ( 
.A(n_4235),
.B(n_3990),
.Y(n_4355)
);

AOI22xp5_ASAP7_75t_L g4356 ( 
.A1(n_4140),
.A2(n_4084),
.B1(n_4076),
.B2(n_3957),
.Y(n_4356)
);

OR2x2_ASAP7_75t_L g4357 ( 
.A(n_4209),
.B(n_3688),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4246),
.B(n_3723),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4190),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4191),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4147),
.B(n_3688),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4228),
.B(n_3724),
.Y(n_4362)
);

HB1xp67_ASAP7_75t_L g4363 ( 
.A(n_4227),
.Y(n_4363)
);

NAND3xp33_ASAP7_75t_L g4364 ( 
.A(n_4200),
.B(n_3940),
.C(n_3949),
.Y(n_4364)
);

AOI221xp5_ASAP7_75t_L g4365 ( 
.A1(n_4234),
.A2(n_3909),
.B1(n_3977),
.B2(n_3983),
.C(n_3981),
.Y(n_4365)
);

OR2x2_ASAP7_75t_L g4366 ( 
.A(n_4276),
.B(n_4242),
.Y(n_4366)
);

OR2x2_ASAP7_75t_L g4367 ( 
.A(n_4363),
.B(n_4223),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4271),
.B(n_4241),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4268),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4344),
.B(n_4315),
.Y(n_4370)
);

INVx3_ASAP7_75t_L g4371 ( 
.A(n_4272),
.Y(n_4371)
);

OR2x2_ASAP7_75t_L g4372 ( 
.A(n_4328),
.B(n_4217),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4280),
.B(n_4213),
.Y(n_4373)
);

NAND2x1_ASAP7_75t_L g4374 ( 
.A(n_4272),
.B(n_4235),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4285),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4268),
.Y(n_4376)
);

AND2x4_ASAP7_75t_L g4377 ( 
.A(n_4364),
.B(n_4261),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4342),
.Y(n_4378)
);

OR2x2_ASAP7_75t_L g4379 ( 
.A(n_4279),
.B(n_4229),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4309),
.B(n_4260),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4317),
.B(n_4289),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4301),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4301),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4291),
.B(n_4219),
.Y(n_4384)
);

INVx1_ASAP7_75t_SL g4385 ( 
.A(n_4322),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4297),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4313),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4331),
.B(n_4261),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4318),
.B(n_4237),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4313),
.Y(n_4390)
);

NAND2x1p5_ASAP7_75t_L g4391 ( 
.A(n_4275),
.B(n_4251),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4310),
.B(n_4237),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4359),
.Y(n_4393)
);

INVx2_ASAP7_75t_SL g4394 ( 
.A(n_4298),
.Y(n_4394)
);

OR2x2_ASAP7_75t_L g4395 ( 
.A(n_4269),
.B(n_4146),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4312),
.B(n_4238),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4359),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4282),
.B(n_4240),
.Y(n_4398)
);

AND2x4_ASAP7_75t_L g4399 ( 
.A(n_4275),
.B(n_4238),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4360),
.Y(n_4400)
);

AND2x4_ASAP7_75t_L g4401 ( 
.A(n_4275),
.B(n_4233),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4360),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4273),
.Y(n_4403)
);

INVx1_ASAP7_75t_SL g4404 ( 
.A(n_4302),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4343),
.B(n_4251),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4314),
.B(n_4222),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4343),
.B(n_4263),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4274),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4334),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_4284),
.B(n_4265),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4335),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4324),
.B(n_4362),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4341),
.Y(n_4413)
);

INVxp67_ASAP7_75t_L g4414 ( 
.A(n_4336),
.Y(n_4414)
);

AND2x4_ASAP7_75t_L g4415 ( 
.A(n_4307),
.B(n_4216),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4293),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4358),
.B(n_4183),
.Y(n_4417)
);

AND2x4_ASAP7_75t_L g4418 ( 
.A(n_4307),
.B(n_4178),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4354),
.Y(n_4419)
);

OR2x2_ASAP7_75t_L g4420 ( 
.A(n_4292),
.B(n_4200),
.Y(n_4420)
);

BUFx2_ASAP7_75t_L g4421 ( 
.A(n_4355),
.Y(n_4421)
);

AND2x2_ASAP7_75t_L g4422 ( 
.A(n_4287),
.B(n_4192),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4311),
.Y(n_4423)
);

NAND2x1_ASAP7_75t_L g4424 ( 
.A(n_4332),
.B(n_3877),
.Y(n_4424)
);

NAND2x1_ASAP7_75t_L g4425 ( 
.A(n_4352),
.B(n_3938),
.Y(n_4425)
);

OR2x2_ASAP7_75t_L g4426 ( 
.A(n_4347),
.B(n_4149),
.Y(n_4426)
);

OR2x2_ASAP7_75t_L g4427 ( 
.A(n_4357),
.B(n_4149),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4345),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4294),
.B(n_3727),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4325),
.Y(n_4430)
);

OAI221xp5_ASAP7_75t_SL g4431 ( 
.A1(n_4300),
.A2(n_4249),
.B1(n_4210),
.B2(n_3959),
.C(n_4172),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4327),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_4337),
.B(n_4174),
.Y(n_4433)
);

AOI221xp5_ASAP7_75t_L g4434 ( 
.A1(n_4296),
.A2(n_4140),
.B1(n_4256),
.B2(n_4148),
.C(n_4226),
.Y(n_4434)
);

AND2x2_ASAP7_75t_SL g4435 ( 
.A(n_4356),
.B(n_4281),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4303),
.B(n_4043),
.Y(n_4436)
);

OR2x2_ASAP7_75t_L g4437 ( 
.A(n_4283),
.B(n_3690),
.Y(n_4437)
);

INVxp67_ASAP7_75t_L g4438 ( 
.A(n_4278),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4326),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4339),
.Y(n_4440)
);

NAND2x1_ASAP7_75t_L g4441 ( 
.A(n_4290),
.B(n_3922),
.Y(n_4441)
);

OR2x2_ASAP7_75t_L g4442 ( 
.A(n_4286),
.B(n_3690),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4319),
.B(n_3618),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4305),
.B(n_3625),
.Y(n_4444)
);

NOR3xp33_ASAP7_75t_L g4445 ( 
.A(n_4350),
.B(n_4321),
.C(n_4351),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4434),
.B(n_4288),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4428),
.B(n_4323),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4439),
.B(n_4440),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4442),
.Y(n_4449)
);

AO221x2_ASAP7_75t_L g4450 ( 
.A1(n_4424),
.A2(n_4308),
.B1(n_4236),
.B2(n_4329),
.C(n_4365),
.Y(n_4450)
);

INVx4_ASAP7_75t_L g4451 ( 
.A(n_4371),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4384),
.B(n_4361),
.Y(n_4452)
);

OAI221xp5_ASAP7_75t_L g4453 ( 
.A1(n_4445),
.A2(n_4299),
.B1(n_4295),
.B2(n_4306),
.C(n_4338),
.Y(n_4453)
);

INVx1_ASAP7_75t_SL g4454 ( 
.A(n_4436),
.Y(n_4454)
);

OAI22xp33_ASAP7_75t_L g4455 ( 
.A1(n_4424),
.A2(n_3984),
.B1(n_4059),
.B2(n_3928),
.Y(n_4455)
);

AOI22xp5_ASAP7_75t_L g4456 ( 
.A1(n_4435),
.A2(n_4134),
.B1(n_4136),
.B2(n_4106),
.Y(n_4456)
);

OAI22xp33_ASAP7_75t_L g4457 ( 
.A1(n_4425),
.A2(n_3901),
.B1(n_3891),
.B2(n_4090),
.Y(n_4457)
);

AO221x2_ASAP7_75t_L g4458 ( 
.A1(n_4394),
.A2(n_4308),
.B1(n_4304),
.B2(n_4340),
.C(n_4277),
.Y(n_4458)
);

AO221x2_ASAP7_75t_L g4459 ( 
.A1(n_4378),
.A2(n_4093),
.B1(n_4056),
.B2(n_3991),
.C(n_4009),
.Y(n_4459)
);

NOR2xp33_ASAP7_75t_L g4460 ( 
.A(n_4438),
.B(n_4431),
.Y(n_4460)
);

AND2x4_ASAP7_75t_L g4461 ( 
.A(n_4386),
.B(n_4270),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_R g4462 ( 
.A(n_4385),
.B(n_3874),
.Y(n_4462)
);

NAND2xp33_ASAP7_75t_SL g4463 ( 
.A(n_4421),
.B(n_4060),
.Y(n_4463)
);

INVxp33_ASAP7_75t_SL g4464 ( 
.A(n_4404),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_4444),
.B(n_4316),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4414),
.B(n_4320),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4429),
.B(n_4330),
.Y(n_4467)
);

NOR2xp33_ASAP7_75t_L g4468 ( 
.A(n_4433),
.B(n_4346),
.Y(n_4468)
);

NAND2xp33_ASAP7_75t_SL g4469 ( 
.A(n_4374),
.B(n_4015),
.Y(n_4469)
);

OAI221xp5_ASAP7_75t_L g4470 ( 
.A1(n_4441),
.A2(n_4256),
.B1(n_4249),
.B2(n_3892),
.C(n_3915),
.Y(n_4470)
);

CKINVDCx8_ASAP7_75t_R g4471 ( 
.A(n_4399),
.Y(n_4471)
);

INVx2_ASAP7_75t_SL g4472 ( 
.A(n_4405),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4417),
.B(n_4333),
.Y(n_4473)
);

HB1xp67_ASAP7_75t_L g4474 ( 
.A(n_4367),
.Y(n_4474)
);

OAI22xp33_ASAP7_75t_L g4475 ( 
.A1(n_4425),
.A2(n_4096),
.B1(n_4100),
.B2(n_4097),
.Y(n_4475)
);

CKINVDCx5p33_ASAP7_75t_R g4476 ( 
.A(n_4381),
.Y(n_4476)
);

INVx3_ASAP7_75t_L g4477 ( 
.A(n_4399),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4416),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4375),
.B(n_4348),
.Y(n_4479)
);

NOR2xp33_ASAP7_75t_L g4480 ( 
.A(n_4406),
.B(n_4373),
.Y(n_4480)
);

INVxp33_ASAP7_75t_SL g4481 ( 
.A(n_4389),
.Y(n_4481)
);

NOR2xp33_ASAP7_75t_L g4482 ( 
.A(n_4370),
.B(n_3885),
.Y(n_4482)
);

AND2x4_ASAP7_75t_L g4483 ( 
.A(n_4415),
.B(n_4202),
.Y(n_4483)
);

AOI22xp5_ASAP7_75t_L g4484 ( 
.A1(n_4377),
.A2(n_3960),
.B1(n_3943),
.B2(n_4105),
.Y(n_4484)
);

OR2x2_ASAP7_75t_L g4485 ( 
.A(n_4426),
.B(n_4349),
.Y(n_4485)
);

OAI22xp33_ASAP7_75t_L g4486 ( 
.A1(n_4391),
.A2(n_4101),
.B1(n_4127),
.B2(n_4115),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_4366),
.B(n_4353),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_R g4488 ( 
.A(n_4418),
.B(n_3926),
.Y(n_4488)
);

AOI22xp5_ASAP7_75t_SL g4489 ( 
.A1(n_4418),
.A2(n_4064),
.B1(n_4063),
.B2(n_4016),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4377),
.B(n_4018),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4427),
.B(n_3625),
.Y(n_4491)
);

AO221x2_ASAP7_75t_L g4492 ( 
.A1(n_4412),
.A2(n_4031),
.B1(n_4027),
.B2(n_3889),
.C(n_4095),
.Y(n_4492)
);

NAND2xp33_ASAP7_75t_R g4493 ( 
.A(n_4401),
.B(n_3969),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4369),
.B(n_4104),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4423),
.Y(n_4495)
);

A2O1A1Ixp33_ASAP7_75t_L g4496 ( 
.A1(n_4415),
.A2(n_4003),
.B(n_3963),
.C(n_4098),
.Y(n_4496)
);

OAI22xp33_ASAP7_75t_L g4497 ( 
.A1(n_4395),
.A2(n_4101),
.B1(n_4115),
.B2(n_4116),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4376),
.B(n_4030),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4382),
.B(n_4113),
.Y(n_4499)
);

OAI22xp33_ASAP7_75t_L g4500 ( 
.A1(n_4401),
.A2(n_4116),
.B1(n_3862),
.B2(n_3864),
.Y(n_4500)
);

INVx2_ASAP7_75t_L g4501 ( 
.A(n_4474),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_4491),
.B(n_4420),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4448),
.Y(n_4503)
);

INVx3_ASAP7_75t_L g4504 ( 
.A(n_4458),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4473),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_4447),
.B(n_4383),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4477),
.B(n_4407),
.Y(n_4507)
);

AOI22xp33_ASAP7_75t_L g4508 ( 
.A1(n_4450),
.A2(n_4422),
.B1(n_4410),
.B2(n_4103),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4451),
.B(n_4388),
.Y(n_4509)
);

OR2x2_ASAP7_75t_L g4510 ( 
.A(n_4465),
.B(n_4379),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4449),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_4487),
.B(n_4372),
.Y(n_4512)
);

INVx1_ASAP7_75t_SL g4513 ( 
.A(n_4464),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4466),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4452),
.Y(n_4515)
);

OR2x2_ASAP7_75t_L g4516 ( 
.A(n_4485),
.B(n_4437),
.Y(n_4516)
);

INVxp67_ASAP7_75t_SL g4517 ( 
.A(n_4489),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4498),
.Y(n_4518)
);

AOI22xp33_ASAP7_75t_L g4519 ( 
.A1(n_4450),
.A2(n_4112),
.B1(n_3972),
.B2(n_4398),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4458),
.B(n_4392),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4467),
.Y(n_4521)
);

HB1xp67_ASAP7_75t_L g4522 ( 
.A(n_4478),
.Y(n_4522)
);

OR2x2_ASAP7_75t_L g4523 ( 
.A(n_4446),
.B(n_4443),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4479),
.Y(n_4524)
);

OR2x2_ASAP7_75t_L g4525 ( 
.A(n_4494),
.B(n_4387),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4499),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4472),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4460),
.B(n_4403),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4495),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4490),
.B(n_4396),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4480),
.B(n_4484),
.Y(n_4531)
);

NAND2x1_ASAP7_75t_SL g4532 ( 
.A(n_4456),
.B(n_4408),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4454),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4471),
.Y(n_4534)
);

AOI22xp33_ASAP7_75t_SL g4535 ( 
.A1(n_4459),
.A2(n_4409),
.B1(n_4413),
.B2(n_4411),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4475),
.B(n_4419),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4476),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4468),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4483),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4488),
.B(n_4368),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4461),
.Y(n_4541)
);

AND3x1_ASAP7_75t_L g4542 ( 
.A(n_4459),
.B(n_4432),
.C(n_4430),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4482),
.B(n_4380),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4496),
.B(n_4390),
.Y(n_4544)
);

INVx1_ASAP7_75t_SL g4545 ( 
.A(n_4462),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4463),
.Y(n_4546)
);

INVx1_ASAP7_75t_SL g4547 ( 
.A(n_4469),
.Y(n_4547)
);

INVxp67_ASAP7_75t_L g4548 ( 
.A(n_4453),
.Y(n_4548)
);

CKINVDCx5p33_ASAP7_75t_R g4549 ( 
.A(n_4493),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4492),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4481),
.Y(n_4551)
);

INVx1_ASAP7_75t_SL g4552 ( 
.A(n_4492),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4455),
.B(n_4402),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4470),
.Y(n_4554)
);

INVx3_ASAP7_75t_L g4555 ( 
.A(n_4457),
.Y(n_4555)
);

OAI21x1_ASAP7_75t_L g4556 ( 
.A1(n_4486),
.A2(n_4397),
.B(n_4393),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4497),
.B(n_4400),
.Y(n_4557)
);

AND2x4_ASAP7_75t_L g4558 ( 
.A(n_4500),
.B(n_4120),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4501),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4533),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4554),
.B(n_3855),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_4505),
.B(n_3855),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4524),
.Y(n_4563)
);

OAI22xp5_ASAP7_75t_L g4564 ( 
.A1(n_4519),
.A2(n_4081),
.B1(n_4010),
.B2(n_4022),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4510),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4534),
.B(n_3995),
.Y(n_4566)
);

INVx1_ASAP7_75t_SL g4567 ( 
.A(n_4545),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4521),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4503),
.B(n_4514),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4551),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4516),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4518),
.Y(n_4572)
);

OAI322xp33_ASAP7_75t_L g4573 ( 
.A1(n_4548),
.A2(n_3964),
.A3(n_3816),
.B1(n_3975),
.B2(n_3985),
.C1(n_3905),
.C2(n_3354),
.Y(n_4573)
);

AOI22xp5_ASAP7_75t_L g4574 ( 
.A1(n_4517),
.A2(n_4126),
.B1(n_3883),
.B2(n_3887),
.Y(n_4574)
);

NOR4xp25_ASAP7_75t_L g4575 ( 
.A(n_4552),
.B(n_3184),
.C(n_3229),
.D(n_3377),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4512),
.Y(n_4576)
);

NAND3xp33_ASAP7_75t_L g4577 ( 
.A(n_4555),
.B(n_3270),
.C(n_3591),
.Y(n_4577)
);

OR4x1_ASAP7_75t_L g4578 ( 
.A(n_4546),
.B(n_3580),
.C(n_3815),
.D(n_3814),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4520),
.B(n_3946),
.Y(n_4579)
);

AOI322xp5_ASAP7_75t_L g4580 ( 
.A1(n_4504),
.A2(n_4128),
.A3(n_3820),
.B1(n_3822),
.B2(n_3757),
.C1(n_3760),
.C2(n_4135),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4515),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4538),
.B(n_3855),
.Y(n_4582)
);

AOI332xp33_ASAP7_75t_L g4583 ( 
.A1(n_4504),
.A2(n_3790),
.A3(n_3841),
.B1(n_3840),
.B2(n_3839),
.B3(n_3830),
.C1(n_3821),
.C2(n_3811),
.Y(n_4583)
);

AOI21xp33_ASAP7_75t_SL g4584 ( 
.A1(n_4549),
.A2(n_861),
.B(n_862),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4526),
.B(n_4085),
.Y(n_4585)
);

NOR4xp25_ASAP7_75t_L g4586 ( 
.A(n_4552),
.B(n_3406),
.C(n_4087),
.D(n_3850),
.Y(n_4586)
);

OAI211xp5_ASAP7_75t_SL g4587 ( 
.A1(n_4508),
.A2(n_4555),
.B(n_4535),
.C(n_4547),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_4522),
.Y(n_4588)
);

OAI32xp33_ASAP7_75t_L g4589 ( 
.A1(n_4547),
.A2(n_3807),
.A3(n_4124),
.B1(n_3793),
.B2(n_3796),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4511),
.Y(n_4590)
);

AO22x1_ASAP7_75t_L g4591 ( 
.A1(n_4550),
.A2(n_4132),
.B1(n_4130),
.B2(n_3807),
.Y(n_4591)
);

NOR2x1_ASAP7_75t_L g4592 ( 
.A(n_4545),
.B(n_3411),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_SL g4593 ( 
.A(n_4542),
.B(n_3941),
.Y(n_4593)
);

NOR2xp33_ASAP7_75t_L g4594 ( 
.A(n_4513),
.B(n_861),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4527),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4525),
.Y(n_4596)
);

AOI22xp5_ASAP7_75t_L g4597 ( 
.A1(n_4587),
.A2(n_4542),
.B1(n_4513),
.B2(n_4528),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4576),
.B(n_4570),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_4565),
.B(n_4506),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4560),
.B(n_4536),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4571),
.Y(n_4601)
);

NAND2x1_ASAP7_75t_L g4602 ( 
.A(n_4588),
.B(n_4509),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_SL g4603 ( 
.A(n_4586),
.B(n_4537),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4561),
.B(n_4506),
.Y(n_4604)
);

HB1xp67_ASAP7_75t_L g4605 ( 
.A(n_4559),
.Y(n_4605)
);

OAI22xp5_ASAP7_75t_L g4606 ( 
.A1(n_4574),
.A2(n_4531),
.B1(n_4523),
.B2(n_4539),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4567),
.B(n_4596),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4595),
.B(n_4553),
.Y(n_4608)
);

INVx1_ASAP7_75t_SL g4609 ( 
.A(n_4566),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4563),
.B(n_4544),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4569),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4581),
.Y(n_4612)
);

AOI22xp33_ASAP7_75t_L g4613 ( 
.A1(n_4564),
.A2(n_4577),
.B1(n_4579),
.B2(n_4568),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4578),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4572),
.B(n_4529),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_SL g4616 ( 
.A(n_4593),
.B(n_4556),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4590),
.Y(n_4617)
);

BUFx6f_ASAP7_75t_L g4618 ( 
.A(n_4594),
.Y(n_4618)
);

OAI21xp33_ASAP7_75t_L g4619 ( 
.A1(n_4574),
.A2(n_4532),
.B(n_4557),
.Y(n_4619)
);

NOR2x1_ASAP7_75t_L g4620 ( 
.A(n_4585),
.B(n_4540),
.Y(n_4620)
);

NOR2xp33_ASAP7_75t_L g4621 ( 
.A(n_4573),
.B(n_4541),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4582),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_4580),
.B(n_4502),
.Y(n_4623)
);

NOR2xp33_ASAP7_75t_L g4624 ( 
.A(n_4584),
.B(n_4543),
.Y(n_4624)
);

AND2x2_ASAP7_75t_SL g4625 ( 
.A(n_4575),
.B(n_4558),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4601),
.B(n_4562),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4607),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4605),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4609),
.Y(n_4629)
);

CKINVDCx5p33_ASAP7_75t_R g4630 ( 
.A(n_4618),
.Y(n_4630)
);

INVx2_ASAP7_75t_SL g4631 ( 
.A(n_4602),
.Y(n_4631)
);

INVx1_ASAP7_75t_SL g4632 ( 
.A(n_4618),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4598),
.Y(n_4633)
);

CKINVDCx20_ASAP7_75t_R g4634 ( 
.A(n_4618),
.Y(n_4634)
);

CKINVDCx16_ASAP7_75t_R g4635 ( 
.A(n_4620),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4615),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4621),
.B(n_4592),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4599),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4614),
.Y(n_4639)
);

CKINVDCx20_ASAP7_75t_R g4640 ( 
.A(n_4603),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4612),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4617),
.Y(n_4642)
);

INVx1_ASAP7_75t_SL g4643 ( 
.A(n_4611),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4604),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4600),
.Y(n_4645)
);

HB1xp67_ASAP7_75t_SL g4646 ( 
.A(n_4625),
.Y(n_4646)
);

NOR2xp33_ASAP7_75t_L g4647 ( 
.A(n_4597),
.B(n_4589),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4622),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4608),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4610),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4606),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4623),
.Y(n_4652)
);

AND4x1_ASAP7_75t_L g4653 ( 
.A(n_4651),
.B(n_4624),
.C(n_4613),
.D(n_4619),
.Y(n_4653)
);

AOI22xp33_ASAP7_75t_SL g4654 ( 
.A1(n_4635),
.A2(n_4558),
.B1(n_4616),
.B2(n_4507),
.Y(n_4654)
);

NAND4xp25_ASAP7_75t_L g4655 ( 
.A(n_4652),
.B(n_3279),
.C(n_3429),
.D(n_3201),
.Y(n_4655)
);

OAI21xp33_ASAP7_75t_SL g4656 ( 
.A1(n_4631),
.A2(n_4530),
.B(n_4591),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4639),
.B(n_4583),
.Y(n_4657)
);

NAND3xp33_ASAP7_75t_L g4658 ( 
.A(n_4630),
.B(n_3402),
.C(n_3399),
.Y(n_4658)
);

NOR2xp33_ASAP7_75t_L g4659 ( 
.A(n_4646),
.B(n_4583),
.Y(n_4659)
);

NAND4xp25_ASAP7_75t_L g4660 ( 
.A(n_4629),
.B(n_4627),
.C(n_4647),
.D(n_4632),
.Y(n_4660)
);

AOI22xp5_ASAP7_75t_SL g4661 ( 
.A1(n_4640),
.A2(n_3411),
.B1(n_3179),
.B2(n_3321),
.Y(n_4661)
);

NAND4xp25_ASAP7_75t_L g4662 ( 
.A(n_4632),
.B(n_3297),
.C(n_865),
.D(n_862),
.Y(n_4662)
);

AOI21xp33_ASAP7_75t_L g4663 ( 
.A1(n_4643),
.A2(n_863),
.B(n_865),
.Y(n_4663)
);

NOR2xp33_ASAP7_75t_SL g4664 ( 
.A(n_4634),
.B(n_4628),
.Y(n_4664)
);

AOI222xp33_ASAP7_75t_L g4665 ( 
.A1(n_4643),
.A2(n_3803),
.B1(n_3818),
.B2(n_3810),
.C1(n_3838),
.C2(n_3825),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4645),
.B(n_863),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4638),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_SL g4668 ( 
.A(n_4637),
.B(n_4137),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_L g4669 ( 
.A(n_4644),
.B(n_866),
.Y(n_4669)
);

OAI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4637),
.A2(n_3464),
.B(n_3460),
.Y(n_4670)
);

NAND3xp33_ASAP7_75t_L g4671 ( 
.A(n_4633),
.B(n_3835),
.C(n_3824),
.Y(n_4671)
);

AOI21xp5_ASAP7_75t_L g4672 ( 
.A1(n_4664),
.A2(n_4648),
.B(n_4642),
.Y(n_4672)
);

OAI322xp33_ASAP7_75t_L g4673 ( 
.A1(n_4667),
.A2(n_4636),
.A3(n_4649),
.B1(n_4650),
.B2(n_4641),
.C1(n_4626),
.C2(n_3844),
.Y(n_4673)
);

NAND3xp33_ASAP7_75t_SL g4674 ( 
.A(n_4653),
.B(n_4626),
.C(n_867),
.Y(n_4674)
);

AOI222xp33_ASAP7_75t_L g4675 ( 
.A1(n_4659),
.A2(n_4657),
.B1(n_4668),
.B2(n_4669),
.C1(n_4666),
.C2(n_4656),
.Y(n_4675)
);

AOI221xp5_ASAP7_75t_L g4676 ( 
.A1(n_4660),
.A2(n_4663),
.B1(n_4654),
.B2(n_4662),
.C(n_4671),
.Y(n_4676)
);

OAI221xp5_ASAP7_75t_L g4677 ( 
.A1(n_4661),
.A2(n_3556),
.B1(n_3369),
.B2(n_3575),
.C(n_3404),
.Y(n_4677)
);

AOI22xp5_ASAP7_75t_L g4678 ( 
.A1(n_4665),
.A2(n_3150),
.B1(n_3963),
.B2(n_3575),
.Y(n_4678)
);

OAI211xp5_ASAP7_75t_SL g4679 ( 
.A1(n_4670),
.A2(n_869),
.B(n_867),
.C(n_868),
.Y(n_4679)
);

NAND5xp2_ASAP7_75t_L g4680 ( 
.A(n_4658),
.B(n_3142),
.C(n_870),
.D(n_868),
.E(n_869),
.Y(n_4680)
);

OAI211xp5_ASAP7_75t_SL g4681 ( 
.A1(n_4655),
.A2(n_874),
.B(n_871),
.C(n_872),
.Y(n_4681)
);

AOI22xp5_ASAP7_75t_L g4682 ( 
.A1(n_4664),
.A2(n_3556),
.B1(n_3369),
.B2(n_3952),
.Y(n_4682)
);

AOI21xp33_ASAP7_75t_L g4683 ( 
.A1(n_4664),
.A2(n_871),
.B(n_872),
.Y(n_4683)
);

AOI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4664),
.A2(n_3574),
.B1(n_3835),
.B2(n_3276),
.Y(n_4684)
);

O2A1O1Ixp33_ASAP7_75t_L g4685 ( 
.A1(n_4664),
.A2(n_877),
.B(n_875),
.C(n_876),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4667),
.Y(n_4686)
);

OAI221xp5_ASAP7_75t_SL g4687 ( 
.A1(n_4653),
.A2(n_3735),
.B1(n_3771),
.B2(n_3768),
.C(n_3766),
.Y(n_4687)
);

OAI22xp33_ASAP7_75t_L g4688 ( 
.A1(n_4664),
.A2(n_4048),
.B1(n_3835),
.B2(n_3791),
.Y(n_4688)
);

NAND4xp75_ASAP7_75t_L g4689 ( 
.A(n_4672),
.B(n_878),
.C(n_875),
.D(n_876),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4686),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4685),
.Y(n_4691)
);

NAND4xp75_ASAP7_75t_L g4692 ( 
.A(n_4676),
.B(n_882),
.C(n_880),
.D(n_881),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4673),
.Y(n_4693)
);

INVx2_ASAP7_75t_SL g4694 ( 
.A(n_4678),
.Y(n_4694)
);

NAND4xp75_ASAP7_75t_L g4695 ( 
.A(n_4683),
.B(n_885),
.C(n_881),
.D(n_883),
.Y(n_4695)
);

INVxp67_ASAP7_75t_SL g4696 ( 
.A(n_4688),
.Y(n_4696)
);

AOI22xp5_ASAP7_75t_L g4697 ( 
.A1(n_4674),
.A2(n_4048),
.B1(n_3276),
.B2(n_3488),
.Y(n_4697)
);

XNOR2x1_ASAP7_75t_L g4698 ( 
.A(n_4695),
.B(n_4681),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_SL g4699 ( 
.A(n_4693),
.B(n_4675),
.Y(n_4699)
);

XNOR2x1_ASAP7_75t_L g4700 ( 
.A(n_4692),
.B(n_4680),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_SL g4701 ( 
.A(n_4691),
.B(n_4682),
.Y(n_4701)
);

NOR2xp33_ASAP7_75t_R g4702 ( 
.A(n_4690),
.B(n_883),
.Y(n_4702)
);

NOR2xp33_ASAP7_75t_R g4703 ( 
.A(n_4694),
.B(n_885),
.Y(n_4703)
);

NOR2xp33_ASAP7_75t_R g4704 ( 
.A(n_4689),
.B(n_886),
.Y(n_4704)
);

INVxp33_ASAP7_75t_SL g4705 ( 
.A(n_4704),
.Y(n_4705)
);

AOI22x1_ASAP7_75t_L g4706 ( 
.A1(n_4703),
.A2(n_4696),
.B1(n_4687),
.B2(n_4697),
.Y(n_4706)
);

XNOR2xp5_ASAP7_75t_L g4707 ( 
.A(n_4700),
.B(n_4684),
.Y(n_4707)
);

AOI21xp5_ASAP7_75t_L g4708 ( 
.A1(n_4699),
.A2(n_4679),
.B(n_4677),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4698),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4709),
.Y(n_4710)
);

NAND3xp33_ASAP7_75t_L g4711 ( 
.A(n_4707),
.B(n_4701),
.C(n_4702),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4710),
.Y(n_4712)
);

AOI31xp33_ASAP7_75t_L g4713 ( 
.A1(n_4712),
.A2(n_4711),
.A3(n_4708),
.B(n_4705),
.Y(n_4713)
);

OAI322xp33_ASAP7_75t_L g4714 ( 
.A1(n_4713),
.A2(n_4706),
.A3(n_888),
.B1(n_889),
.B2(n_890),
.C1(n_891),
.C2(n_892),
.Y(n_4714)
);

OAI22xp5_ASAP7_75t_SL g4715 ( 
.A1(n_4713),
.A2(n_889),
.B1(n_887),
.B2(n_888),
.Y(n_4715)
);

OAI21xp5_ASAP7_75t_L g4716 ( 
.A1(n_4714),
.A2(n_3485),
.B(n_3471),
.Y(n_4716)
);

INVx2_ASAP7_75t_SL g4717 ( 
.A(n_4716),
.Y(n_4717)
);

OAI221xp5_ASAP7_75t_R g4718 ( 
.A1(n_4717),
.A2(n_4715),
.B1(n_893),
.B2(n_891),
.C(n_892),
.Y(n_4718)
);

AOI211xp5_ASAP7_75t_L g4719 ( 
.A1(n_4718),
.A2(n_895),
.B(n_893),
.C(n_894),
.Y(n_4719)
);


endmodule