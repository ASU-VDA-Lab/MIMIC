module fake_netlist_1_7680_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_30;
wire n_26;
wire n_13;
wire n_33;
wire n_16;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_0), .B(n_7), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_14), .B(n_1), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_13), .A2(n_9), .B(n_2), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_14), .A2(n_1), .B(n_2), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_19), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_19), .B(n_14), .Y(n_25) );
NAND2xp33_ASAP7_75t_R g26 ( .A(n_18), .B(n_17), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_15), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_25), .B(n_15), .Y(n_29) );
OAI21xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_23), .B(n_24), .Y(n_30) );
OAI211xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_28), .B(n_29), .C(n_22), .Y(n_31) );
OAI221xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_26), .B1(n_29), .B2(n_11), .C(n_21), .Y(n_32) );
O2A1O1Ixp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_26), .B(n_4), .C(n_5), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_33), .B(n_3), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_32), .B1(n_12), .B2(n_16), .Y(n_35) );
endmodule