module fake_jpeg_11084_n_515 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_56),
.B(n_61),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_17),
.C(n_1),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_57),
.B(n_28),
.C(n_49),
.Y(n_157)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_60),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_31),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_77),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_1),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_66),
.B(n_84),
.Y(n_162)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_69),
.Y(n_166)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_18),
.Y(n_75)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_25),
.B(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_2),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_25),
.B(n_2),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_2),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_93),
.Y(n_137)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_12),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_92),
.B(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_30),
.B(n_3),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_104),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_95),
.Y(n_195)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_3),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_4),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_110),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

NAND2x1_ASAP7_75t_SL g107 ( 
.A(n_45),
.B(n_33),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_107),
.Y(n_183)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_116),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_45),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_112),
.Y(n_144)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_114),
.Y(n_165)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_119),
.Y(n_155)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_5),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_19),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_83),
.A2(n_27),
.B1(n_40),
.B2(n_35),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_129),
.A2(n_143),
.B1(n_158),
.B2(n_184),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_53),
.B1(n_52),
.B2(n_37),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_130),
.A2(n_148),
.B1(n_150),
.B2(n_153),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_77),
.B(n_32),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_40),
.B1(n_35),
.B2(n_46),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_78),
.A2(n_53),
.B1(n_37),
.B2(n_28),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_79),
.A2(n_29),
.B1(n_46),
.B2(n_43),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_87),
.A2(n_106),
.B1(n_100),
.B2(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_58),
.B(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_156),
.B(n_170),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_157),
.B(n_163),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_98),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_101),
.A2(n_26),
.B1(n_41),
.B2(n_33),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_161),
.A2(n_167),
.B1(n_188),
.B2(n_201),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_60),
.B(n_40),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_19),
.B1(n_32),
.B2(n_29),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_63),
.B1(n_89),
.B2(n_139),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_76),
.A2(n_26),
.B1(n_47),
.B2(n_40),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_86),
.B(n_5),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_68),
.B(n_5),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_67),
.B(n_6),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_91),
.B(n_6),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_194),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_114),
.A2(n_47),
.B1(n_8),
.B2(n_10),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_95),
.B(n_6),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_191),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_111),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_95),
.B(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_72),
.B(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_59),
.B(n_11),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_144),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_99),
.A2(n_12),
.B1(n_102),
.B2(n_64),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_200),
.B1(n_154),
.B2(n_166),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_69),
.A2(n_12),
.B1(n_97),
.B2(n_63),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_71),
.A2(n_115),
.B1(n_80),
.B2(n_108),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_138),
.B1(n_157),
.B2(n_181),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_205),
.A2(n_247),
.B1(n_264),
.B2(n_240),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_132),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_206),
.B(n_223),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_119),
.B1(n_112),
.B2(n_113),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_207),
.A2(n_253),
.B1(n_265),
.B2(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

NAND2x1_ASAP7_75t_L g218 ( 
.A(n_156),
.B(n_89),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_218),
.A2(n_227),
.B(n_231),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_242),
.B1(n_128),
.B2(n_260),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_132),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g299 ( 
.A1(n_224),
.A2(n_237),
.B1(n_258),
.B2(n_269),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_162),
.B(n_194),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_181),
.C(n_170),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_229),
.B(n_231),
.C(n_238),
.Y(n_289)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_163),
.C(n_123),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_232),
.B(n_233),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_155),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_159),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_234),
.B(n_243),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_177),
.B(n_126),
.CI(n_163),
.CON(n_235),
.SN(n_235)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_235),
.A2(n_213),
.B(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_188),
.A2(n_166),
.B1(n_146),
.B2(n_174),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_131),
.B(n_179),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_131),
.B(n_179),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_240),
.B(n_249),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_137),
.B(n_136),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_136),
.A2(n_174),
.B1(n_193),
.B2(n_168),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_140),
.B(n_141),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_248),
.Y(n_307)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_150),
.A2(n_148),
.B1(n_185),
.B2(n_125),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_147),
.A2(n_152),
.B(n_186),
.C(n_142),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_144),
.B(n_152),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_149),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_250),
.B(n_254),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_133),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_193),
.B(n_151),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_267),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_168),
.A2(n_202),
.B1(n_127),
.B2(n_176),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_169),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_259),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_127),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_266),
.C(n_271),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_169),
.A2(n_146),
.B(n_192),
.C(n_151),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_257),
.A2(n_262),
.B(n_264),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_135),
.A2(n_154),
.B1(n_171),
.B2(n_189),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_178),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_264),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_189),
.A2(n_199),
.B1(n_149),
.B2(n_165),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_263),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_182),
.B(n_178),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_134),
.A2(n_202),
.B1(n_176),
.B2(n_125),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_173),
.B(n_165),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_134),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_268),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_173),
.A2(n_185),
.B1(n_199),
.B2(n_149),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_262),
.B1(n_219),
.B2(n_216),
.Y(n_288)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_128),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_221),
.B(n_197),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_276),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_277),
.A2(n_287),
.B1(n_317),
.B2(n_320),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_222),
.B(n_221),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_291),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_283),
.A2(n_311),
.B(n_287),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_227),
.A2(n_219),
.B1(n_216),
.B2(n_222),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_288),
.A2(n_268),
.B1(n_211),
.B2(n_215),
.Y(n_326)
);

AO22x2_ASAP7_75t_L g291 ( 
.A1(n_218),
.A2(n_248),
.B1(n_209),
.B2(n_227),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_226),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_296),
.B(n_303),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_212),
.A2(n_218),
.B1(n_267),
.B2(n_241),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_298),
.A2(n_246),
.B1(n_245),
.B2(n_250),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_299),
.A2(n_214),
.B1(n_230),
.B2(n_256),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_235),
.B(n_212),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_204),
.B(n_235),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_308),
.C(n_303),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_225),
.B(n_252),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_239),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_249),
.B(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_314),
.B(n_298),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_238),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_322),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_242),
.A2(n_240),
.B1(n_238),
.B2(n_257),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_321),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_255),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_277),
.B1(n_320),
.B2(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_261),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_329),
.B(n_330),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_285),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_339),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_259),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_337),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_210),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_347),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_304),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_280),
.B(n_217),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_342),
.B(n_301),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_318),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_352),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_344),
.A2(n_360),
.B1(n_319),
.B2(n_279),
.Y(n_392)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_283),
.C(n_296),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_280),
.B(n_272),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_L g393 ( 
.A1(n_349),
.A2(n_356),
.B(n_302),
.Y(n_393)
);

INVx8_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_307),
.A2(n_317),
.B(n_288),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_351),
.A2(n_358),
.B(n_291),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_289),
.B(n_281),
.C(n_272),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_355),
.Y(n_388)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_306),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_309),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_357),
.A2(n_319),
.B(n_275),
.Y(n_379)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

BUFx12f_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_345),
.A2(n_339),
.B1(n_333),
.B2(n_341),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_362),
.A2(n_374),
.B1(n_381),
.B2(n_383),
.Y(n_417)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_325),
.A2(n_291),
.B1(n_311),
.B2(n_276),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_370),
.A2(n_373),
.B1(n_334),
.B2(n_353),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_325),
.A2(n_291),
.B1(n_276),
.B2(n_314),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_291),
.B1(n_299),
.B2(n_301),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_335),
.B(n_359),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_336),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_393),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_345),
.B1(n_334),
.B2(n_356),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_351),
.A2(n_273),
.B1(n_275),
.B2(n_278),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_351),
.A2(n_278),
.B1(n_284),
.B2(n_279),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_385),
.A2(n_324),
.B1(n_343),
.B2(n_329),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_337),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_327),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_294),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_391),
.A2(n_324),
.B(n_342),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_363),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_415),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_381),
.A2(n_358),
.B1(n_349),
.B2(n_348),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_396),
.A2(n_373),
.B1(n_365),
.B2(n_389),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_347),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_409),
.C(n_420),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_398),
.A2(n_412),
.B(n_413),
.Y(n_433)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_363),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_400),
.B(n_410),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_401),
.B(n_411),
.Y(n_442)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_405),
.A2(n_375),
.B1(n_382),
.B2(n_367),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_406),
.A2(n_416),
.B1(n_418),
.B2(n_383),
.Y(n_431)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_408),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_338),
.C(n_331),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_388),
.B(n_331),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_384),
.A2(n_323),
.B(n_357),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_378),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_419),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_391),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_370),
.A2(n_328),
.B1(n_332),
.B2(n_350),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_368),
.A2(n_350),
.B1(n_359),
.B2(n_330),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_360),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_422),
.A2(n_434),
.B1(n_437),
.B2(n_439),
.Y(n_447)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_377),
.C(n_365),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_428),
.C(n_435),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_377),
.C(n_376),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_412),
.B(n_367),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_404),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_431),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_386),
.B1(n_382),
.B2(n_375),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_374),
.C(n_378),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_379),
.C(n_387),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_404),
.C(n_401),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_402),
.A2(n_385),
.B1(n_392),
.B2(n_362),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_395),
.A2(n_390),
.B1(n_391),
.B2(n_387),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_441),
.A2(n_415),
.B1(n_416),
.B2(n_398),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_432),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_455),
.Y(n_464)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_411),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_457),
.Y(n_473)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_436),
.A2(n_402),
.B1(n_405),
.B2(n_394),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_451),
.A2(n_439),
.B1(n_437),
.B2(n_441),
.Y(n_475)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_453),
.A2(n_431),
.B1(n_417),
.B2(n_421),
.Y(n_469)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_424),
.Y(n_454)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_454),
.Y(n_471)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_396),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_460),
.Y(n_467)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_461),
.B(n_428),
.C(n_427),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_456),
.A2(n_433),
.B(n_413),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_456),
.B(n_434),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_468),
.C(n_408),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_435),
.C(n_438),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_469),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_461),
.B(n_442),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_433),
.C(n_422),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_450),
.C(n_447),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_475),
.A2(n_459),
.B1(n_419),
.B2(n_407),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_476),
.B(n_479),
.Y(n_493)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_478),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_450),
.C(n_447),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_452),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_480),
.B(n_482),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_489)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_449),
.C(n_453),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_449),
.C(n_442),
.Y(n_484)
);

AO221x1_ASAP7_75t_L g485 ( 
.A1(n_470),
.A2(n_448),
.B1(n_421),
.B2(n_443),
.C(n_390),
.Y(n_485)
);

OAI321xp33_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_470),
.A3(n_403),
.B1(n_471),
.B2(n_380),
.C(n_361),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_469),
.B1(n_466),
.B2(n_474),
.Y(n_488)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_488),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_477),
.A2(n_463),
.B(n_462),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_492),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_476),
.A2(n_472),
.B(n_467),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_361),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_483),
.A2(n_475),
.B1(n_471),
.B2(n_468),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_495),
.Y(n_497)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_490),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_500),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_366),
.B(n_372),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_479),
.C(n_484),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_SL g502 ( 
.A1(n_495),
.A2(n_481),
.B(n_380),
.C(n_361),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_502),
.A2(n_380),
.B1(n_294),
.B2(n_489),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_498),
.A2(n_489),
.B(n_487),
.Y(n_503)
);

AOI21x1_ASAP7_75t_L g508 ( 
.A1(n_503),
.A2(n_506),
.B(n_497),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_372),
.C(n_346),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_501),
.A2(n_290),
.B(n_372),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_505),
.A2(n_502),
.B(n_366),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_508),
.A2(n_505),
.B(n_507),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_510),
.B(n_312),
.Y(n_512)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_511),
.A2(n_512),
.B(n_302),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_312),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_310),
.B(n_499),
.Y(n_515)
);


endmodule