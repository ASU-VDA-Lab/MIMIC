module fake_jpeg_304_n_214 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_1),
.B(n_39),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_67),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_65),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_84),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_60),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_55),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_68),
.B1(n_60),
.B2(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_96),
.B1(n_70),
.B2(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_66),
.B1(n_68),
.B2(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_52),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_112),
.Y(n_122)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_0),
.Y(n_128)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_4),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_64),
.Y(n_118)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_70),
.C(n_56),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_87),
.C(n_58),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_131),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_58),
.B1(n_89),
.B2(n_87),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_98),
.Y(n_141)
);

BUFx16f_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_58),
.B1(n_74),
.B2(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_31),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_72),
.B1(n_61),
.B2(n_74),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_74),
.B1(n_61),
.B2(n_75),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_3),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_75),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_136),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_136)
);

AO21x1_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_99),
.B(n_103),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_143),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_149),
.C(n_150),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_114),
.B(n_75),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_14),
.B(n_15),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_27),
.C(n_47),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_25),
.C(n_45),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_8),
.B(n_10),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_144),
.B(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_160),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_159),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_35),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_11),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_174),
.B1(n_178),
.B2(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_177),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_24),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_145),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_17),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_48),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_19),
.B1(n_20),
.B2(n_36),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_150),
.C(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.C(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_162),
.B(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_197),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_169),
.B(n_180),
.C(n_166),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_173),
.C(n_170),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_173),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_199),
.B(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_204),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_197),
.B(n_164),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_195),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_201),
.B1(n_182),
.B2(n_185),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_206),
.B(n_204),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_38),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_40),
.Y(n_214)
);


endmodule