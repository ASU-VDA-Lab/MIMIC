module real_aes_1945_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_639;
wire n_587;
wire n_546;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_0), .A2(n_39), .B1(n_440), .B2(n_582), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_1), .B(n_296), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_2), .A2(n_82), .B1(n_375), .B2(n_399), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_3), .A2(n_7), .B1(n_525), .B2(n_633), .Y(n_632) );
AO22x2_ASAP7_75t_L g268 ( .A1(n_4), .A2(n_177), .B1(n_265), .B2(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g678 ( .A(n_4), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_5), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_6), .A2(n_18), .B1(n_316), .B2(n_557), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_8), .A2(n_42), .B1(n_443), .B2(n_445), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_9), .A2(n_161), .B1(n_314), .B2(n_316), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_10), .A2(n_60), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_11), .A2(n_106), .B1(n_318), .B2(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_12), .A2(n_226), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_13), .A2(n_126), .B1(n_321), .B2(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_14), .A2(n_217), .B1(n_359), .B2(n_360), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_15), .A2(n_110), .B1(n_377), .B2(n_378), .Y(n_508) );
AOI22x1_ASAP7_75t_L g401 ( .A1(n_16), .A2(n_104), .B1(n_377), .B2(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_17), .A2(n_210), .B1(n_367), .B2(n_368), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_19), .A2(n_100), .B1(n_336), .B2(n_339), .Y(n_335) );
AO22x2_ASAP7_75t_L g264 ( .A1(n_20), .A2(n_57), .B1(n_265), .B2(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_20), .B(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_21), .A2(n_109), .B1(n_458), .B2(n_553), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_22), .A2(n_127), .B1(n_261), .B2(n_430), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_23), .A2(n_221), .B1(n_370), .B2(n_371), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_24), .A2(n_169), .B1(n_314), .B2(n_318), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_25), .A2(n_199), .B1(n_321), .B2(n_325), .Y(n_320) );
XNOR2xp5_ASAP7_75t_L g379 ( .A(n_26), .B(n_380), .Y(n_379) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_26), .B(n_380), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_27), .A2(n_30), .B1(n_377), .B2(n_378), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_28), .A2(n_40), .B1(n_321), .B2(n_333), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_29), .A2(n_196), .B1(n_532), .B2(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_31), .A2(n_192), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g426 ( .A1(n_32), .A2(n_146), .B1(n_209), .B2(n_427), .C1(n_428), .C2(n_430), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_33), .A2(n_191), .B1(n_422), .B2(n_525), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_34), .A2(n_223), .B1(n_360), .B2(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_35), .B(n_296), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_36), .A2(n_90), .B1(n_375), .B2(n_399), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_37), .A2(n_117), .B1(n_238), .B2(n_303), .C1(n_307), .C2(n_427), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_38), .A2(n_164), .B1(n_359), .B2(n_360), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_41), .A2(n_107), .B1(n_484), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_43), .A2(n_74), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_44), .A2(n_154), .B1(n_416), .B2(n_417), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_45), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_46), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_47), .A2(n_143), .B1(n_303), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_48), .A2(n_232), .B1(n_284), .B2(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_49), .A2(n_125), .B1(n_465), .B2(n_467), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_50), .A2(n_227), .B1(n_430), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_51), .A2(n_166), .B1(n_629), .B2(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_52), .A2(n_685), .B1(n_703), .B2(n_704), .Y(n_702) );
INVxp67_ASAP7_75t_L g704 ( .A(n_52), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_53), .A2(n_188), .B1(n_389), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_54), .A2(n_129), .B1(n_413), .B2(n_582), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_55), .A2(n_230), .B1(n_447), .B2(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_56), .B(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_58), .A2(n_86), .B1(n_362), .B2(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_59), .A2(n_113), .B1(n_410), .B2(n_411), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_61), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_62), .A2(n_208), .B1(n_367), .B2(n_368), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_63), .A2(n_118), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g644 ( .A(n_64), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_65), .A2(n_105), .B1(n_362), .B2(n_363), .Y(n_502) );
INVx3_ASAP7_75t_L g265 ( .A(n_66), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_67), .A2(n_144), .B1(n_303), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_68), .A2(n_170), .B1(n_330), .B2(n_333), .Y(n_329) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_69), .A2(n_434), .B(n_469), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_69), .B(n_436), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_70), .A2(n_72), .B1(n_460), .B2(n_462), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_71), .A2(n_178), .B1(n_411), .B2(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_73), .A2(n_225), .B1(n_658), .B2(n_659), .Y(n_657) );
XOR2x2_ASAP7_75t_L g517 ( .A(n_75), .B(n_518), .Y(n_517) );
AO222x2_ASAP7_75t_L g353 ( .A1(n_76), .A2(n_124), .B1(n_151), .B2(n_354), .C1(n_355), .C2(n_356), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_77), .A2(n_179), .B1(n_325), .B2(n_444), .Y(n_637) );
INVx1_ASAP7_75t_L g431 ( .A(n_78), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_79), .A2(n_222), .B1(n_261), .B2(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_80), .A2(n_131), .B1(n_362), .B2(n_363), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_81), .A2(n_163), .B1(n_368), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_SL g273 ( .A(n_83), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_83), .B(n_111), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_84), .Y(n_385) );
INVx2_ASAP7_75t_L g249 ( .A(n_85), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_87), .A2(n_158), .B1(n_537), .B2(n_539), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_88), .A2(n_130), .B1(n_411), .B2(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_89), .A2(n_218), .B1(n_374), .B2(n_375), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_91), .A2(n_207), .B1(n_487), .B2(n_489), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_92), .A2(n_214), .B1(n_522), .B2(n_602), .Y(n_653) );
OA22x2_ASAP7_75t_L g256 ( .A1(n_93), .A2(n_257), .B1(n_342), .B2(n_343), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_93), .Y(n_342) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_94), .A2(n_101), .B1(n_284), .B2(n_484), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_95), .A2(n_233), .B1(n_492), .B2(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_96), .A2(n_156), .B1(n_410), .B2(n_413), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_97), .A2(n_172), .B1(n_330), .B2(n_419), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_98), .A2(n_174), .B1(n_416), .B2(n_607), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_99), .A2(n_120), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_102), .A2(n_198), .B1(n_402), .B2(n_451), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_103), .A2(n_147), .B1(n_334), .B2(n_534), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_108), .A2(n_121), .B1(n_410), .B2(n_487), .Y(n_528) );
AO22x2_ASAP7_75t_L g276 ( .A1(n_111), .A2(n_186), .B1(n_265), .B2(n_277), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_112), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_114), .A2(n_204), .B1(n_419), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_115), .A2(n_136), .B1(n_422), .B2(n_483), .Y(n_551) );
OA22x2_ASAP7_75t_L g647 ( .A1(n_116), .A2(n_648), .B1(n_649), .B2(n_668), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_116), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_119), .A2(n_216), .B1(n_321), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_122), .A2(n_148), .B1(n_325), .B2(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_123), .A2(n_142), .B1(n_284), .B2(n_290), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_128), .A2(n_138), .B1(n_316), .B2(n_416), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_132), .A2(n_194), .B1(n_303), .B2(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g274 ( .A(n_133), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_134), .A2(n_168), .B1(n_321), .B2(n_487), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_135), .A2(n_202), .B1(n_355), .B2(n_356), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_137), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_139), .A2(n_141), .B1(n_417), .B2(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_140), .A2(n_159), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_145), .A2(n_187), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_149), .A2(n_184), .B1(n_416), .B2(n_417), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_150), .A2(n_190), .B1(n_303), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_152), .A2(n_211), .B1(n_425), .B2(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g592 ( .A(n_153), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_155), .A2(n_683), .B1(n_684), .B2(n_698), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_155), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_157), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_160), .A2(n_180), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_162), .A2(n_228), .B1(n_303), .B2(n_578), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_165), .A2(n_183), .B1(n_261), .B2(n_278), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_167), .B(n_455), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_171), .A2(n_234), .B1(n_451), .B2(n_535), .Y(n_667) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_173), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_175), .B(n_296), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_176), .A2(n_189), .B1(n_483), .B2(n_484), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_181), .A2(n_200), .B1(n_612), .B2(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_182), .A2(n_197), .B1(n_370), .B2(n_378), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_185), .A2(n_235), .B1(n_532), .B2(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_193), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g674 ( .A(n_193), .Y(n_674) );
OA22x2_ASAP7_75t_L g474 ( .A1(n_195), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_195), .Y(n_475) );
INVx1_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
AND2x2_ASAP7_75t_R g700 ( .A(n_201), .B(n_674), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_203), .A2(n_240), .B1(n_250), .B2(n_680), .C(n_681), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_205), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_206), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_212), .A2(n_237), .B1(n_261), .B2(n_430), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_213), .A2(n_229), .B1(n_261), .B2(n_430), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_215), .B(n_248), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_219), .A2(n_236), .B1(n_375), .B2(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_220), .B(n_354), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_224), .B(n_455), .Y(n_454) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_231), .B(n_544), .Y(n_543) );
CKINVDCx6p67_ASAP7_75t_R g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_244), .B(n_247), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g708 ( .A(n_245), .B(n_247), .Y(n_708) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_246), .B(n_674), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_513), .B(n_671), .Y(n_250) );
OR2x2_ASAP7_75t_L g680 ( .A(n_251), .B(n_513), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_253), .B1(n_472), .B2(n_473), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_345), .B1(n_346), .B2(n_471), .Y(n_253) );
INVx1_ASAP7_75t_SL g471 ( .A(n_254), .Y(n_471) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_311), .Y(n_257) );
NOR3xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_294), .C(n_301), .Y(n_258) );
NOR4xp25_ASAP7_75t_L g343 ( .A(n_259), .B(n_312), .C(n_328), .D(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_283), .Y(n_259) );
BUFx5_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g429 ( .A(n_262), .Y(n_429) );
BUFx3_ASAP7_75t_L g461 ( .A(n_262), .Y(n_461) );
BUFx3_ASAP7_75t_L g656 ( .A(n_262), .Y(n_656) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
AND2x4_ASAP7_75t_L g304 ( .A(n_263), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g341 ( .A(n_263), .B(n_324), .Y(n_341) );
AND2x4_ASAP7_75t_L g356 ( .A(n_263), .B(n_270), .Y(n_356) );
AND2x2_ASAP7_75t_L g359 ( .A(n_263), .B(n_305), .Y(n_359) );
AND2x2_ASAP7_75t_L g371 ( .A(n_263), .B(n_324), .Y(n_371) );
AND2x2_ASAP7_75t_L g392 ( .A(n_263), .B(n_305), .Y(n_392) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
AND2x2_ASAP7_75t_L g281 ( .A(n_264), .B(n_268), .Y(n_281) );
INVx1_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
INVx1_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
INVx2_ASAP7_75t_L g266 ( .A(n_265), .Y(n_266) );
INVx1_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
OAI22x1_ASAP7_75t_L g271 ( .A1(n_265), .A2(n_272), .B1(n_273), .B2(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_265), .Y(n_272) );
INVx1_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
AND2x4_ASAP7_75t_L g299 ( .A(n_267), .B(n_300), .Y(n_299) );
INVxp67_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g293 ( .A(n_268), .B(n_289), .Y(n_293) );
AND2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g332 ( .A(n_270), .B(n_299), .Y(n_332) );
AND2x4_ASAP7_75t_L g362 ( .A(n_270), .B(n_293), .Y(n_362) );
AND2x2_ASAP7_75t_L g374 ( .A(n_270), .B(n_299), .Y(n_374) );
AND2x2_ASAP7_75t_L g399 ( .A(n_270), .B(n_299), .Y(n_399) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
AND2x2_ASAP7_75t_L g286 ( .A(n_271), .B(n_276), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_271), .Y(n_306) );
AND2x4_ASAP7_75t_L g324 ( .A(n_275), .B(n_306), .Y(n_324) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g305 ( .A(n_276), .B(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g319 ( .A(n_276), .Y(n_319) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g463 ( .A(n_279), .Y(n_463) );
INVx2_ASAP7_75t_L g481 ( .A(n_279), .Y(n_481) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_280), .Y(n_430) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x4_ASAP7_75t_L g318 ( .A(n_281), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g334 ( .A(n_281), .B(n_324), .Y(n_334) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_281), .B(n_282), .Y(n_355) );
AND2x4_ASAP7_75t_L g368 ( .A(n_281), .B(n_319), .Y(n_368) );
AND2x4_ASAP7_75t_L g375 ( .A(n_281), .B(n_324), .Y(n_375) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_281), .B(n_282), .Y(n_389) );
BUFx2_ASAP7_75t_SL g659 ( .A(n_284), .Y(n_659) );
BUFx6f_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
BUFx3_ASAP7_75t_L g468 ( .A(n_285), .Y(n_468) );
BUFx4f_ASAP7_75t_L g483 ( .A(n_285), .Y(n_483) );
INVx2_ASAP7_75t_L g526 ( .A(n_285), .Y(n_526) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g298 ( .A(n_286), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g309 ( .A(n_286), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g354 ( .A(n_286), .B(n_299), .Y(n_354) );
AND2x2_ASAP7_75t_L g360 ( .A(n_286), .B(n_310), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_286), .B(n_287), .Y(n_363) );
AND2x2_ASAP7_75t_L g394 ( .A(n_286), .B(n_287), .Y(n_394) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g466 ( .A(n_291), .Y(n_466) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_292), .Y(n_422) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_292), .Y(n_484) );
AND2x2_ASAP7_75t_L g315 ( .A(n_293), .B(n_305), .Y(n_315) );
AND2x4_ASAP7_75t_L g327 ( .A(n_293), .B(n_324), .Y(n_327) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_293), .B(n_305), .Y(n_367) );
AND2x6_ASAP7_75t_L g378 ( .A(n_293), .B(n_324), .Y(n_378) );
AND2x2_ASAP7_75t_L g507 ( .A(n_293), .B(n_305), .Y(n_507) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_295), .B(n_302), .Y(n_344) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_296), .Y(n_652) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx4_ASAP7_75t_SL g427 ( .A(n_297), .Y(n_427) );
INVx3_ASAP7_75t_L g455 ( .A(n_297), .Y(n_455) );
INVx3_ASAP7_75t_SL g626 ( .A(n_297), .Y(n_626) );
INVx6_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_L g323 ( .A(n_299), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g338 ( .A(n_299), .B(n_305), .Y(n_338) );
AND2x2_ASAP7_75t_L g370 ( .A(n_299), .B(n_324), .Y(n_370) );
AND2x6_ASAP7_75t_L g377 ( .A(n_299), .B(n_305), .Y(n_377) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g424 ( .A(n_304), .Y(n_424) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_304), .Y(n_458) );
BUFx2_ASAP7_75t_L g602 ( .A(n_304), .Y(n_602) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g425 ( .A(n_308), .Y(n_425) );
INVx1_ASAP7_75t_L g522 ( .A(n_308), .Y(n_522) );
INVx2_ASAP7_75t_SL g553 ( .A(n_308), .Y(n_553) );
INVx2_ASAP7_75t_L g578 ( .A(n_308), .Y(n_578) );
INVx2_ASAP7_75t_L g603 ( .A(n_308), .Y(n_603) );
INVx2_ASAP7_75t_L g689 ( .A(n_308), .Y(n_689) );
INVx6_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_328), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_320), .Y(n_312) );
BUFx2_ASAP7_75t_L g665 ( .A(n_314), .Y(n_665) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_315), .Y(n_416) );
INVx2_ASAP7_75t_L g449 ( .A(n_315), .Y(n_449) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g417 ( .A(n_317), .Y(n_417) );
INVx5_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g539 ( .A(n_318), .Y(n_539) );
BUFx2_ASAP7_75t_L g607 ( .A(n_318), .Y(n_607) );
BUFx3_ASAP7_75t_L g639 ( .A(n_318), .Y(n_639) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx4_ASAP7_75t_L g439 ( .A(n_322), .Y(n_439) );
INVx2_ASAP7_75t_L g587 ( .A(n_322), .Y(n_587) );
INVx3_ASAP7_75t_SL g612 ( .A(n_322), .Y(n_612) );
INVx2_ASAP7_75t_SL g663 ( .A(n_322), .Y(n_663) );
INVx8_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g413 ( .A(n_326), .Y(n_413) );
INVx2_ASAP7_75t_L g445 ( .A(n_326), .Y(n_445) );
INVx2_ASAP7_75t_SL g487 ( .A(n_326), .Y(n_487) );
INVx2_ASAP7_75t_SL g583 ( .A(n_326), .Y(n_583) );
INVx8_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_335), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g492 ( .A(n_331), .Y(n_492) );
INVx3_ASAP7_75t_L g534 ( .A(n_331), .Y(n_534) );
INVx6_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g451 ( .A(n_332), .Y(n_451) );
BUFx3_ASAP7_75t_L g696 ( .A(n_332), .Y(n_696) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g419 ( .A(n_334), .Y(n_419) );
BUFx2_ASAP7_75t_SL g452 ( .A(n_334), .Y(n_452) );
INVx2_ASAP7_75t_L g494 ( .A(n_334), .Y(n_494) );
BUFx2_ASAP7_75t_SL g562 ( .A(n_334), .Y(n_562) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
INVx2_ASAP7_75t_SL g489 ( .A(n_337), .Y(n_489) );
INVx3_ASAP7_75t_L g582 ( .A(n_337), .Y(n_582) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g444 ( .A(n_338), .Y(n_444) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_341), .Y(n_402) );
BUFx3_ASAP7_75t_L g411 ( .A(n_341), .Y(n_411) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_341), .Y(n_532) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI22x1_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_432), .B1(n_433), .B2(n_470), .Y(n_346) );
INVx2_ASAP7_75t_L g470 ( .A(n_347), .Y(n_470) );
XNOR2x1_ASAP7_75t_L g347 ( .A(n_348), .B(n_406), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_379), .B(n_404), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_349), .B(n_405), .Y(n_404) );
XNOR2x1_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_364), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_357), .Y(n_352) );
INVx2_ASAP7_75t_SL g384 ( .A(n_354), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_356), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_372), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_381), .B(n_395), .Y(n_380) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_390), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_385), .B2(n_386), .C1(n_387), .C2(n_388), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_384), .A2(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_386), .Y(n_598) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx2_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
XOR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_431), .Y(n_406) );
NAND4xp75_ASAP7_75t_L g407 ( .A(n_408), .B(n_414), .C(n_420), .D(n_426), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .Y(n_408) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
BUFx6f_ASAP7_75t_SL g633 ( .A(n_422), .Y(n_633) );
INVx1_ASAP7_75t_L g547 ( .A(n_427), .Y(n_547) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g573 ( .A(n_429), .Y(n_573) );
BUFx3_ASAP7_75t_L g629 ( .A(n_430), .Y(n_629) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_453), .Y(n_436) );
NAND4xp25_ASAP7_75t_SL g437 ( .A(n_438), .B(n_442), .C(n_446), .D(n_450), .Y(n_437) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_439), .Y(n_564) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g538 ( .A(n_449), .Y(n_538) );
NAND4xp25_ASAP7_75t_SL g453 ( .A(n_454), .B(n_456), .C(n_459), .D(n_464), .Y(n_453) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx6f_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
XNOR2x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_495), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .C(n_482), .Y(n_478) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_484), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .C(n_490), .D(n_491), .Y(n_485) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g535 ( .A(n_494), .Y(n_535) );
XOR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_512), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g496 ( .A(n_497), .B(n_504), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
AOI22xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_615), .B1(n_616), .B2(n_670), .Y(n_513) );
INVx1_ASAP7_75t_L g670 ( .A(n_514), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_566), .B1(n_613), .B2(n_614), .Y(n_514) );
INVx1_ASAP7_75t_L g613 ( .A(n_515), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_540), .B1(n_541), .B2(n_565), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
NOR2xp67_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
NAND4xp25_ASAP7_75t_SL g519 ( .A(n_520), .B(n_521), .C(n_523), .D(n_524), .Y(n_519) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .C(n_533), .D(n_536), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_532), .Y(n_642) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g558 ( .A(n_538), .Y(n_558) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
OAI21xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_548), .B(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g614 ( .A(n_566), .Y(n_614) );
OA22x2_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_590), .B2(n_591), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_589), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_579), .Y(n_569) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
XNOR2x1_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_604), .Y(n_593) );
NOR2xp67_ASAP7_75t_L g594 ( .A(n_595), .B(n_599), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_609), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_645), .B1(n_646), .B2(n_669), .Y(n_616) );
INVx3_ASAP7_75t_L g669 ( .A(n_617), .Y(n_669) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_644), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_619), .B(n_635), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_631), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B1(n_624), .B2(n_627), .C1(n_628), .C2(n_630), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_640), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g668 ( .A(n_649), .Y(n_668) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_660), .Y(n_649) );
NAND4xp25_ASAP7_75t_SL g650 ( .A(n_651), .B(n_653), .C(n_654), .D(n_657), .Y(n_650) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .C(n_666), .D(n_667), .Y(n_660) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_673), .B(n_676), .Y(n_707) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI222xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_699), .B1(n_701), .B2(n_704), .C1(n_705), .C2(n_708), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g703 ( .A(n_685), .Y(n_703) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_686), .B(n_692), .Y(n_685) );
NAND4xp25_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .C(n_690), .D(n_691), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .C(n_695), .D(n_697), .Y(n_692) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
CKINVDCx6p67_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
endmodule