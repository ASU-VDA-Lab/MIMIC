module fake_netlist_5_566_n_2040 (n_137, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2040);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2040;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_96),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_11),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_82),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_158),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_166),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_32),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_62),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_107),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_97),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_48),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_7),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_10),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_119),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_144),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_208),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_151),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_85),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_114),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_10),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_20),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_26),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_110),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_104),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_52),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_25),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_33),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_159),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_50),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_160),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_112),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_115),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_150),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_63),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_66),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_178),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_125),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_21),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_128),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_111),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_155),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_108),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_60),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_94),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_141),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_124),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_181),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_17),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_86),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_44),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_176),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_133),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_31),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_36),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_72),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_106),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_37),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_74),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_54),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_56),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_80),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_89),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_182),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_34),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_19),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_126),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_91),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_170),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_51),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_59),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_113),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_75),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_116),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_88),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_193),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_57),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_180),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_77),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_93),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_54),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_24),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_95),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_46),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_194),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_37),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_29),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_27),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_67),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_129),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_117),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_61),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_22),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_103),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_140),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_29),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_83),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_57),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_109),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_207),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_49),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_162),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_130),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_17),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_120),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_161),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_65),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_15),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_92),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_8),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_135),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_90),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_69),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_209),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_73),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_62),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_1),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_201),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_99),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_79),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_71),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_87),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_138),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_72),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_197),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_0),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_74),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_105),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_16),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_184),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_199),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_189),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_147),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_8),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_142),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_98),
.Y(n_364)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_172),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_202),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_46),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_35),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_35),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_43),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_9),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_139),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_18),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_206),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_59),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_70),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_41),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_5),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_58),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_169),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_23),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_7),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_63),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_31),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_171),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_56),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_131),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_9),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_67),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_25),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_175),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_42),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_165),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_185),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_5),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_148),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_179),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_164),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_156),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_177),
.Y(n_401)
);

BUFx8_ASAP7_75t_SL g402 ( 
.A(n_21),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_42),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_32),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_187),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_47),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_4),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_200),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_146),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_41),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_134),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_30),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_6),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_30),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_43),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_228),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_402),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_218),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_245),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_218),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_218),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_245),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_210),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_218),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_213),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_218),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_278),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_290),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_214),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_273),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_231),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_391),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_246),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_407),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_215),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_407),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_219),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_220),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_273),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_216),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_224),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_268),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_216),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_212),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_268),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_295),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_226),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_227),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_289),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_229),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_295),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_302),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_302),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_222),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_222),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_239),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_240),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_393),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_308),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_235),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_328),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_235),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_403),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_242),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_248),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_237),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_249),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_251),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_237),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_254),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_241),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_365),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_258),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_241),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_330),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_211),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_252),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_261),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_252),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_263),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_264),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_322),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_263),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_383),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_278),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_280),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_280),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_281),
.Y(n_505)
);

INVxp33_ASAP7_75t_SL g506 ( 
.A(n_221),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_281),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_223),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_282),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_336),
.Y(n_510)
);

INVxp33_ASAP7_75t_SL g511 ( 
.A(n_232),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_266),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_267),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_282),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_269),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_287),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_278),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_287),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_288),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_288),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_418),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_418),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_420),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_423),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_421),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_425),
.B(n_290),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_436),
.B(n_336),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_427),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_475),
.A2(n_292),
.B1(n_343),
.B2(n_277),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_R g538 ( 
.A(n_416),
.B(n_270),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_493),
.B(n_339),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_436),
.B(n_339),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_456),
.B(n_411),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_429),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_SL g544 ( 
.A(n_480),
.B(n_247),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_419),
.A2(n_369),
.B1(n_344),
.B2(n_374),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_438),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_432),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_433),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_434),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_454),
.A2(n_238),
.B1(n_243),
.B2(n_236),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_446),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_417),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_448),
.B(n_296),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_435),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_456),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_435),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_437),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

AND2x2_ASAP7_75t_SL g571 ( 
.A(n_502),
.B(n_411),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_R g572 ( 
.A(n_478),
.B(n_274),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_428),
.B(n_247),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_517),
.B(n_294),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_441),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_457),
.A2(n_253),
.B1(n_257),
.B2(n_244),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_506),
.B(n_316),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_510),
.A2(n_271),
.B1(n_276),
.B2(n_259),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_467),
.A2(n_415),
.B1(n_414),
.B2(n_413),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_449),
.B(n_296),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_422),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_445),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_453),
.B(n_459),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_463),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_460),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_462),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_479),
.B(n_330),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_447),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_447),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_499),
.B(n_217),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_450),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_489),
.B(n_394),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_489),
.B(n_394),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_509),
.B(n_348),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_473),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_511),
.B(n_316),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_474),
.B(n_392),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_539),
.B(n_481),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_596),
.B(n_487),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_599),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_522),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_524),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_578),
.B(n_498),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_522),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_524),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_523),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_530),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_605),
.B(n_513),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_525),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_530),
.Y(n_618)
);

INVx8_ASAP7_75t_L g619 ( 
.A(n_526),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_572),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_523),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_596),
.B(n_515),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_532),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_535),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_596),
.B(n_501),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_525),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_535),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_604),
.B(n_392),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_528),
.B(n_563),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_527),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_599),
.B(n_305),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_599),
.B(n_275),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_536),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_599),
.B(n_279),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_600),
.B(n_285),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_529),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_556),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_602),
.B(n_592),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_574),
.B(n_428),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_538),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_531),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_542),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_600),
.B(n_291),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_571),
.B(n_482),
.Y(n_651)
);

INVx6_ASAP7_75t_L g652 ( 
.A(n_600),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_600),
.A2(n_540),
.B1(n_533),
.B2(n_602),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_582),
.B(n_300),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_587),
.B(n_301),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_558),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_546),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_558),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_533),
.B(n_303),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_592),
.B(n_452),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_567),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_567),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_571),
.B(n_484),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_547),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_SL g666 ( 
.A1(n_541),
.A2(n_560),
.B1(n_580),
.B2(n_576),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_542),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_546),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_589),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_543),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_530),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_540),
.A2(n_439),
.B1(n_451),
.B2(n_348),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_543),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_545),
.B(n_304),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_546),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_571),
.A2(n_283),
.B1(n_298),
.B2(n_293),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_550),
.B(n_485),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_546),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_588),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_545),
.B(n_311),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_576),
.A2(n_307),
.B1(n_312),
.B2(n_310),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_551),
.B(n_320),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_588),
.Y(n_684)
);

NOR2x1p5_ASAP7_75t_L g685 ( 
.A(n_573),
.B(n_569),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_588),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_321),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g688 ( 
.A(n_565),
.B(n_490),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_561),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_598),
.A2(n_314),
.B1(n_315),
.B2(n_297),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_573),
.B(n_365),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_590),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_555),
.B(n_564),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_598),
.A2(n_314),
.B1(n_315),
.B2(n_297),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_549),
.B(n_495),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_603),
.B(n_512),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_569),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_591),
.Y(n_701)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_564),
.A2(n_230),
.B(n_225),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_SL g703 ( 
.A1(n_580),
.A2(n_225),
.B1(n_234),
.B2(n_230),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_568),
.B(n_323),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_568),
.B(n_325),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_562),
.B(n_494),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_570),
.B(n_329),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_570),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_565),
.B(n_294),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_588),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_575),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_575),
.B(n_332),
.Y(n_712)
);

AND3x2_ASAP7_75t_L g713 ( 
.A(n_521),
.B(n_233),
.C(n_217),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_547),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_577),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_SL g716 ( 
.A1(n_537),
.A2(n_440),
.B1(n_461),
.B2(n_442),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_548),
.A2(n_331),
.B1(n_313),
.B2(n_324),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_577),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_585),
.A2(n_334),
.B1(n_384),
.B2(n_385),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_601),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_601),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_562),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_579),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_530),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_548),
.B(n_233),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_579),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_581),
.B(n_505),
.C(n_327),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_544),
.B(n_335),
.C(n_318),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_530),
.Y(n_729)
);

BUFx6f_ASAP7_75t_SL g730 ( 
.A(n_583),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_SL g731 ( 
.A(n_537),
.B(n_470),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_583),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_584),
.Y(n_733)
);

HB1xp67_ASAP7_75t_SL g734 ( 
.A(n_584),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_586),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_586),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_593),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_593),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_594),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_534),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_594),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_534),
.A2(n_372),
.B1(n_387),
.B2(n_342),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_534),
.B(n_472),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_534),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_534),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_552),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_552),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_552),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_552),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_552),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_553),
.B(n_333),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_553),
.Y(n_752)
);

BUFx4f_ASAP7_75t_L g753 ( 
.A(n_553),
.Y(n_753)
);

AO22x2_ASAP7_75t_L g754 ( 
.A1(n_553),
.A2(n_319),
.B1(n_337),
.B2(n_406),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_553),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_559),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_559),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_608),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_630),
.B(n_354),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_355),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_616),
.B(n_597),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_611),
.B(n_607),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_653),
.B(n_362),
.C(n_357),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_608),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_666),
.B(n_338),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_SL g767 ( 
.A(n_652),
.B(n_338),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_720),
.B(n_597),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_725),
.A2(n_341),
.B1(n_409),
.B2(n_265),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_720),
.B(n_597),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_721),
.B(n_597),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_658),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_652),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_623),
.B(n_368),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_643),
.A2(n_345),
.B1(n_346),
.B2(n_408),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_643),
.B(n_703),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_656),
.B(n_370),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_721),
.B(n_559),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_626),
.B(n_378),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_620),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_629),
.B(n_597),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_699),
.B(n_338),
.Y(n_782)
);

NAND2x1_ASAP7_75t_L g783 ( 
.A(n_652),
.B(n_559),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_665),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_652),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_699),
.B(n_338),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_619),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_655),
.B(n_559),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_677),
.B(n_380),
.C(n_379),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_610),
.B(n_595),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_725),
.A2(n_389),
.B(n_319),
.C(n_337),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_610),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_736),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_736),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_615),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_714),
.B(n_472),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_714),
.B(n_278),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_685),
.A2(n_347),
.B1(n_350),
.B2(n_405),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_644),
.B(n_734),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_613),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_613),
.B(n_566),
.Y(n_801)
);

O2A1O1Ixp5_ASAP7_75t_L g802 ( 
.A1(n_634),
.A2(n_627),
.B(n_631),
.C(n_617),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_658),
.B(n_338),
.Y(n_803)
);

INVx6_ASAP7_75t_L g804 ( 
.A(n_736),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_718),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_617),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_658),
.B(n_397),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_627),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_647),
.B(n_382),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_665),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_631),
.B(n_595),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_677),
.B(n_412),
.C(n_250),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_632),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_632),
.B(n_566),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_735),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_633),
.B(n_566),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_725),
.A2(n_265),
.B1(n_409),
.B2(n_272),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_633),
.B(n_640),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_735),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_635),
.B(n_397),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_737),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_737),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_682),
.B(n_250),
.C(n_234),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_640),
.B(n_566),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_L g825 ( 
.A(n_685),
.B(n_365),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_697),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_738),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_645),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_645),
.B(n_566),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_692),
.A2(n_358),
.B1(n_360),
.B2(n_361),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_620),
.B(n_294),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_660),
.B(n_363),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_692),
.A2(n_272),
.B1(n_286),
.B2(n_341),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_709),
.B(n_727),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_661),
.A2(n_286),
.B1(n_256),
.B2(n_260),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_637),
.B(n_397),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_648),
.B(n_649),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_648),
.B(n_595),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_738),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_741),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_638),
.B(n_397),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_690),
.B(n_364),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_667),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_667),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_671),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_671),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_674),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_674),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_719),
.B(n_367),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_689),
.B(n_595),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_689),
.B(n_595),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_694),
.B(n_255),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_694),
.B(n_255),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_690),
.B(n_373),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_700),
.B(n_256),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_708),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_708),
.B(n_260),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_661),
.B(n_477),
.Y(n_859)
);

AND2x6_ASAP7_75t_SL g860 ( 
.A(n_706),
.B(n_340),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_711),
.B(n_262),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_711),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_650),
.B(n_397),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_715),
.A2(n_262),
.B1(n_284),
.B2(n_401),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_651),
.B(n_381),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_664),
.B(n_386),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_715),
.B(n_365),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_619),
.B(n_284),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_723),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_723),
.B(n_365),
.Y(n_870)
);

AOI221xp5_ASAP7_75t_L g871 ( 
.A1(n_717),
.A2(n_673),
.B1(n_691),
.B2(n_696),
.C(n_682),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_726),
.B(n_483),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_728),
.B(n_388),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_726),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_732),
.B(n_365),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_732),
.B(n_733),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_733),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_739),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_739),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_754),
.B(n_483),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_748),
.B(n_365),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_743),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_609),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_675),
.B(n_299),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_743),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_713),
.B(n_299),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_695),
.Y(n_887)
);

AOI221xp5_ASAP7_75t_L g888 ( 
.A1(n_717),
.A2(n_404),
.B1(n_340),
.B2(n_352),
.C(n_366),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_688),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_609),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_748),
.B(n_306),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_701),
.B(n_486),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_701),
.B(n_486),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_678),
.B(n_395),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_619),
.Y(n_895)
);

OAI21xp33_ASAP7_75t_SL g896 ( 
.A1(n_681),
.A2(n_687),
.B(n_683),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_698),
.B(n_742),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_704),
.B(n_306),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_749),
.B(n_365),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_705),
.B(n_707),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_712),
.A2(n_401),
.B1(n_309),
.B2(n_317),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_L g902 ( 
.A(n_749),
.B(n_309),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_754),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_612),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_729),
.B(n_756),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_750),
.B(n_398),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_751),
.B(n_317),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_612),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_754),
.B(n_488),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_619),
.B(n_326),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_614),
.Y(n_911)
);

OAI22xp33_ASAP7_75t_L g912 ( 
.A1(n_731),
.A2(n_326),
.B1(n_349),
.B2(n_359),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_614),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_730),
.A2(n_399),
.B1(n_349),
.B2(n_353),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_754),
.B(n_488),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_621),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_621),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_744),
.B(n_353),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_693),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_622),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_622),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_744),
.B(n_356),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_624),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_750),
.B(n_356),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_730),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_763),
.B(n_752),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_856),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_856),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_857),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_795),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_760),
.A2(n_730),
.B1(n_746),
.B2(n_745),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_759),
.B(n_745),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_857),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_896),
.B(n_752),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_758),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_758),
.Y(n_936)
);

INVxp33_ASAP7_75t_SL g937 ( 
.A(n_919),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_862),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_887),
.B(n_746),
.Y(n_939)
);

BUFx10_ASAP7_75t_L g940 ( 
.A(n_809),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_900),
.B(n_757),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_793),
.B(n_757),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_766),
.A2(n_352),
.B1(n_404),
.B2(n_366),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_834),
.A2(n_693),
.B1(n_755),
.B2(n_716),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_871),
.A2(n_888),
.B(n_791),
.C(n_823),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_862),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_877),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_793),
.B(n_693),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_777),
.B(n_747),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_826),
.B(n_693),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_879),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_879),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_761),
.Y(n_953)
);

OR2x6_ASAP7_75t_L g954 ( 
.A(n_787),
.B(n_706),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_758),
.A2(n_400),
.B1(n_359),
.B2(n_753),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_761),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_832),
.B(n_747),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_792),
.B(n_800),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_805),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_815),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_815),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_880),
.B(n_400),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_804),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_787),
.B(n_706),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_895),
.B(n_491),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_806),
.B(n_747),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_819),
.Y(n_967)
);

OR2x2_ASAP7_75t_SL g968 ( 
.A(n_812),
.B(n_376),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_808),
.B(n_813),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_895),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_892),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_819),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_828),
.B(n_755),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_821),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_804),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_882),
.B(n_491),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_794),
.B(n_753),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_762),
.A2(n_753),
.B(n_618),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_885),
.B(n_676),
.Y(n_979)
);

AND2x4_ASAP7_75t_SL g980 ( 
.A(n_893),
.B(n_722),
.Y(n_980)
);

BUFx8_ASAP7_75t_L g981 ( 
.A(n_797),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_843),
.B(n_679),
.Y(n_982)
);

AND3x1_ASAP7_75t_L g983 ( 
.A(n_799),
.B(n_376),
.C(n_377),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_776),
.A2(n_897),
.B1(n_825),
.B2(n_774),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_794),
.B(n_496),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_769),
.A2(n_628),
.B1(n_624),
.B2(n_639),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_802),
.B(n_679),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_821),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_804),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_919),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_859),
.B(n_722),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_776),
.A2(n_680),
.B1(n_684),
.B2(n_686),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_844),
.B(n_680),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_859),
.B(n_496),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_822),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_780),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_780),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_822),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_791),
.A2(n_396),
.B(n_377),
.C(n_406),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_827),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_903),
.B(n_784),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_827),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_795),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_839),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_785),
.B(n_684),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_766),
.A2(n_817),
.B1(n_903),
.B2(n_880),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_839),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_785),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_840),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_796),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_889),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_909),
.A2(n_396),
.B(n_389),
.C(n_390),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_845),
.B(n_686),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_840),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_846),
.B(n_710),
.Y(n_1015)
);

AND2x6_ASAP7_75t_L g1016 ( 
.A(n_909),
.B(n_710),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_860),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_810),
.B(n_722),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_795),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_883),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_847),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_848),
.Y(n_1022)
);

OR2x6_ASAP7_75t_SL g1023 ( 
.A(n_789),
.B(n_390),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_785),
.B(n_740),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_795),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_779),
.B(n_497),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_869),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_915),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_868),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_874),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_SL g1031 ( 
.A(n_831),
.B(n_925),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_890),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_878),
.B(n_625),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_908),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_818),
.B(n_625),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_890),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_911),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_842),
.B(n_702),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_837),
.B(n_628),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_904),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_915),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_868),
.B(n_497),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_912),
.A2(n_663),
.B1(n_646),
.B2(n_636),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_886),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_904),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_917),
.Y(n_1046)
);

BUFx8_ASAP7_75t_SL g1047 ( 
.A(n_868),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_785),
.B(n_615),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_833),
.A2(n_663),
.B1(n_646),
.B2(n_636),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_825),
.A2(n_618),
.B1(n_662),
.B2(n_659),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_920),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_886),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_921),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_773),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_872),
.Y(n_1055)
);

NOR2x2_ASAP7_75t_L g1056 ( 
.A(n_868),
.B(n_294),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_913),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_788),
.A2(n_618),
.B(n_724),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_765),
.A2(n_662),
.B1(n_641),
.B2(n_642),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_872),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_773),
.B(n_615),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_913),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_916),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_773),
.B(n_615),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_876),
.B(n_639),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_916),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_910),
.B(n_500),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_886),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_923),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_SL g1070 ( 
.A1(n_865),
.A2(n_351),
.B1(n_516),
.B2(n_514),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_907),
.A2(n_702),
.B(n_642),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_910),
.B(n_500),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_923),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_884),
.B(n_898),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_852),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_891),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_910),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_891),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_772),
.B(n_641),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_853),
.B(n_855),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_866),
.B(n_740),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_858),
.B(n_654),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_891),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_781),
.B(n_740),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_783),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_790),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_924),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_905),
.A2(n_615),
.B(n_724),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_801),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_861),
.B(n_654),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_835),
.A2(n_764),
.B1(n_775),
.B2(n_849),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_811),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_924),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_873),
.B(n_78),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_768),
.B(n_657),
.Y(n_1095)
);

AO22x1_ASAP7_75t_L g1096 ( 
.A1(n_924),
.A2(n_507),
.B1(n_518),
.B2(n_516),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_770),
.B(n_657),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_924),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_798),
.B(n_914),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_814),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_816),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_824),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_829),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_771),
.B(n_659),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_778),
.B(n_669),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_924),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_838),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_924),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_850),
.B(n_669),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_851),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_918),
.B(n_670),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_975),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_L g1113 ( 
.A(n_971),
.B(n_854),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_996),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_950),
.A2(n_1099),
.B(n_767),
.C(n_1071),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_944),
.B(n_894),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_927),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1006),
.A2(n_864),
.B1(n_910),
.B2(n_922),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1099),
.A2(n_901),
.B1(n_906),
.B2(n_867),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_975),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_991),
.B(n_830),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_927),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1011),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1074),
.B(n_867),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_984),
.B(n_906),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_945),
.A2(n_875),
.B(n_870),
.C(n_786),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1006),
.A2(n_841),
.B1(n_820),
.B2(n_836),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_989),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1010),
.B(n_782),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_957),
.A2(n_820),
.B(n_836),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1025),
.A2(n_841),
.B(n_863),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1017),
.A2(n_937),
.B1(n_983),
.B2(n_996),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_933),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1055),
.B(n_786),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_945),
.A2(n_863),
.B(n_875),
.C(n_870),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_940),
.B(n_351),
.Y(n_1137)
);

INVx5_ASAP7_75t_L g1138 ( 
.A(n_1016),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1060),
.B(n_670),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_940),
.B(n_803),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_933),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_951),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1091),
.A2(n_899),
.B1(n_881),
.B2(n_902),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1025),
.A2(n_672),
.B(n_740),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1025),
.A2(n_672),
.B(n_740),
.Y(n_1145)
);

INVx6_ASAP7_75t_L g1146 ( 
.A(n_963),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_952),
.Y(n_1148)
);

CKINVDCx16_ASAP7_75t_R g1149 ( 
.A(n_997),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_950),
.B(n_351),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1087),
.A2(n_1093),
.B(n_1108),
.C(n_1106),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1075),
.B(n_807),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_994),
.B(n_902),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_943),
.A2(n_899),
.B1(n_504),
.B2(n_503),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_994),
.B(n_672),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_997),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_952),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_928),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_943),
.A2(n_503),
.B1(n_504),
.B2(n_507),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1081),
.A2(n_468),
.B(n_452),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_929),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1028),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_963),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1041),
.A2(n_968),
.B1(n_969),
.B2(n_958),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1012),
.A2(n_520),
.B(n_519),
.C(n_518),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_985),
.B(n_965),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_985),
.B(n_351),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1025),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1041),
.B(n_672),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1083),
.A2(n_1070),
.B1(n_1021),
.B2(n_1027),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_976),
.B(n_514),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_938),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1081),
.A2(n_724),
.B(n_672),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_989),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_1016),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_978),
.A2(n_724),
.B(n_668),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1020),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1083),
.A2(n_519),
.B1(n_520),
.B2(n_455),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_981),
.B(n_466),
.C(n_458),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1022),
.B(n_1030),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1020),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_937),
.B(n_724),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_981),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1016),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_965),
.B(n_1031),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1080),
.A2(n_668),
.B(n_469),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1052),
.B(n_970),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1023),
.A2(n_465),
.B1(n_469),
.B2(n_468),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1044),
.A2(n_668),
.B1(n_466),
.B2(n_465),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1086),
.B(n_668),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1001),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1058),
.A2(n_464),
.B(n_458),
.Y(n_1192)
);

AO21x1_ASAP7_75t_L g1193 ( 
.A1(n_934),
.A2(n_926),
.B(n_932),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_977),
.A2(n_464),
.B(n_455),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_931),
.A2(n_668),
.B(n_2),
.C(n_3),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_1029),
.B(n_84),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1001),
.B(n_1),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1089),
.A2(n_668),
.B(n_3),
.C(n_4),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_2),
.B(n_6),
.C(n_12),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1008),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1101),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1100),
.B(n_205),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1012),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_949),
.A2(n_198),
.B(n_192),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_R g1205 ( 
.A(n_990),
.B(n_191),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1102),
.B(n_1107),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1110),
.A2(n_16),
.B(n_18),
.C(n_20),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1100),
.B(n_22),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1076),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_946),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1067),
.B(n_190),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1078),
.A2(n_28),
.B(n_38),
.C(n_39),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_930),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_980),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_947),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1001),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1032),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_L g1218 ( 
.A1(n_977),
.A2(n_188),
.B(n_186),
.C(n_173),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_970),
.B(n_127),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1068),
.B(n_40),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_976),
.B(n_40),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1103),
.B(n_44),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_962),
.A2(n_154),
.B1(n_153),
.B2(n_152),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_953),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_999),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_941),
.A2(n_149),
.B(n_143),
.Y(n_1226)
);

NOR3xp33_ASAP7_75t_SL g1227 ( 
.A(n_999),
.B(n_45),
.C(n_49),
.Y(n_1227)
);

OAI21xp33_ASAP7_75t_SL g1228 ( 
.A1(n_941),
.A2(n_50),
.B(n_51),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_980),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1035),
.A2(n_137),
.B(n_136),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_990),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1077),
.B(n_53),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1072),
.B(n_123),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1039),
.A2(n_1065),
.B(n_1088),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1103),
.B(n_53),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1072),
.B(n_1094),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1084),
.A2(n_122),
.B(n_121),
.Y(n_1237)
);

AOI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_939),
.A2(n_55),
.B(n_58),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_926),
.A2(n_118),
.B(n_102),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_SL g1240 ( 
.A1(n_1087),
.A2(n_101),
.B(n_100),
.C(n_64),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1084),
.A2(n_60),
.B(n_61),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_948),
.B(n_64),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_979),
.B(n_65),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_948),
.B(n_66),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_930),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1038),
.A2(n_1034),
.B(n_1053),
.C(n_1046),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1079),
.A2(n_1105),
.B(n_1104),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_SL g1248 ( 
.A1(n_1093),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1095),
.A2(n_68),
.B(n_73),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_930),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1094),
.B(n_76),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_935),
.A2(n_76),
.B1(n_936),
.B2(n_1043),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_979),
.B(n_1016),
.Y(n_1253)
);

NOR3xp33_ASAP7_75t_SL g1254 ( 
.A(n_942),
.B(n_1056),
.C(n_1051),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1097),
.A2(n_1109),
.B(n_1082),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_979),
.B(n_1016),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1090),
.A2(n_1111),
.B(n_1061),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1018),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_935),
.A2(n_936),
.B1(n_1043),
.B2(n_1042),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1061),
.A2(n_1064),
.B(n_1048),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_955),
.A2(n_1037),
.B(n_973),
.C(n_1033),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1047),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1032),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_956),
.B(n_1007),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1024),
.A2(n_1005),
.B(n_987),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_964),
.B(n_1042),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_SL g1267 ( 
.A1(n_954),
.A2(n_1018),
.B1(n_964),
.B2(n_1042),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1018),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1234),
.A2(n_987),
.B(n_930),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1206),
.B(n_962),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1127),
.B(n_1166),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1125),
.A2(n_986),
.B(n_992),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1180),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1193),
.A2(n_1002),
.A3(n_1007),
.B(n_956),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1116),
.A2(n_942),
.B(n_954),
.C(n_966),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1112),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1170),
.A2(n_1252),
.B1(n_1195),
.B2(n_1128),
.C(n_1244),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1124),
.B(n_962),
.Y(n_1278)
);

AOI211x1_ASAP7_75t_L g1279 ( 
.A1(n_1164),
.A2(n_1096),
.B(n_1015),
.C(n_1013),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1136),
.A2(n_1050),
.B(n_993),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1124),
.B(n_962),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1164),
.B(n_962),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1231),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1224),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1173),
.A2(n_1108),
.B(n_982),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1156),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1149),
.B(n_1003),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1187),
.B(n_1229),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1255),
.A2(n_1019),
.B(n_1003),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1128),
.A2(n_988),
.A3(n_1014),
.B(n_960),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1185),
.B(n_1047),
.Y(n_1291)
);

NAND2x1_ASAP7_75t_L g1292 ( 
.A(n_1168),
.B(n_1003),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1246),
.A2(n_988),
.A3(n_1014),
.B(n_960),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1114),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1112),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1117),
.B(n_1002),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1134),
.B(n_972),
.Y(n_1297)
);

NOR2x1_ASAP7_75t_R g1298 ( 
.A(n_1123),
.B(n_1008),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1232),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1122),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1142),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1170),
.A2(n_961),
.A3(n_959),
.B(n_1009),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1131),
.A2(n_998),
.B(n_967),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1112),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1148),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1115),
.A2(n_1059),
.B(n_974),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1260),
.A2(n_1036),
.B(n_1069),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1252),
.A2(n_1019),
.B(n_1003),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1262),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1120),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1120),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1141),
.B(n_1045),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1187),
.B(n_954),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1168),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1120),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1118),
.A2(n_1049),
.B1(n_1019),
.B2(n_1004),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1177),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_1073),
.B(n_1069),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1147),
.B(n_1040),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1197),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1160),
.A2(n_995),
.B(n_1000),
.Y(n_1321)
);

OAI21xp33_ASAP7_75t_L g1322 ( 
.A1(n_1171),
.A2(n_1220),
.B(n_1221),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1118),
.A2(n_1049),
.B1(n_1066),
.B2(n_1063),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1119),
.A2(n_1054),
.B(n_1085),
.C(n_1057),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1257),
.A2(n_1054),
.B(n_1098),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1121),
.A2(n_1045),
.B1(n_1057),
.B2(n_1062),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1191),
.B(n_1062),
.Y(n_1327)
);

AO32x2_ASAP7_75t_L g1328 ( 
.A1(n_1209),
.A2(n_1098),
.A3(n_1259),
.B1(n_1216),
.B2(n_1178),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1192),
.A2(n_1098),
.B(n_1132),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1144),
.A2(n_1145),
.B(n_1202),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1242),
.A2(n_1098),
.B(n_1126),
.C(n_1261),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1202),
.A2(n_1264),
.B(n_1259),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1146),
.B(n_1267),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1129),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1157),
.B(n_1158),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1266),
.B(n_1254),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1181),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1161),
.B(n_1172),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1186),
.A2(n_1237),
.B(n_1143),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1210),
.B(n_1215),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1138),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1251),
.B(n_1238),
.C(n_1249),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1169),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1228),
.A2(n_1218),
.B(n_1226),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1138),
.A2(n_1184),
.B1(n_1175),
.B2(n_1153),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1208),
.A2(n_1222),
.B(n_1235),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1129),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1239),
.A2(n_1190),
.B(n_1256),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1183),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1129),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1139),
.B(n_1217),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1146),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1263),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1198),
.A2(n_1201),
.A3(n_1207),
.B(n_1199),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1241),
.A2(n_1212),
.A3(n_1178),
.B(n_1204),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1253),
.A2(n_1230),
.B(n_1155),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1167),
.B(n_1236),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1135),
.B(n_1152),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1138),
.A2(n_1175),
.B(n_1184),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1174),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1133),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1243),
.Y(n_1362)
);

NAND2x1_ASAP7_75t_L g1363 ( 
.A(n_1146),
.B(n_1200),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_SL g1364 ( 
.A1(n_1151),
.A2(n_1240),
.B(n_1211),
.C(n_1233),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1154),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1138),
.A2(n_1175),
.B(n_1184),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1154),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1174),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1140),
.B(n_1130),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1175),
.B(n_1184),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1182),
.B(n_1245),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1248),
.A2(n_1150),
.B(n_1238),
.C(n_1137),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1174),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1223),
.A2(n_1225),
.B(n_1165),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1216),
.A2(n_1205),
.B1(n_1179),
.B2(n_1196),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1203),
.A2(n_1189),
.B(n_1113),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1219),
.B(n_1250),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1209),
.A2(n_1188),
.B(n_1159),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1188),
.A2(n_1159),
.B(n_1268),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1219),
.A2(n_1213),
.B(n_1250),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1258),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1227),
.A2(n_1213),
.B(n_1250),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1163),
.A2(n_1193),
.A3(n_1128),
.B(n_1246),
.Y(n_1383)
);

AOI221x1_ASAP7_75t_L g1384 ( 
.A1(n_1213),
.A2(n_1170),
.B1(n_1252),
.B2(n_1195),
.C(n_945),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1163),
.B(n_1214),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1247),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1265),
.A2(n_1173),
.B(n_1176),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1162),
.B(n_971),
.Y(n_1388)
);

NOR3xp33_ASAP7_75t_L g1389 ( 
.A(n_1137),
.B(n_760),
.C(n_697),
.Y(n_1389)
);

NAND3x1_ASAP7_75t_L g1390 ( 
.A(n_1232),
.B(n_677),
.C(n_717),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1180),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1125),
.A2(n_984),
.B(n_1136),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1127),
.B(n_892),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1125),
.A2(n_984),
.B(n_1136),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1112),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1114),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_SL g1398 ( 
.A1(n_1239),
.A2(n_1226),
.B(n_1193),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1123),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1180),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1247),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1116),
.A2(n_760),
.B(n_759),
.C(n_826),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1125),
.A2(n_934),
.B(n_1116),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1116),
.A2(n_760),
.B1(n_826),
.B2(n_697),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1252),
.A2(n_984),
.B(n_895),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1265),
.A2(n_1173),
.B(n_1176),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1193),
.A2(n_1246),
.B(n_1125),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1180),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1193),
.A2(n_1246),
.B(n_1125),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1247),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1125),
.A2(n_934),
.B(n_1116),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1231),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1114),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1138),
.B(n_1175),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1180),
.Y(n_1419)
);

OAI22x1_ASAP7_75t_L g1420 ( 
.A1(n_1242),
.A2(n_677),
.B1(n_944),
.B2(n_664),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1247),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1206),
.B(n_1127),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1112),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1180),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1247),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1127),
.B(n_940),
.Y(n_1428)
);

AO22x2_ASAP7_75t_L g1429 ( 
.A1(n_1170),
.A2(n_1252),
.B1(n_1216),
.B2(n_1091),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1369),
.B(n_1299),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1404),
.A2(n_1369),
.B1(n_1390),
.B2(n_1375),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1386),
.A2(n_1411),
.B(n_1401),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1313),
.B(n_1377),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1423),
.A2(n_1427),
.B(n_1394),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

AOI222xp33_ASAP7_75t_L g1436 ( 
.A1(n_1420),
.A2(n_1322),
.B1(n_1429),
.B2(n_1393),
.C1(n_1392),
.C2(n_1394),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1314),
.B(n_1352),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1294),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1285),
.A2(n_1406),
.B(n_1387),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1309),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1389),
.A2(n_1357),
.B1(n_1336),
.B2(n_1291),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_SL g1442 ( 
.A1(n_1331),
.A2(n_1281),
.B(n_1278),
.C(n_1270),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1392),
.A2(n_1402),
.B(n_1405),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1270),
.B(n_1275),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1398),
.A2(n_1344),
.B(n_1403),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1304),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1271),
.B(n_1362),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1313),
.B(n_1377),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1307),
.A2(n_1289),
.B(n_1356),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1339),
.A2(n_1413),
.B(n_1318),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1346),
.A2(n_1321),
.B(n_1282),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1332),
.A2(n_1348),
.B(n_1272),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1340),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1272),
.A2(n_1280),
.B(n_1303),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1282),
.A2(n_1316),
.B(n_1323),
.Y(n_1456)
);

INVxp67_ASAP7_75t_SL g1457 ( 
.A(n_1316),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1280),
.A2(n_1308),
.B(n_1324),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1342),
.A2(n_1344),
.B(n_1378),
.C(n_1426),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1315),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1359),
.A2(n_1366),
.B(n_1277),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1293),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1278),
.A2(n_1281),
.B(n_1376),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1293),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1359),
.A2(n_1366),
.B(n_1380),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1333),
.B(n_1380),
.Y(n_1467)
);

OAI211xp5_ASAP7_75t_L g1468 ( 
.A1(n_1384),
.A2(n_1372),
.B(n_1414),
.C(n_1424),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1352),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1374),
.A2(n_1379),
.B(n_1367),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1412),
.B(n_1414),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1323),
.A2(n_1365),
.A3(n_1345),
.B(n_1358),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1286),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1294),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1276),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1358),
.A2(n_1296),
.A3(n_1319),
.B(n_1297),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1284),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1429),
.A2(n_1273),
.B1(n_1391),
.B2(n_1400),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1333),
.B(n_1341),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1407),
.A2(n_1410),
.B(n_1296),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1407),
.A2(n_1410),
.B(n_1297),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1353),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1347),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1314),
.B(n_1341),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1335),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1409),
.A2(n_1419),
.B(n_1424),
.C(n_1422),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1412),
.B(n_1422),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1417),
.A2(n_1421),
.B1(n_1333),
.B2(n_1397),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1361),
.A2(n_1417),
.B1(n_1421),
.B2(n_1416),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1335),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1312),
.A2(n_1319),
.B(n_1418),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1312),
.A2(n_1418),
.B(n_1370),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1343),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1370),
.A2(n_1326),
.B(n_1351),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1388),
.B(n_1327),
.Y(n_1495)
);

CKINVDCx6p67_ASAP7_75t_R g1496 ( 
.A(n_1276),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1306),
.A2(n_1364),
.B(n_1371),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1351),
.A2(n_1371),
.B(n_1300),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1302),
.Y(n_1499)
);

NAND2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1314),
.B(n_1363),
.Y(n_1500)
);

AO31x2_ASAP7_75t_L g1501 ( 
.A1(n_1290),
.A2(n_1383),
.A3(n_1337),
.B(n_1317),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1292),
.A2(n_1305),
.B(n_1301),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1360),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1382),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1320),
.A2(n_1428),
.B1(n_1381),
.B2(n_1287),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1382),
.Y(n_1506)
);

AO32x2_ASAP7_75t_L g1507 ( 
.A1(n_1290),
.A2(n_1328),
.A3(n_1274),
.B1(n_1383),
.B2(n_1354),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1288),
.B(n_1373),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1274),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1306),
.A2(n_1279),
.B(n_1355),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1355),
.A2(n_1354),
.B(n_1328),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1354),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1288),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1349),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1320),
.B(n_1350),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1328),
.A2(n_1334),
.B(n_1295),
.C(n_1368),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1355),
.A2(n_1314),
.B(n_1385),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1385),
.A2(n_1276),
.B(n_1425),
.Y(n_1518)
);

AOI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1385),
.A2(n_1283),
.B(n_1415),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1310),
.B(n_1311),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1311),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1395),
.Y(n_1522)
);

AO31x2_ASAP7_75t_L g1523 ( 
.A1(n_1395),
.A2(n_1277),
.A3(n_1193),
.B(n_1386),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1395),
.B(n_1425),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1425),
.A2(n_1401),
.B(n_1386),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1298),
.A2(n_1401),
.B(n_1386),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1393),
.B(n_1396),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1308),
.B(n_1405),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1293),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1293),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1293),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1314),
.B(n_1138),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1308),
.B(n_1405),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1293),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1389),
.A2(n_760),
.B(n_1402),
.C(n_759),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1386),
.A2(n_1411),
.B(n_1401),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1399),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1393),
.B(n_1396),
.Y(n_1538)
);

NAND2x1_ASAP7_75t_L g1539 ( 
.A(n_1308),
.B(n_1168),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1402),
.A2(n_760),
.B(n_759),
.Y(n_1540)
);

CKINVDCx11_ASAP7_75t_R g1541 ( 
.A(n_1320),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1338),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1329),
.A2(n_1330),
.B(n_1387),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_SL g1545 ( 
.A1(n_1275),
.A2(n_1270),
.B(n_1346),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1402),
.A2(n_760),
.B(n_759),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1314),
.B(n_1138),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1393),
.B(n_1396),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1404),
.A2(n_1299),
.B1(n_760),
.B2(n_826),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1402),
.A2(n_760),
.B(n_759),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1392),
.A2(n_1394),
.B(n_984),
.C(n_759),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1293),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1329),
.A2(n_1269),
.B(n_1325),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1393),
.B(n_1271),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1293),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1302),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1393),
.B(n_1271),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_R g1558 ( 
.A(n_1399),
.B(n_690),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_L g1559 ( 
.A(n_1399),
.B(n_1123),
.Y(n_1559)
);

AND2x6_ASAP7_75t_L g1560 ( 
.A(n_1341),
.B(n_1278),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1369),
.B(n_760),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1293),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1404),
.B(n_760),
.C(n_1389),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1404),
.A2(n_1277),
.B1(n_677),
.B2(n_731),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1386),
.A2(n_1411),
.B(n_1401),
.Y(n_1565)
);

AO31x2_ASAP7_75t_L g1566 ( 
.A1(n_1277),
.A2(n_1193),
.A3(n_1401),
.B(n_1386),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1293),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1304),
.Y(n_1568)
);

AOI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1403),
.A2(n_1116),
.B(n_934),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1314),
.B(n_1138),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1294),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_SL g1572 ( 
.A1(n_1331),
.A2(n_945),
.B(n_1195),
.C(n_1116),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1386),
.A2(n_1411),
.B(n_1401),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1286),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1313),
.B(n_1377),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1352),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1329),
.A2(n_1330),
.B(n_1387),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1495),
.B(n_1527),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1535),
.A2(n_1550),
.B(n_1546),
.C(n_1540),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1563),
.A2(n_1441),
.B1(n_1561),
.B2(n_1564),
.Y(n_1581)
);

A2O1A1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1561),
.A2(n_1458),
.B(n_1551),
.C(n_1443),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1450),
.B(n_1461),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1489),
.B(n_1433),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1433),
.B(n_1448),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1564),
.A2(n_1431),
.B(n_1549),
.C(n_1551),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1470),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1434),
.A2(n_1462),
.B(n_1573),
.Y(n_1588)
);

CKINVDCx6p67_ASAP7_75t_R g1589 ( 
.A(n_1514),
.Y(n_1589)
);

O2A1O1Ixp5_ASAP7_75t_L g1590 ( 
.A1(n_1444),
.A2(n_1468),
.B(n_1459),
.C(n_1464),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1433),
.B(n_1448),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1538),
.B(n_1548),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1446),
.Y(n_1593)
);

O2A1O1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1572),
.A2(n_1486),
.B(n_1444),
.C(n_1459),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1505),
.A2(n_1430),
.B1(n_1447),
.B2(n_1478),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1522),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1510),
.A2(n_1453),
.B(n_1455),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1471),
.B(n_1543),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1467),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1474),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1487),
.B(n_1447),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1488),
.B(n_1438),
.Y(n_1602)
);

OAI211xp5_ASAP7_75t_L g1603 ( 
.A1(n_1436),
.A2(n_1572),
.B(n_1430),
.C(n_1505),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1478),
.A2(n_1493),
.B1(n_1486),
.B2(n_1533),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1571),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1435),
.B(n_1454),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1575),
.B(n_1513),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1528),
.A2(n_1533),
.B1(n_1457),
.B2(n_1542),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1432),
.A2(n_1536),
.B(n_1565),
.Y(n_1609)
);

OA21x2_ASAP7_75t_L g1610 ( 
.A1(n_1480),
.A2(n_1481),
.B(n_1451),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1482),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1432),
.A2(n_1536),
.B(n_1565),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1479),
.A2(n_1515),
.B1(n_1485),
.B2(n_1490),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1498),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1508),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1503),
.B(n_1498),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1565),
.A2(n_1526),
.B(n_1525),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1479),
.A2(n_1515),
.B1(n_1574),
.B2(n_1473),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1470),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1483),
.Y(n_1620)
);

A2O1A1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1516),
.A2(n_1511),
.B(n_1539),
.C(n_1517),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1498),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1541),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1476),
.B(n_1472),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1442),
.A2(n_1545),
.B(n_1466),
.C(n_1518),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1476),
.B(n_1472),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1520),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1442),
.A2(n_1516),
.B(n_1521),
.C(n_1504),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1519),
.A2(n_1514),
.B1(n_1460),
.B2(n_1568),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1520),
.B(n_1524),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1512),
.A2(n_1556),
.B1(n_1499),
.B2(n_1445),
.C(n_1506),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1446),
.A2(n_1460),
.B1(n_1568),
.B2(n_1469),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1501),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1476),
.B(n_1472),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1532),
.A2(n_1547),
.B(n_1570),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1532),
.A2(n_1547),
.B(n_1570),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1440),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_1440),
.Y(n_1638)
);

NOR2xp67_ASAP7_75t_L g1639 ( 
.A(n_1537),
.B(n_1559),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1475),
.B(n_1469),
.Y(n_1640)
);

BUFx8_ASAP7_75t_SL g1641 ( 
.A(n_1537),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1470),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1497),
.A2(n_1576),
.B(n_1500),
.C(n_1484),
.Y(n_1643)
);

O2A1O1Ixp5_ASAP7_75t_L g1644 ( 
.A1(n_1456),
.A2(n_1569),
.B(n_1452),
.C(n_1552),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1500),
.A2(n_1437),
.B1(n_1496),
.B2(n_1484),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1523),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1472),
.B(n_1560),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1507),
.B(n_1523),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1560),
.B(n_1523),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1507),
.B(n_1566),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1492),
.B(n_1560),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_1522),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1439),
.A2(n_1449),
.B(n_1577),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1558),
.A2(n_1534),
.B(n_1463),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1463),
.A2(n_1529),
.B1(n_1465),
.B2(n_1555),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1494),
.A2(n_1491),
.B(n_1502),
.C(n_1465),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1560),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1529),
.A2(n_1552),
.B1(n_1567),
.B2(n_1562),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1530),
.A2(n_1567),
.B1(n_1531),
.B2(n_1509),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1577),
.A2(n_1544),
.B(n_1553),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1566),
.A2(n_1551),
.B(n_1252),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1512),
.B(n_1464),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1663)
);

AND2x2_ASAP7_75t_SL g1664 ( 
.A(n_1467),
.B(n_1389),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1467),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1564),
.A2(n_1561),
.B1(n_666),
.B2(n_1563),
.C(n_760),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1563),
.A2(n_1375),
.B1(n_1404),
.B2(n_1441),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1551),
.A2(n_1252),
.B(n_1493),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1477),
.Y(n_1669)
);

O2A1O1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1535),
.A2(n_1546),
.B(n_1550),
.C(n_1540),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1495),
.B(n_1527),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1467),
.B(n_1479),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1561),
.A2(n_1540),
.B(n_1550),
.C(n_1546),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1561),
.B(n_1450),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1561),
.B(n_1450),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1434),
.A2(n_1462),
.B(n_1573),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1493),
.Y(n_1678)
);

AOI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1563),
.A2(n_1564),
.B(n_1389),
.C(n_760),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1540),
.A2(n_1550),
.B(n_1546),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_SL g1681 ( 
.A1(n_1540),
.A2(n_1546),
.B(n_1550),
.C(n_1535),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1561),
.B(n_1450),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1563),
.A2(n_1375),
.B1(n_1404),
.B2(n_1441),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1563),
.B(n_1535),
.C(n_760),
.Y(n_1685)
);

OA22x2_ASAP7_75t_L g1686 ( 
.A1(n_1441),
.A2(n_1420),
.B1(n_1431),
.B2(n_1404),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1441),
.A2(n_571),
.B1(n_1431),
.B2(n_1561),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1477),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1563),
.A2(n_1375),
.B1(n_1404),
.B2(n_1441),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1551),
.A2(n_1252),
.B(n_1493),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1477),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1563),
.A2(n_1375),
.B1(n_1404),
.B2(n_1441),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1680),
.B(n_1661),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1616),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1674),
.A2(n_1670),
.B(n_1579),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1647),
.B(n_1624),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1626),
.B(n_1634),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1614),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1649),
.B(n_1662),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1609),
.A2(n_1612),
.B(n_1617),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1622),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1599),
.B(n_1665),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1675),
.B(n_1676),
.Y(n_1703)
);

NAND2x1p5_ASAP7_75t_L g1704 ( 
.A(n_1657),
.B(n_1664),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1633),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1665),
.B(n_1673),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1581),
.A2(n_1666),
.B1(n_1687),
.B2(n_1692),
.C(n_1667),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1673),
.B(n_1648),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1691),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1684),
.A2(n_1689),
.B1(n_1686),
.B2(n_1685),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1686),
.A2(n_1679),
.B1(n_1603),
.B2(n_1595),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1669),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1674),
.A2(n_1681),
.B(n_1582),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1673),
.B(n_1648),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1688),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1611),
.Y(n_1717)
);

AO21x2_ASAP7_75t_L g1718 ( 
.A1(n_1656),
.A2(n_1621),
.B(n_1582),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1654),
.B(n_1643),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1650),
.B(n_1585),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1644),
.A2(n_1590),
.B(n_1631),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1650),
.B(n_1591),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1664),
.A2(n_1584),
.B1(n_1629),
.B2(n_1602),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1587),
.A2(n_1642),
.B(n_1619),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1678),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1683),
.B(n_1592),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1613),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1620),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1610),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_SL g1730 ( 
.A(n_1604),
.B(n_1608),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1655),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1598),
.B(n_1646),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1658),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1660),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1659),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1606),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1660),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1583),
.B(n_1601),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1615),
.B(n_1671),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1628),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1607),
.B(n_1630),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1593),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1698),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1696),
.B(n_1677),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1701),
.Y(n_1745)
);

INVx3_ASAP7_75t_SL g1746 ( 
.A(n_1693),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1713),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1708),
.B(n_1715),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1707),
.A2(n_1586),
.B(n_1594),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1734),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1713),
.B(n_1640),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1720),
.B(n_1588),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1713),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1696),
.B(n_1597),
.Y(n_1755)
);

AO21x2_ASAP7_75t_L g1756 ( 
.A1(n_1700),
.A2(n_1625),
.B(n_1668),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1705),
.Y(n_1757)
);

AO21x2_ASAP7_75t_L g1758 ( 
.A1(n_1700),
.A2(n_1690),
.B(n_1668),
.Y(n_1758)
);

NAND2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1710),
.B(n_1596),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1694),
.B(n_1578),
.Y(n_1760)
);

OR2x6_ASAP7_75t_SL g1761 ( 
.A(n_1699),
.B(n_1618),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1707),
.A2(n_1580),
.B1(n_1663),
.B2(n_1682),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1722),
.B(n_1653),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1724),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1711),
.A2(n_1690),
.B1(n_1600),
.B2(n_1672),
.C(n_1605),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1694),
.B(n_1736),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1724),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1711),
.A2(n_1623),
.B1(n_1639),
.B2(n_1654),
.C(n_1645),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1699),
.B(n_1627),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1693),
.B(n_1593),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1750),
.A2(n_1729),
.B(n_1737),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1752),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1743),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1759),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1769),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1749),
.A2(n_1695),
.B1(n_1714),
.B2(n_1723),
.C(n_1693),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1760),
.B(n_1638),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1749),
.A2(n_1695),
.B1(n_1714),
.B2(n_1693),
.C(n_1704),
.Y(n_1778)
);

AOI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1768),
.A2(n_1703),
.B(n_1740),
.C(n_1726),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1759),
.A2(n_1693),
.B1(n_1704),
.B2(n_1718),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1743),
.Y(n_1781)
);

OAI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1765),
.A2(n_1740),
.B(n_1721),
.C(n_1719),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1768),
.A2(n_1704),
.B1(n_1718),
.B2(n_1727),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1760),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1755),
.B(n_1732),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1765),
.B(n_1721),
.C(n_1719),
.Y(n_1786)
);

NAND2xp33_ASAP7_75t_R g1787 ( 
.A(n_1766),
.B(n_1738),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1761),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1743),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1745),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1758),
.A2(n_1718),
.B1(n_1741),
.B2(n_1706),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1754),
.B(n_1747),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1745),
.Y(n_1793)
);

AOI31xp33_ASAP7_75t_L g1794 ( 
.A1(n_1762),
.A2(n_1738),
.A3(n_1632),
.B(n_1736),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1766),
.B(n_1725),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1769),
.B(n_1739),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1769),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1755),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1758),
.A2(n_1730),
.B(n_1636),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1750),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1748),
.B(n_1702),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1739),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1758),
.A2(n_1741),
.B1(n_1728),
.B2(n_1721),
.Y(n_1803)
);

OAI21xp33_ASAP7_75t_SL g1804 ( 
.A1(n_1770),
.A2(n_1716),
.B(n_1712),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1762),
.B(n_1721),
.C(n_1731),
.Y(n_1805)
);

NAND4xp25_ASAP7_75t_L g1806 ( 
.A(n_1744),
.B(n_1732),
.C(n_1697),
.D(n_1731),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1751),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1744),
.B(n_1721),
.C(n_1735),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1756),
.A2(n_1709),
.B1(n_1717),
.B2(n_1716),
.C(n_1712),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1757),
.Y(n_1810)
);

AO21x1_ASAP7_75t_SL g1811 ( 
.A1(n_1757),
.A2(n_1733),
.B(n_1735),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1746),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1770),
.A2(n_1728),
.B1(n_1742),
.B2(n_1589),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1761),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1773),
.Y(n_1815)
);

OR2x6_ASAP7_75t_L g1816 ( 
.A(n_1799),
.B(n_1747),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1771),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1771),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1771),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1773),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1792),
.B(n_1763),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1786),
.A2(n_1756),
.B(n_1596),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1781),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1804),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1790),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1812),
.Y(n_1826)
);

OA21x2_ASAP7_75t_L g1827 ( 
.A1(n_1808),
.A2(n_1767),
.B(n_1764),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1812),
.Y(n_1828)
);

CKINVDCx20_ASAP7_75t_R g1829 ( 
.A(n_1774),
.Y(n_1829)
);

OA21x2_ASAP7_75t_L g1830 ( 
.A1(n_1809),
.A2(n_1767),
.B(n_1764),
.Y(n_1830)
);

OAI21xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1776),
.A2(n_1778),
.B(n_1805),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1800),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1807),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1785),
.B(n_1755),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1789),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1811),
.Y(n_1836)
);

INVx4_ASAP7_75t_SL g1837 ( 
.A(n_1812),
.Y(n_1837)
);

INVx4_ASAP7_75t_SL g1838 ( 
.A(n_1812),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1793),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1810),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1792),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1828),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1829),
.B(n_1641),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1826),
.B(n_1772),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1820),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1820),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

INVx3_ASAP7_75t_R g1848 ( 
.A(n_1828),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1825),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1825),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1833),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1834),
.B(n_1806),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1826),
.B(n_1772),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1831),
.A2(n_1782),
.B(n_1783),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1826),
.B(n_1814),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1831),
.B(n_1784),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1833),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1817),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1815),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1826),
.B(n_1792),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1837),
.B(n_1812),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1835),
.B(n_1798),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1835),
.B(n_1797),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1828),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1837),
.B(n_1754),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1839),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1815),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1834),
.B(n_1785),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1836),
.B(n_1801),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1839),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1834),
.B(n_1824),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1822),
.B(n_1788),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1840),
.B(n_1788),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1754),
.Y(n_1874)
);

NAND2x1_ASAP7_75t_SL g1875 ( 
.A(n_1827),
.B(n_1830),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1837),
.B(n_1775),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1817),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1817),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1837),
.B(n_1794),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1824),
.B(n_1802),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1836),
.B(n_1801),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1824),
.B(n_1796),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1837),
.B(n_1811),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1840),
.B(n_1795),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1754),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1838),
.B(n_1754),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1838),
.B(n_1754),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1875),
.Y(n_1888)
);

INVxp67_ASAP7_75t_SL g1889 ( 
.A(n_1871),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1854),
.B(n_1779),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1854),
.B(n_1777),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1875),
.Y(n_1894)
);

AND2x2_ASAP7_75t_SL g1895 ( 
.A(n_1856),
.B(n_1596),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1856),
.B(n_1748),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1866),
.Y(n_1897)
);

OAI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1872),
.A2(n_1787),
.B1(n_1774),
.B2(n_1746),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1870),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1843),
.B(n_1829),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1859),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1859),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1867),
.Y(n_1904)
);

NOR2xp67_ASAP7_75t_L g1905 ( 
.A(n_1883),
.B(n_1841),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1882),
.B(n_1815),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1855),
.B(n_1748),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1855),
.B(n_1838),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1883),
.B(n_1838),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1861),
.B(n_1841),
.Y(n_1910)
);

OAI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1879),
.A2(n_1746),
.B1(n_1816),
.B2(n_1841),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1873),
.A2(n_1816),
.B(n_1827),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1873),
.B(n_1821),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1860),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1847),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1842),
.B(n_1821),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1845),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1857),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1847),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1882),
.B(n_1823),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1869),
.B(n_1881),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1871),
.B(n_1823),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1852),
.B(n_1880),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1865),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1895),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1895),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1889),
.Y(n_1927)
);

INVx1_ASAP7_75t_SL g1928 ( 
.A(n_1923),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1922),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1922),
.Y(n_1930)
);

INVx3_ASAP7_75t_SL g1931 ( 
.A(n_1890),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1923),
.B(n_1842),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1890),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1921),
.B(n_1909),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1890),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1891),
.B(n_1869),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1921),
.B(n_1881),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1906),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1906),
.Y(n_1939)
);

AO22x1_ASAP7_75t_L g1940 ( 
.A1(n_1892),
.A2(n_1864),
.B1(n_1848),
.B2(n_1596),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1909),
.B(n_1860),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1902),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1898),
.A2(n_1913),
.B1(n_1896),
.B2(n_1911),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1893),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1903),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1893),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1893),
.B(n_1844),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1900),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1900),
.B(n_1864),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1904),
.Y(n_1950)
);

AO21x2_ASAP7_75t_L g1951 ( 
.A1(n_1888),
.A2(n_1848),
.B(n_1846),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1900),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1927),
.A2(n_1894),
.B(n_1888),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1932),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1940),
.A2(n_1901),
.B(n_1912),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1944),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1944),
.B(n_1934),
.Y(n_1957)
);

AOI222xp33_ASAP7_75t_L g1958 ( 
.A1(n_1928),
.A2(n_1918),
.B1(n_1917),
.B2(n_1897),
.C1(n_1899),
.C2(n_1894),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1932),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1943),
.A2(n_1908),
.B1(n_1914),
.B2(n_1905),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1937),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1940),
.A2(n_1918),
.B(n_1917),
.Y(n_1962)
);

INVxp67_ASAP7_75t_L g1963 ( 
.A(n_1934),
.Y(n_1963)
);

OAI322xp33_ASAP7_75t_L g1964 ( 
.A1(n_1925),
.A2(n_1897),
.A3(n_1899),
.B1(n_1914),
.B2(n_1920),
.C1(n_1916),
.C2(n_1852),
.Y(n_1964)
);

NAND3xp33_ASAP7_75t_L g1965 ( 
.A(n_1927),
.B(n_1910),
.C(n_1920),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1937),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1926),
.A2(n_1756),
.B1(n_1780),
.B2(n_1910),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1936),
.A2(n_1887),
.B(n_1886),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1929),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1929),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1933),
.B(n_1907),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1935),
.A2(n_1849),
.B1(n_1851),
.B2(n_1846),
.C(n_1850),
.Y(n_1972)
);

AOI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1946),
.A2(n_1924),
.B(n_1876),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1931),
.A2(n_1880),
.B1(n_1803),
.B2(n_1791),
.Y(n_1974)
);

NOR2x1_ASAP7_75t_L g1975 ( 
.A(n_1953),
.B(n_1951),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1958),
.B(n_1930),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1961),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1966),
.B(n_1930),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1957),
.B(n_1948),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1954),
.B(n_1938),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1957),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1963),
.B(n_1947),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1956),
.B(n_1947),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1959),
.B(n_1941),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1964),
.B(n_1952),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1971),
.B(n_1941),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1973),
.B(n_1931),
.Y(n_1987)
);

INVx2_ASAP7_75t_SL g1988 ( 
.A(n_1953),
.Y(n_1988)
);

AOI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1975),
.A2(n_1962),
.B(n_1955),
.Y(n_1989)
);

AOI322xp5_ASAP7_75t_L g1990 ( 
.A1(n_1985),
.A2(n_1972),
.A3(n_1967),
.B1(n_1970),
.B2(n_1969),
.C1(n_1938),
.C2(n_1939),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1981),
.B(n_1983),
.Y(n_1991)
);

AOI211xp5_ASAP7_75t_SL g1992 ( 
.A1(n_1976),
.A2(n_1960),
.B(n_1974),
.C(n_1949),
.Y(n_1992)
);

A2O1A1Ixp33_ASAP7_75t_L g1993 ( 
.A1(n_1976),
.A2(n_1967),
.B(n_1965),
.C(n_1968),
.Y(n_1993)
);

NAND3xp33_ASAP7_75t_L g1994 ( 
.A(n_1987),
.B(n_1949),
.C(n_1939),
.Y(n_1994)
);

OAI33xp33_ASAP7_75t_L g1995 ( 
.A1(n_1978),
.A2(n_1942),
.A3(n_1950),
.B1(n_1945),
.B2(n_1851),
.B3(n_1849),
.Y(n_1995)
);

NAND4xp25_ASAP7_75t_L g1996 ( 
.A(n_1979),
.B(n_1949),
.C(n_1950),
.D(n_1942),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1984),
.B(n_1931),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1983),
.B(n_1986),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_L g1999 ( 
.A(n_1980),
.B(n_1949),
.C(n_1945),
.Y(n_1999)
);

OAI221xp5_ASAP7_75t_SL g2000 ( 
.A1(n_1988),
.A2(n_1924),
.B1(n_1816),
.B2(n_1951),
.C(n_1813),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_L g2001 ( 
.A1(n_1980),
.A2(n_1951),
.B1(n_1924),
.B2(n_1850),
.C(n_1915),
.Y(n_2001)
);

AOI222xp33_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_1993),
.B1(n_1994),
.B2(n_1999),
.C1(n_1995),
.C2(n_1991),
.Y(n_2002)
);

AOI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_2000),
.A2(n_1977),
.B1(n_1982),
.B2(n_1978),
.C(n_1919),
.Y(n_2003)
);

NOR2x1_ASAP7_75t_L g2004 ( 
.A(n_1998),
.B(n_1652),
.Y(n_2004)
);

NOR3x1_ASAP7_75t_L g2005 ( 
.A(n_1996),
.B(n_1863),
.C(n_1862),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1992),
.A2(n_1919),
.B(n_1915),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1997),
.B(n_1844),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1990),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_SL g2009 ( 
.A1(n_1989),
.A2(n_1858),
.B(n_1847),
.C(n_1877),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_2004),
.B(n_1865),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_2006),
.B(n_1652),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_2007),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_2008),
.B(n_1853),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2005),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2003),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2002),
.Y(n_2016)
);

NOR2xp67_ASAP7_75t_L g2017 ( 
.A(n_2009),
.B(n_1865),
.Y(n_2017)
);

AOI322xp5_ASAP7_75t_L g2018 ( 
.A1(n_2016),
.A2(n_1819),
.A3(n_1878),
.B1(n_1877),
.B2(n_1858),
.C1(n_1874),
.C2(n_1885),
.Y(n_2018)
);

CKINVDCx16_ASAP7_75t_R g2019 ( 
.A(n_2013),
.Y(n_2019)
);

AND2x2_ASAP7_75t_SL g2020 ( 
.A(n_2012),
.B(n_1641),
.Y(n_2020)
);

NAND4xp75_ASAP7_75t_L g2021 ( 
.A(n_2011),
.B(n_1887),
.C(n_1886),
.D(n_1827),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_2010),
.A2(n_1637),
.B(n_1865),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_2015),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2019),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2020),
.B(n_2014),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_2021),
.Y(n_2026)
);

AND2x2_ASAP7_75t_SL g2027 ( 
.A(n_2024),
.B(n_2023),
.Y(n_2027)
);

AOI322xp5_ASAP7_75t_L g2028 ( 
.A1(n_2027),
.A2(n_2025),
.A3(n_2026),
.B1(n_2022),
.B2(n_2017),
.C1(n_2018),
.C2(n_1858),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_2028),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2028),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2030),
.A2(n_2025),
.B1(n_1637),
.B2(n_1877),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2029),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_SL g2033 ( 
.A1(n_2032),
.A2(n_1589),
.B1(n_1885),
.B2(n_1874),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_2031),
.A2(n_1878),
.B1(n_1863),
.B2(n_1867),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_2033),
.A2(n_1878),
.B1(n_1885),
.B2(n_1874),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_SL g2036 ( 
.A1(n_2035),
.A2(n_2034),
.B1(n_1885),
.B2(n_1874),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_2036),
.B(n_1862),
.Y(n_2037)
);

OAI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_2037),
.A2(n_1884),
.B(n_1853),
.Y(n_2038)
);

AOI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_2038),
.A2(n_1819),
.B1(n_1884),
.B2(n_1818),
.C(n_1832),
.Y(n_2039)
);

AOI211xp5_ASAP7_75t_L g2040 ( 
.A1(n_2039),
.A2(n_1635),
.B(n_1868),
.C(n_1818),
.Y(n_2040)
);


endmodule