module fake_jpeg_2788_n_9 (n_0, n_1, n_9);

input n_0;
input n_1;

output n_9;

wire n_3;
wire n_2;
wire n_4;
wire n_8;
wire n_6;
wire n_5;
wire n_7;

CKINVDCx16_ASAP7_75t_R g2 ( 
.A(n_1),
.Y(n_2)
);

INVx4_ASAP7_75t_L g3 ( 
.A(n_0),
.Y(n_3)
);

BUFx2_ASAP7_75t_L g4 ( 
.A(n_3),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_4),
.Y(n_5)
);

AOI22xp33_ASAP7_75t_L g6 ( 
.A1(n_5),
.A2(n_3),
.B1(n_2),
.B2(n_0),
.Y(n_6)
);

OAI21x1_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_2),
.B(n_3),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_7),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);


endmodule