module fake_netlist_1_6525_n_686 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_686);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_686;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_76), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_72), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_59), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_55), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_48), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_60), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_57), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_20), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_66), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_71), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_56), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_62), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_17), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_31), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_73), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_20), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_67), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_32), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_34), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_80), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_49), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_11), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_45), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_23), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_50), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_53), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_42), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_51), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_38), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_64), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
INVxp33_ASAP7_75t_SL g126 ( .A(n_41), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_27), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_16), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_125), .B(n_1), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_94), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_125), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_112), .Y(n_137) );
NAND2xp33_ASAP7_75t_R g138 ( .A(n_105), .B(n_25), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_102), .B(n_1), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_92), .B(n_2), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_90), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_115), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_106), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_90), .Y(n_146) );
NOR2xp33_ASAP7_75t_R g147 ( .A(n_83), .B(n_30), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_120), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_122), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_117), .B(n_3), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_115), .B(n_3), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_126), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_90), .B(n_4), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
NOR2xp33_ASAP7_75t_R g157 ( .A(n_93), .B(n_33), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_117), .B(n_4), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_85), .B(n_35), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_128), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_106), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_124), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_86), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_81), .B(n_28), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_86), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_89), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_81), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_88), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_88), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_85), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_87), .B(n_5), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_130), .B(n_121), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_160), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_161), .B(n_103), .Y(n_176) );
INVx8_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_172), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_136), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_172), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_161), .A2(n_129), .B1(n_87), .B2(n_110), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_130), .B(n_114), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_155), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_131), .Y(n_189) );
NOR2x1p5_ASAP7_75t_L g190 ( .A(n_135), .B(n_129), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_130), .B(n_110), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_153), .B(n_127), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_155), .B(n_109), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_134), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVxp67_ASAP7_75t_SL g201 ( .A(n_169), .Y(n_201) );
INVxp33_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
NAND3xp33_ASAP7_75t_L g204 ( .A(n_139), .B(n_109), .C(n_116), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_164), .B(n_124), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_156), .B(n_121), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_142), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_145), .B(n_118), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_151), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_133), .Y(n_215) );
INVxp67_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_156), .B(n_118), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_133), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_143), .A2(n_116), .B1(n_97), .B2(n_111), .Y(n_220) );
OR2x2_ASAP7_75t_SL g221 ( .A(n_152), .B(n_127), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_133), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_136), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_137), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_166), .B(n_123), .Y(n_226) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_173), .B(n_123), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_162), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_144), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_144), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_158), .B(n_119), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_158), .B(n_97), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_136), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_173), .B(n_119), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_171), .B(n_104), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_177), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_216), .B(n_149), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_233), .B(n_165), .Y(n_239) );
NOR3xp33_ASAP7_75t_SL g240 ( .A(n_185), .B(n_132), .C(n_150), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_208), .Y(n_241) );
NOR2xp33_ASAP7_75t_R g242 ( .A(n_177), .B(n_146), .Y(n_242) );
OR2x6_ASAP7_75t_L g243 ( .A(n_177), .B(n_166), .Y(n_243) );
NOR3xp33_ASAP7_75t_SL g244 ( .A(n_205), .B(n_154), .C(n_140), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_233), .B(n_171), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_226), .B(n_159), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_194), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_226), .B(n_170), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_233), .B(n_170), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_225), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_226), .B(n_167), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_176), .A2(n_165), .B(n_167), .C(n_166), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_235), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_182), .B(n_85), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_236), .B(n_144), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_200), .A2(n_160), .B1(n_108), .B2(n_91), .Y(n_259) );
BUFx10_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_227), .A2(n_104), .B1(n_111), .B2(n_95), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_200), .A2(n_107), .B(n_91), .C(n_95), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_226), .B(n_160), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_204), .B(n_138), .C(n_100), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_236), .B(n_147), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_174), .B(n_160), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_201), .B(n_157), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_235), .B(n_160), .Y(n_269) );
BUFx6f_ASAP7_75t_SL g270 ( .A(n_227), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_194), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_212), .B(n_96), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
BUFx4_ASAP7_75t_SL g275 ( .A(n_206), .Y(n_275) );
OR2x6_ASAP7_75t_L g276 ( .A(n_235), .B(n_107), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_230), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_220), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_179), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_176), .B(n_5), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_207), .B(n_160), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_232), .B(n_96), .C(n_100), .Y(n_282) );
NOR3xp33_ASAP7_75t_SL g283 ( .A(n_217), .B(n_101), .C(n_108), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_194), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_203), .A2(n_114), .B1(n_113), .B2(n_101), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_228), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_187), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_190), .Y(n_291) );
NOR3xp33_ASAP7_75t_SL g292 ( .A(n_217), .B(n_113), .C(n_7), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_180), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_207), .B(n_99), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_230), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_188), .A2(n_99), .B(n_136), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_187), .B(n_99), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_210), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_207), .B(n_89), .Y(n_300) );
INVx5_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_218), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_187), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_242), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_272), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_281), .A2(n_188), .B(n_203), .Y(n_307) );
OAI22xp5_ASAP7_75t_SL g308 ( .A1(n_278), .A2(n_221), .B1(n_202), .B2(n_174), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_274), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_269), .A2(n_197), .B(n_193), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g311 ( .A1(n_270), .A2(n_212), .B1(n_174), .B2(n_193), .Y(n_311) );
OAI21xp33_ASAP7_75t_SL g312 ( .A1(n_276), .A2(n_195), .B(n_181), .Y(n_312) );
BUFx2_ASAP7_75t_SL g313 ( .A(n_249), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_298), .A2(n_197), .B(n_193), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_250), .B(n_218), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_252), .B(n_221), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_250), .B(n_253), .Y(n_318) );
NOR2xp33_ASAP7_75t_SL g319 ( .A(n_287), .B(n_175), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_262), .A2(n_195), .B(n_197), .C(n_222), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_250), .B(n_186), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_279), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_253), .B(n_186), .Y(n_323) );
INVx8_ASAP7_75t_L g324 ( .A(n_253), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_279), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_248), .B(n_184), .Y(n_327) );
CKINVDCx11_ASAP7_75t_R g328 ( .A(n_276), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_276), .A2(n_222), .B1(n_231), .B2(n_219), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_237), .Y(n_330) );
AOI21x1_ASAP7_75t_L g331 ( .A1(n_298), .A2(n_181), .B(n_178), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_257), .A2(n_175), .B(n_184), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_275), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_249), .B(n_178), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_257), .A2(n_175), .B(n_231), .Y(n_337) );
INVx6_ASAP7_75t_L g338 ( .A(n_260), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_248), .B(n_191), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_271), .B(n_223), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_271), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_284), .B(n_191), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_258), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_276), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_284), .B(n_223), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_241), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_248), .B(n_199), .Y(n_348) );
BUFx4_ASAP7_75t_SL g349 ( .A(n_291), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_237), .Y(n_350) );
INVx5_ASAP7_75t_L g351 ( .A(n_272), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_256), .B(n_199), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_255), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_289), .A2(n_219), .B1(n_211), .B2(n_214), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_270), .A2(n_261), .B1(n_243), .B2(n_278), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_273), .B(n_213), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_265), .Y(n_358) );
CKINVDCx6p67_ASAP7_75t_R g359 ( .A(n_328), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_260), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_310), .A2(n_266), .B(n_288), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_308), .A2(n_243), .B1(n_260), .B2(n_263), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
CKINVDCx8_ASAP7_75t_R g364 ( .A(n_313), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_324), .B(n_280), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_307), .A2(n_290), .B(n_299), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_318), .A2(n_243), .B1(n_286), .B2(n_263), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_314), .A2(n_246), .B(n_251), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_324), .B(n_239), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_305), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_345), .A2(n_311), .B1(n_315), .B2(n_356), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_358), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_309), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_334), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_357), .B(n_263), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_357), .B(n_245), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_325), .Y(n_383) );
BUFx12f_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_321), .A2(n_323), .B1(n_341), .B2(n_346), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_335), .B(n_286), .Y(n_386) );
AOI32xp33_ASAP7_75t_L g387 ( .A1(n_312), .A2(n_291), .A3(n_268), .B1(n_259), .B2(n_267), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_341), .B(n_245), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_317), .B(n_238), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_335), .B(n_283), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_340), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_343), .A2(n_243), .B1(n_242), .B2(n_267), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_377), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_384), .A2(n_344), .B1(n_313), .B2(n_339), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_366), .A2(n_320), .B(n_316), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_384), .A2(n_348), .B1(n_343), .B2(n_327), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_385), .A2(n_346), .B1(n_341), .B2(n_329), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_361), .A2(n_331), .B(n_254), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_380), .B(n_309), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_369), .A2(n_262), .B(n_331), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_381), .B(n_346), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_376), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_389), .A2(n_240), .B1(n_282), .B2(n_244), .C(n_292), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_381), .B(n_346), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_373), .B(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
AND2x4_ASAP7_75t_SL g412 ( .A(n_368), .B(n_342), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_380), .B(n_316), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_367), .A2(n_305), .B1(n_294), .B2(n_350), .Y(n_414) );
INVx4_ASAP7_75t_L g415 ( .A(n_363), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_390), .A2(n_350), .B1(n_300), .B2(n_211), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_364), .A2(n_354), .B1(n_352), .B2(n_319), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_372), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_362), .A2(n_213), .B1(n_214), .B2(n_342), .Y(n_419) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_359), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_386), .A2(n_342), .B1(n_322), .B2(n_326), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_412), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_398), .A2(n_388), .B1(n_360), .B2(n_368), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_404), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_408), .A2(n_359), .B1(n_392), .B2(n_365), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_415), .B(n_379), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_398), .A2(n_364), .B1(n_363), .B2(n_371), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_414), .A2(n_388), .B1(n_387), .B2(n_370), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_404), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_420), .A2(n_360), .B1(n_374), .B2(n_391), .C1(n_383), .C2(n_371), .Y(n_432) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_395), .A2(n_297), .B(n_264), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_420), .A2(n_378), .B1(n_388), .B2(n_363), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_405), .A2(n_378), .B1(n_259), .B2(n_338), .C(n_330), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g436 ( .A1(n_417), .A2(n_363), .B(n_342), .C(n_267), .Y(n_436) );
OAI33xp33_ASAP7_75t_L g437 ( .A1(n_418), .A2(n_215), .A3(n_229), .B1(n_189), .B2(n_196), .B3(n_12), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_404), .Y(n_439) );
BUFx2_ASAP7_75t_SL g440 ( .A(n_402), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_415), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_393), .B(n_322), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_393), .B(n_326), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_414), .A2(n_363), .B1(n_338), .B2(n_330), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
OAI33xp33_ASAP7_75t_L g446 ( .A1(n_418), .A2(n_215), .A3(n_229), .B1(n_189), .B2(n_196), .B3(n_12), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_405), .B(n_89), .C(n_168), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_379), .Y(n_448) );
AOI322xp5_ASAP7_75t_L g449 ( .A1(n_408), .A2(n_6), .A3(n_8), .B1(n_9), .B2(n_11), .C1(n_13), .C2(n_14), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
NAND2x1_ASAP7_75t_L g451 ( .A(n_393), .B(n_379), .Y(n_451) );
OAI31xp33_ASAP7_75t_L g452 ( .A1(n_417), .A2(n_396), .A3(n_394), .B(n_402), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_338), .B1(n_272), .B2(n_301), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g454 ( .A1(n_394), .A2(n_301), .B(n_89), .C(n_351), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_397), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_397), .B(n_336), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_409), .B(n_336), .Y(n_457) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_455), .B(n_403), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_435), .A2(n_409), .B(n_411), .C(n_396), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_430), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_422), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_429), .B(n_397), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_429), .B(n_397), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_438), .B(n_406), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_425), .B(n_411), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_438), .B(n_406), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_434), .B(n_415), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_432), .B(n_406), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_450), .B(n_400), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_442), .B(n_400), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_439), .B(n_403), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_439), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_442), .B(n_400), .Y(n_476) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_449), .A2(n_423), .B(n_452), .C(n_436), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_427), .A2(n_407), .B1(n_403), .B2(n_413), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_422), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_443), .B(n_413), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_448), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_434), .B(n_403), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_448), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_451), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_456), .B(n_449), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_456), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g487 ( .A1(n_436), .A2(n_416), .B(n_419), .C(n_415), .Y(n_487) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_454), .A2(n_416), .B(n_419), .C(n_415), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_457), .B(n_413), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
OR2x6_ASAP7_75t_L g491 ( .A(n_440), .B(n_407), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_447), .A2(n_395), .B(n_399), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g493 ( .A(n_428), .B(n_421), .C(n_407), .D(n_403), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_445), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_445), .B(n_407), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_441), .B(n_426), .Y(n_497) );
OAI33xp33_ASAP7_75t_L g498 ( .A1(n_444), .A2(n_6), .A3(n_8), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_498) );
AOI33xp33_ASAP7_75t_L g499 ( .A1(n_453), .A2(n_421), .A3(n_407), .B1(n_403), .B2(n_412), .B3(n_21), .Y(n_499) );
NAND2x1_ASAP7_75t_L g500 ( .A(n_441), .B(n_407), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_440), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_441), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_426), .B(n_402), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_426), .B(n_402), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_471), .B(n_468), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_472), .B(n_16), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_459), .B(n_460), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_479), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_474), .B(n_431), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_477), .A2(n_89), .B(n_168), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_459), .B(n_401), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_464), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_476), .B(n_412), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_481), .B(n_401), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_476), .B(n_89), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_497), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_474), .B(n_17), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_499), .B(n_168), .C(n_401), .Y(n_523) );
OAI32xp33_ASAP7_75t_L g524 ( .A1(n_482), .A2(n_446), .A3(n_437), .B1(n_21), .B2(n_22), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_480), .B(n_18), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_461), .B(n_168), .C(n_401), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_480), .B(n_18), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_486), .B(n_19), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_465), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_481), .B(n_401), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_465), .Y(n_533) );
NAND2x2_ASAP7_75t_L g534 ( .A(n_485), .B(n_349), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_458), .B(n_19), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_465), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_467), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_489), .B(n_22), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_497), .Y(n_539) );
NOR4xp25_ASAP7_75t_SL g540 ( .A(n_502), .B(n_23), .C(n_433), .D(n_401), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_486), .B(n_399), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_467), .Y(n_542) );
OR2x6_ASAP7_75t_L g543 ( .A(n_491), .B(n_399), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_502), .B(n_168), .C(n_351), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_463), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_458), .B(n_433), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_463), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_483), .B(n_433), .Y(n_548) );
NOR4xp25_ASAP7_75t_SL g549 ( .A(n_498), .B(n_37), .C(n_40), .D(n_43), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_469), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_473), .B(n_333), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_462), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_493), .A2(n_333), .B1(n_338), .B2(n_306), .C(n_351), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_496), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_462), .B(n_168), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_462), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_458), .B(n_351), .Y(n_557) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_493), .A2(n_332), .B(n_337), .C(n_296), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_466), .B(n_351), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_491), .B(n_306), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_466), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_466), .B(n_306), .Y(n_562) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_553), .A2(n_470), .B(n_478), .C(n_487), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_519), .B(n_484), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_553), .A2(n_488), .B(n_500), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_534), .A2(n_523), .B1(n_529), .B2(n_535), .Y(n_567) );
AOI221x1_ASAP7_75t_L g568 ( .A1(n_512), .A2(n_492), .B1(n_490), .B2(n_484), .C(n_503), .Y(n_568) );
AOI211xp5_ASAP7_75t_SL g569 ( .A1(n_507), .A2(n_506), .B(n_505), .C(n_495), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_509), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_552), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_542), .B(n_503), .Y(n_572) );
NOR2xp33_ASAP7_75t_SL g573 ( .A(n_510), .B(n_494), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_520), .B(n_494), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_522), .A2(n_491), .B1(n_500), .B2(n_501), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_554), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_509), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
AOI211xp5_ASAP7_75t_L g579 ( .A1(n_525), .A2(n_490), .B(n_484), .C(n_504), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_537), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_527), .B(n_490), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_550), .B(n_504), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_538), .A2(n_503), .B(n_501), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_508), .A2(n_504), .B(n_501), .C(n_491), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_547), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_533), .B(n_491), .Y(n_586) );
AOI32xp33_ASAP7_75t_L g587 ( .A1(n_516), .A2(n_285), .A3(n_247), .B1(n_296), .B2(n_52), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_545), .B(n_44), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_521), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_539), .B(n_554), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_548), .B(n_46), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_524), .A2(n_247), .B(n_285), .C(n_58), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_530), .A2(n_301), .B1(n_272), .B2(n_183), .C(n_192), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_546), .A2(n_301), .B1(n_285), .B2(n_247), .Y(n_595) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_548), .A2(n_47), .B(n_54), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_536), .B(n_61), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_561), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_541), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_528), .B(n_514), .Y(n_600) );
AOI321xp33_ASAP7_75t_L g601 ( .A1(n_518), .A2(n_63), .A3(n_65), .B1(n_68), .B2(n_69), .C(n_70), .Y(n_601) );
XNOR2x1_ASAP7_75t_L g602 ( .A(n_551), .B(n_74), .Y(n_602) );
NOR2xp67_ASAP7_75t_L g603 ( .A(n_544), .B(n_78), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_511), .B(n_224), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_526), .A2(n_175), .B1(n_183), .B2(n_192), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_555), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_567), .A2(n_543), .B1(n_557), .B2(n_531), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_599), .B(n_532), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_589), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_602), .A2(n_559), .B(n_543), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_566), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_579), .B(n_560), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_600), .B(n_543), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_585), .B(n_560), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_571), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_570), .B(n_513), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_564), .B(n_559), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_578), .Y(n_619) );
NOR2x1_ASAP7_75t_L g620 ( .A(n_603), .B(n_562), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_577), .B(n_562), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_576), .A2(n_558), .B(n_549), .Y(n_622) );
NOR2xp33_ASAP7_75t_R g623 ( .A(n_573), .B(n_540), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_564), .B(n_224), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_580), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_584), .B(n_602), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_563), .A2(n_224), .B1(n_183), .B2(n_192), .C(n_198), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_590), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_581), .B(n_224), .Y(n_629) );
NOR4xp25_ASAP7_75t_SL g630 ( .A(n_576), .B(n_183), .C(n_192), .D(n_198), .Y(n_630) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_569), .B(n_175), .Y(n_631) );
NOR3xp33_ASAP7_75t_SL g632 ( .A(n_583), .B(n_183), .C(n_192), .Y(n_632) );
NOR4xp25_ASAP7_75t_SL g633 ( .A(n_594), .B(n_198), .C(n_234), .D(n_277), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_571), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_581), .B(n_234), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_592), .Y(n_636) );
XNOR2xp5_ASAP7_75t_L g637 ( .A(n_574), .B(n_234), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_598), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_565), .A2(n_593), .B(n_587), .Y(n_639) );
BUFx3_ASAP7_75t_L g640 ( .A(n_610), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_608), .B(n_606), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_626), .A2(n_575), .B1(n_595), .B2(n_572), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_611), .A2(n_595), .B1(n_586), .B2(n_582), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_638), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_613), .A2(n_588), .B(n_591), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_639), .B(n_601), .C(n_568), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_620), .B(n_597), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_636), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_619), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_632), .A2(n_597), .B(n_605), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_613), .A2(n_596), .B(n_605), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_637), .B(n_607), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_625), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_612), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_622), .A2(n_604), .B(n_234), .Y(n_655) );
AOI221xp5_ASAP7_75t_SL g656 ( .A1(n_628), .A2(n_277), .B1(n_295), .B2(n_614), .C(n_615), .Y(n_656) );
AOI221x1_ASAP7_75t_SL g657 ( .A1(n_642), .A2(n_621), .B1(n_609), .B2(n_617), .C(n_634), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_640), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_648), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_651), .A2(n_627), .B(n_633), .Y(n_660) );
AOI322xp5_ASAP7_75t_L g661 ( .A1(n_652), .A2(n_618), .A3(n_634), .B1(n_616), .B2(n_635), .C1(n_629), .C2(n_624), .Y(n_661) );
XOR2x2_ASAP7_75t_L g662 ( .A(n_643), .B(n_631), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_643), .A2(n_646), .B1(n_641), .B2(n_655), .C(n_653), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_649), .Y(n_664) );
BUFx3_ASAP7_75t_L g665 ( .A(n_654), .Y(n_665) );
NOR3x1_ASAP7_75t_L g666 ( .A(n_650), .B(n_623), .C(n_616), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_656), .B(n_624), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_656), .A2(n_647), .B1(n_645), .B2(n_650), .C(n_644), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_641), .B(n_629), .C(n_635), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_647), .A2(n_631), .B(n_630), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_642), .A2(n_295), .B1(n_643), .B2(n_646), .C(n_507), .Y(n_671) );
NAND2xp33_ASAP7_75t_L g672 ( .A(n_642), .B(n_626), .Y(n_672) );
NOR2x1p5_ASAP7_75t_L g673 ( .A(n_658), .B(n_666), .Y(n_673) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_665), .B(n_667), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_657), .B(n_671), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_663), .B(n_662), .Y(n_676) );
INVx1_ASAP7_75t_SL g677 ( .A(n_672), .Y(n_677) );
NOR4xp75_ASAP7_75t_L g678 ( .A(n_676), .B(n_668), .C(n_670), .D(n_663), .Y(n_678) );
NAND4xp25_ASAP7_75t_SL g679 ( .A(n_677), .B(n_661), .C(n_669), .D(n_660), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_675), .A2(n_660), .B(n_664), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_680), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_678), .Y(n_682) );
AOI22xp5_ASAP7_75t_SL g683 ( .A1(n_682), .A2(n_674), .B1(n_673), .B2(n_679), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_681), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_684), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_683), .B(n_659), .Y(n_686) );
endmodule