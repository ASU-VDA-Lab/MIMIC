module fake_netlist_5_1580_n_1919 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1919);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1919;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_27),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_41),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_94),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_97),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_61),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_36),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_167),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_156),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_11),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_56),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_40),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_109),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_110),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_75),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_28),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_76),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_126),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_150),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_103),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_64),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_114),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_170),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_106),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_107),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_31),
.Y(n_245)
);

BUFx2_ASAP7_75t_SL g246 ( 
.A(n_137),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_157),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_111),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_29),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_185),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_79),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_26),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_23),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_83),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_118),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_89),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_129),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_28),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_30),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_59),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_23),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_196),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_191),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_119),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_1),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_112),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_138),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_95),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_175),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_168),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_142),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_5),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_148),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_20),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_65),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_158),
.Y(n_288)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_87),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_35),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_26),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_193),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_64),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_66),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_70),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_202),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_85),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_127),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_37),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_182),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_117),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_84),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_57),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_183),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_57),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_12),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_159),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_42),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_179),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_30),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_169),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_58),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_125),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_147),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_176),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_45),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_115),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_203),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_8),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_67),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_52),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_173),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_120),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_199),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_32),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_42),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_17),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_78),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_74),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_86),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_163),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_8),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_33),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_116),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_63),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_194),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_101),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_7),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_51),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_139),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_92),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_4),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_53),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_4),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_178),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_67),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_132),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_162),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_48),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_165),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_6),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_38),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_47),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_100),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_65),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_50),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_104),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_186),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_62),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_16),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_15),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_54),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_121),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_146),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_39),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_38),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_108),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_124),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_51),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_54),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_19),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_90),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_72),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_31),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_166),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_9),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_59),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_35),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_102),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_73),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_49),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_47),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_1),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_82),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_140),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_192),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_60),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_15),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_18),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_188),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_60),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_180),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_40),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_77),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_43),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_130),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_21),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_155),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_181),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_22),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_274),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_249),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_220),
.B(n_0),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_334),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

BUFx6f_ASAP7_75t_SL g413 ( 
.A(n_231),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_377),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_274),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_0),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_244),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_274),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_274),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_231),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_274),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_324),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_216),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_254),
.B(n_3),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_252),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_330),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_254),
.B(n_3),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_321),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_205),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_258),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_328),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_265),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_265),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_287),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_249),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_207),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_261),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_210),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_213),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_217),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_298),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_374),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_268),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_206),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_269),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_228),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_402),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_208),
.Y(n_452)
);

BUFx2_ASAP7_75t_SL g453 ( 
.A(n_263),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_278),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_226),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_245),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_291),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_335),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_214),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_263),
.B(n_7),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_214),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_303),
.B(n_9),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_257),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_R g464 ( 
.A(n_250),
.B(n_128),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_221),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_230),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_292),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_287),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_220),
.B(n_10),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_251),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_303),
.B(n_10),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_255),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_270),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_260),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_306),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_311),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_214),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_319),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_325),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_279),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_262),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_206),
.B(n_11),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_283),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_286),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_331),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_332),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_294),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_295),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_249),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_214),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_241),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_267),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_247),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_212),
.B(n_14),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_216),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_344),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_223),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_253),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_273),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_315),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_223),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_236),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_372),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_236),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_300),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_301),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_337),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_315),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_315),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_338),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_212),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_339),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_227),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_445),
.B(n_227),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_453),
.B(n_266),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_470),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_472),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_424),
.A2(n_313),
.B1(n_320),
.B2(n_248),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_453),
.B(n_266),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_416),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_423),
.B(n_375),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_420),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_407),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_421),
.B(n_375),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_475),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_482),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_418),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_493),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_R g535 ( 
.A(n_428),
.B(n_209),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_452),
.B(n_302),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_496),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_500),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_431),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_425),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_458),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_435),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_429),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_465),
.B(n_466),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_446),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_492),
.B(n_302),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_433),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_451),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_448),
.Y(n_556)
);

NAND2x1_ASAP7_75t_L g557 ( 
.A(n_514),
.B(n_390),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_390),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_423),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_434),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_455),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_512),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_490),
.A2(n_243),
.B1(n_380),
.B2(n_371),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_421),
.B(n_391),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_512),
.Y(n_567)
);

CKINVDCx6p67_ASAP7_75t_R g568 ( 
.A(n_501),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_512),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_512),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_471),
.A2(n_391),
.B(n_259),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_440),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_436),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_514),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_436),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_433),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_441),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_441),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_447),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_411),
.B(n_256),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_432),
.B(n_271),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_447),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_459),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_449),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_449),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_461),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_461),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_478),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_412),
.B(n_272),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_510),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_454),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_432),
.B(n_276),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_478),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_454),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_R g597 ( 
.A(n_457),
.B(n_209),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_414),
.B(n_285),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_457),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_536),
.B(n_427),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_537),
.B(n_409),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_533),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_583),
.Y(n_603)
);

CKINVDCx16_ASAP7_75t_R g604 ( 
.A(n_531),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_536),
.B(n_430),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_536),
.B(n_460),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_517),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_533),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_536),
.B(n_467),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_548),
.B(n_424),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_526),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_551),
.B(n_462),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_572),
.Y(n_615)
);

AND2x2_ASAP7_75t_SL g616 ( 
.A(n_551),
.B(n_417),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_551),
.B(n_499),
.Y(n_617)
);

AND2x2_ASAP7_75t_SL g618 ( 
.A(n_551),
.B(n_495),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_515),
.B(n_467),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_543),
.B(n_476),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_516),
.B(n_476),
.Y(n_621)
);

INVx4_ASAP7_75t_SL g622 ( 
.A(n_533),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_442),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_575),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_583),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_528),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_575),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_533),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_520),
.B(n_498),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_517),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_558),
.B(n_498),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_533),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_582),
.A2(n_479),
.B1(n_480),
.B2(n_477),
.Y(n_635)
);

AND3x1_ASAP7_75t_L g636 ( 
.A(n_554),
.B(n_503),
.C(n_502),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_550),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_575),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_528),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_594),
.B(n_443),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_547),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_550),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_550),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g644 ( 
.A(n_519),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_594),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_592),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_577),
.B(n_439),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_552),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_561),
.B(n_477),
.Y(n_649)
);

BUFx10_ASAP7_75t_L g650 ( 
.A(n_559),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_594),
.B(n_290),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_594),
.B(n_479),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_557),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_561),
.B(n_480),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_559),
.A2(n_487),
.B1(n_508),
.B2(n_486),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_578),
.B(n_486),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_575),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_566),
.B(n_505),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_569),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_575),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_560),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_578),
.B(n_487),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_522),
.B(n_508),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_557),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_571),
.A2(n_483),
.B1(n_376),
.B2(n_394),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_539),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_569),
.B(n_563),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_521),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_569),
.B(n_511),
.Y(n_671)
);

BUFx4f_ASAP7_75t_L g672 ( 
.A(n_568),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_580),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_571),
.A2(n_376),
.B1(n_394),
.B2(n_372),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_524),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_550),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_591),
.B(n_509),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_580),
.B(n_513),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_598),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_565),
.B(n_513),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_574),
.B(n_444),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_581),
.B(n_408),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_581),
.B(n_305),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_525),
.B(n_413),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_584),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_564),
.B(n_567),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_556),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_585),
.B(n_225),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_556),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_574),
.A2(n_469),
.B1(n_410),
.B2(n_309),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_584),
.B(n_317),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_586),
.B(n_342),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_525),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_585),
.B(n_595),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_535),
.A2(n_413),
.B1(n_354),
.B2(n_242),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_595),
.B(n_541),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_556),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_556),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_542),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_544),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_576),
.A2(n_382),
.B1(n_308),
.B2(n_326),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_576),
.A2(n_367),
.B1(n_358),
.B2(n_362),
.Y(n_704)
);

CKINVDCx6p67_ASAP7_75t_R g705 ( 
.A(n_568),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_541),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_587),
.B(n_415),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_556),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_518),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_553),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_573),
.B(n_450),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_593),
.B(n_596),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_570),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_553),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_573),
.B(n_456),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_544),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_595),
.B(n_312),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_546),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_546),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_599),
.B(n_224),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_579),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_542),
.B(n_264),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_570),
.B(n_343),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_588),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_588),
.B(n_369),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_570),
.B(n_347),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_518),
.B(n_463),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_527),
.Y(n_728)
);

BUFx4f_ASAP7_75t_L g729 ( 
.A(n_570),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_589),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_589),
.Y(n_731)
);

NOR2x1p5_ASAP7_75t_L g732 ( 
.A(n_527),
.B(n_238),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_590),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_590),
.B(n_474),
.Y(n_734)
);

OAI221xp5_ASAP7_75t_L g735 ( 
.A1(n_597),
.A2(n_507),
.B1(n_506),
.B2(n_481),
.C(n_484),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_530),
.B(n_485),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_530),
.B(n_214),
.Y(n_737)
);

INVx3_ASAP7_75t_R g738 ( 
.A(n_562),
.Y(n_738)
);

INVx5_ASAP7_75t_L g739 ( 
.A(n_540),
.Y(n_739)
);

INVx4_ASAP7_75t_SL g740 ( 
.A(n_545),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_545),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_681),
.A2(n_348),
.B1(n_364),
.B2(n_360),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_681),
.B(n_351),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_615),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_618),
.B(n_491),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_618),
.B(n_491),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_611),
.B(n_610),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_600),
.B(n_605),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_703),
.A2(n_341),
.B1(n_388),
.B2(n_383),
.C(n_366),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_683),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_720),
.B(n_549),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_683),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_606),
.B(n_214),
.Y(n_753)
);

BUFx5_ASAP7_75t_L g754 ( 
.A(n_651),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_616),
.A2(n_610),
.B1(n_619),
.B2(n_621),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_603),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_619),
.B(n_534),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_603),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_621),
.B(n_534),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_614),
.B(n_214),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_651),
.B(n_214),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_684),
.B(n_538),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_611),
.B(n_538),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_616),
.A2(n_246),
.B1(n_289),
.B2(n_370),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_666),
.A2(n_400),
.B1(n_381),
.B2(n_392),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_652),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_736),
.B(n_549),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_SL g768 ( 
.A1(n_644),
.A2(n_555),
.B1(n_368),
.B2(n_403),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_736),
.B(n_555),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_645),
.A2(n_356),
.B(n_373),
.C(n_396),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_645),
.B(n_275),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_655),
.B(n_489),
.C(n_488),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_631),
.B(n_238),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_613),
.B(n_437),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_666),
.A2(n_296),
.B1(n_401),
.B2(n_387),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_727),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_683),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_613),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_612),
.B(n_211),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_625),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_617),
.B(n_277),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_695),
.B(n_280),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_706),
.B(n_281),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_406),
.C(n_345),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_675),
.B(n_730),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_707),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_735),
.A2(n_243),
.B1(n_304),
.B2(n_349),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_675),
.B(n_296),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_741),
.B(n_437),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_609),
.A2(n_468),
.B(n_438),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_629),
.A2(n_304),
.B1(n_349),
.B2(n_350),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_722),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_739),
.B(n_282),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_609),
.B(n_215),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_721),
.B(n_296),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_714),
.B(n_284),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_659),
.B(n_215),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_731),
.Y(n_798)
);

INVx6_ASAP7_75t_L g799 ( 
.A(n_739),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_625),
.B(n_438),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_739),
.Y(n_801)
);

INVx8_ASAP7_75t_L g802 ( 
.A(n_739),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_697),
.B(n_218),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_679),
.B(n_601),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_692),
.A2(n_361),
.B1(n_350),
.B2(n_352),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_660),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_678),
.B(n_288),
.Y(n_807)
);

BUFx5_ASAP7_75t_L g808 ( 
.A(n_651),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_678),
.B(n_293),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_682),
.B(n_219),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_731),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_219),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_634),
.B(n_297),
.Y(n_813)
);

BUFx5_ASAP7_75t_L g814 ( 
.A(n_651),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_641),
.B(n_299),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_653),
.A2(n_307),
.B(n_310),
.C(n_314),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_731),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_711),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_648),
.B(n_316),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_685),
.B(n_222),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_662),
.B(n_318),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_620),
.B(n_468),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_653),
.A2(n_296),
.B1(n_359),
.B2(n_352),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_731),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_649),
.Y(n_825)
);

INVxp33_ASAP7_75t_L g826 ( 
.A(n_656),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_692),
.A2(n_361),
.B1(n_355),
.B2(n_359),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_690),
.B(n_322),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_663),
.B(n_473),
.Y(n_829)
);

AND2x2_ASAP7_75t_SL g830 ( 
.A(n_604),
.B(n_473),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_646),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_737),
.B(n_363),
.C(n_232),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_711),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_626),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_717),
.B(n_323),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_725),
.B(n_229),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_724),
.B(n_296),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_660),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_715),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_651),
.B(n_296),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_665),
.B(n_327),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_680),
.B(n_497),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_665),
.B(n_329),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_623),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_685),
.B(n_233),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_623),
.A2(n_333),
.B(n_346),
.C(n_340),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_670),
.B(n_336),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_679),
.B(n_497),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_654),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_SL g851 ( 
.A1(n_674),
.A2(n_371),
.B1(n_355),
.B2(n_365),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_733),
.B(n_296),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_679),
.B(n_601),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_698),
.B(n_296),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_664),
.B(n_233),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_639),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_623),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_640),
.A2(n_384),
.B1(n_393),
.B2(n_368),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_693),
.B(n_234),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_693),
.A2(n_504),
.B(n_464),
.C(n_405),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_694),
.B(n_234),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_640),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_694),
.B(n_235),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_716),
.B(n_235),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_718),
.B(n_237),
.Y(n_865)
);

AOI22x1_ASAP7_75t_L g866 ( 
.A1(n_673),
.A2(n_385),
.B1(n_405),
.B2(n_404),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_676),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_640),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_719),
.B(n_237),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_710),
.A2(n_385),
.B(n_404),
.C(n_240),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_671),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_871)
);

NOR2x1p5_ASAP7_75t_L g872 ( 
.A(n_705),
.B(n_380),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_658),
.B(n_239),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_674),
.B(n_504),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_710),
.A2(n_387),
.B1(n_399),
.B2(n_384),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_658),
.B(n_353),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_667),
.B(n_353),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_732),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_701),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_667),
.B(n_354),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_647),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_669),
.A2(n_395),
.B1(n_399),
.B2(n_393),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_674),
.B(n_395),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_686),
.B(n_398),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_669),
.B(n_398),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_702),
.B(n_386),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_624),
.B(n_386),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_688),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_636),
.B(n_379),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_624),
.B(n_379),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_748),
.A2(n_729),
.B(n_608),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_757),
.B(n_712),
.C(n_630),
.Y(n_892)
);

BUFx4f_ASAP7_75t_L g893 ( 
.A(n_802),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_748),
.A2(n_729),
.B(n_668),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_857),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_785),
.A2(n_632),
.B(n_643),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_755),
.A2(n_644),
.B1(n_723),
.B2(n_726),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_745),
.A2(n_696),
.B(n_726),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_747),
.B(n_687),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_774),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_785),
.A2(n_723),
.B(n_702),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_745),
.A2(n_734),
.B(n_627),
.Y(n_902)
);

OR2x2_ASAP7_75t_SL g903 ( 
.A(n_751),
.B(n_738),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_746),
.A2(n_643),
.B(n_637),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_774),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_888),
.B(n_734),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_746),
.A2(n_628),
.B(n_632),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_756),
.Y(n_908)
);

OAI321xp33_ASAP7_75t_L g909 ( 
.A1(n_810),
.A2(n_703),
.A3(n_704),
.B1(n_397),
.B2(n_403),
.C(n_22),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_753),
.A2(n_628),
.B(n_632),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_776),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_759),
.B(n_607),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_763),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_825),
.B(n_638),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_850),
.B(n_638),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_857),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_812),
.A2(n_672),
.B(n_704),
.C(n_661),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_760),
.A2(n_628),
.B(n_637),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_857),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_800),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_766),
.A2(n_661),
.B1(n_657),
.B2(n_709),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_822),
.B(n_687),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_802),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_760),
.A2(n_643),
.B(n_637),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_842),
.A2(n_602),
.B(n_642),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_743),
.A2(n_699),
.B(n_689),
.C(n_691),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_829),
.B(n_699),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_862),
.B(n_687),
.Y(n_928)
);

AND2x2_ASAP7_75t_SL g929 ( 
.A(n_767),
.B(n_728),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_843),
.B(n_689),
.Y(n_930)
);

OAI321xp33_ASAP7_75t_L g931 ( 
.A1(n_787),
.A2(n_397),
.A3(n_16),
.B1(n_17),
.B2(n_20),
.C(n_24),
.Y(n_931)
);

CKINVDCx10_ASAP7_75t_R g932 ( 
.A(n_831),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_844),
.A2(n_602),
.B(n_642),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_788),
.A2(n_713),
.B(n_708),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_802),
.B(n_705),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_L g936 ( 
.A(n_820),
.B(n_701),
.C(n_650),
.Y(n_936)
);

NOR2x1_ASAP7_75t_L g937 ( 
.A(n_801),
.B(n_677),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_765),
.B(n_642),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_788),
.A2(n_700),
.B(n_633),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_781),
.A2(n_602),
.B(n_677),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_800),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_797),
.B(n_677),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_771),
.A2(n_642),
.B(n_700),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_854),
.A2(n_811),
.B(n_798),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_794),
.B(n_622),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_807),
.A2(n_700),
.B(n_633),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_846),
.B(n_622),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_859),
.B(n_622),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_818),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_809),
.A2(n_633),
.B(n_700),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_833),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_769),
.B(n_650),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_861),
.B(n_740),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_863),
.B(n_740),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_831),
.B(n_728),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_789),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_862),
.B(n_728),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_790),
.A2(n_177),
.B(n_174),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_828),
.B(n_14),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_817),
.A2(n_824),
.B(n_835),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_764),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_831),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_834),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_837),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_890),
.A2(n_80),
.B(n_164),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_887),
.A2(n_161),
.B(n_154),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_SL g967 ( 
.A1(n_816),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_967)
);

AO22x1_ASAP7_75t_L g968 ( 
.A1(n_826),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_782),
.A2(n_81),
.B(n_151),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_758),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_750),
.B(n_752),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_806),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_777),
.A2(n_34),
.B(n_41),
.C(n_43),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_784),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_783),
.A2(n_88),
.B(n_145),
.Y(n_975)
);

AO32x1_ASAP7_75t_L g976 ( 
.A1(n_840),
.A2(n_44),
.A3(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_790),
.B(n_874),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_796),
.A2(n_93),
.B(n_144),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_789),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_870),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_744),
.B(n_867),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_868),
.A2(n_99),
.B1(n_141),
.B2(n_136),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_792),
.B(n_55),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_860),
.A2(n_58),
.B(n_62),
.C(n_63),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_R g985 ( 
.A(n_879),
.B(n_105),
.Y(n_985)
);

OAI21xp33_ASAP7_75t_L g986 ( 
.A1(n_875),
.A2(n_66),
.B(n_68),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_845),
.B(n_113),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_799),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_780),
.B(n_91),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_742),
.A2(n_69),
.B(n_96),
.C(n_123),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_786),
.B(n_133),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_761),
.A2(n_134),
.B(n_152),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_856),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_778),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_778),
.B(n_873),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_778),
.B(n_873),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_841),
.A2(n_813),
.B(n_821),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_775),
.A2(n_823),
.B1(n_858),
.B2(n_851),
.Y(n_998)
);

NOR2x1p5_ASAP7_75t_L g999 ( 
.A(n_804),
.B(n_853),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_815),
.A2(n_819),
.B(n_848),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_795),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_832),
.A2(n_847),
.B(n_886),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_883),
.B(n_830),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_849),
.B(n_876),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_878),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_877),
.B(n_880),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_871),
.A2(n_880),
.B(n_886),
.C(n_885),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_789),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_885),
.A2(n_865),
.B(n_864),
.C(n_869),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_773),
.B(n_762),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_806),
.B(n_839),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_795),
.A2(n_852),
.B(n_838),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_838),
.A2(n_852),
.B(n_865),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_793),
.B(n_872),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_864),
.A2(n_869),
.B(n_836),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_855),
.B(n_768),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_779),
.B(n_799),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_803),
.A2(n_884),
.B(n_770),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_799),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_754),
.A2(n_814),
.B(n_808),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_772),
.B(n_814),
.Y(n_1021)
);

AOI33xp33_ASAP7_75t_L g1022 ( 
.A1(n_791),
.A2(n_882),
.A3(n_827),
.B1(n_805),
.B2(n_749),
.B3(n_881),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_866),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_754),
.A2(n_808),
.B(n_814),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_754),
.A2(n_808),
.B(n_814),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_808),
.A2(n_814),
.B(n_889),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_814),
.B(n_805),
.Y(n_1027)
);

AO22x1_ASAP7_75t_L g1028 ( 
.A1(n_827),
.A2(n_644),
.B1(n_757),
.B2(n_810),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_748),
.B(n_755),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_748),
.B(n_755),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_755),
.A2(n_748),
.B1(n_618),
.B2(n_747),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_755),
.A2(n_765),
.B1(n_748),
.B2(n_764),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_845),
.B(n_868),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_748),
.A2(n_785),
.B(n_746),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_879),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_748),
.A2(n_737),
.B(n_812),
.C(n_810),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_755),
.B(n_747),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_748),
.B(n_755),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_747),
.B(n_610),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_748),
.A2(n_785),
.B(n_746),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_774),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_748),
.A2(n_785),
.B(n_746),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_755),
.B(n_757),
.Y(n_1043)
);

OAI321xp33_ASAP7_75t_L g1044 ( 
.A1(n_755),
.A2(n_810),
.A3(n_812),
.B1(n_787),
.B2(n_742),
.C(n_749),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_748),
.A2(n_737),
.B(n_812),
.C(n_810),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_747),
.B(n_610),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_755),
.A2(n_812),
.B(n_810),
.C(n_748),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_748),
.B(n_755),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_748),
.A2(n_785),
.B(n_746),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_774),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_748),
.A2(n_785),
.B(n_746),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_1036),
.C(n_1047),
.Y(n_1052)
);

AO21x2_ASAP7_75t_L g1053 ( 
.A1(n_939),
.A2(n_934),
.B(n_1002),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1020),
.A2(n_1025),
.B(n_1024),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_949),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_912),
.B(n_952),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_1021),
.A2(n_945),
.B(n_947),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_SL g1059 ( 
.A1(n_1029),
.A2(n_1048),
.B(n_1030),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_910),
.A2(n_924),
.B(n_918),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_997),
.A2(n_1051),
.B(n_1040),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1016),
.A2(n_1032),
.B1(n_1031),
.B2(n_1039),
.Y(n_1062)
);

AO31x2_ASAP7_75t_L g1063 ( 
.A1(n_1009),
.A2(n_1032),
.A3(n_1007),
.B(n_1042),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_934),
.A2(n_939),
.B(n_1034),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1033),
.B(n_987),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1006),
.B(n_1046),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_951),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_940),
.A2(n_933),
.B(n_925),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1006),
.B(n_1049),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_1013),
.A2(n_1012),
.A3(n_984),
.B(n_894),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_897),
.A2(n_906),
.B1(n_1037),
.B2(n_977),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_904),
.A2(n_907),
.B(n_1026),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1004),
.B(n_1001),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1004),
.B(n_995),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_913),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_936),
.B(n_911),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_996),
.B(n_1000),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_998),
.A2(n_1027),
.B1(n_961),
.B2(n_958),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1010),
.B(n_922),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_899),
.B(n_1028),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1003),
.B(n_892),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_891),
.A2(n_927),
.B(n_930),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_L g1083 ( 
.A1(n_1018),
.A2(n_1002),
.B(n_948),
.C(n_959),
.Y(n_1083)
);

INVx3_ASAP7_75t_SL g1084 ( 
.A(n_1035),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_981),
.B(n_964),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_900),
.B(n_920),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_895),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1019),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_898),
.A2(n_901),
.B(n_943),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_971),
.B(n_905),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_941),
.B(n_1050),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1041),
.B(n_914),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_902),
.A2(n_1044),
.B(n_998),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1022),
.A2(n_986),
.B(n_958),
.C(n_917),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_915),
.B(n_942),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_895),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_946),
.A2(n_950),
.B(n_926),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_961),
.A2(n_929),
.B1(n_987),
.B2(n_938),
.Y(n_1098)
);

AOI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_909),
.A2(n_1023),
.B(n_980),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_908),
.B(n_1017),
.Y(n_1100)
);

OAI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_983),
.A2(n_1008),
.B1(n_956),
.B2(n_979),
.C(n_1014),
.Y(n_1101)
);

AOI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_931),
.A2(n_954),
.B(n_953),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_965),
.A2(n_966),
.B(n_963),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_973),
.A2(n_969),
.A3(n_978),
.B(n_975),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1011),
.B(n_991),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1033),
.B(n_999),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_970),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_937),
.A2(n_1011),
.B(n_992),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_962),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_895),
.B(n_916),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_993),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_903),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_916),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_990),
.A2(n_931),
.B(n_928),
.C(n_921),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_919),
.B(n_972),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_970),
.A2(n_919),
.B(n_994),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_970),
.A2(n_919),
.B(n_994),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_970),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_972),
.B(n_968),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_957),
.A2(n_893),
.B(n_923),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_893),
.A2(n_923),
.B(n_972),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_982),
.A2(n_989),
.B(n_967),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1019),
.B(n_974),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1019),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_989),
.A2(n_988),
.B(n_976),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_985),
.B(n_955),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_932),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_976),
.A2(n_955),
.B(n_935),
.C(n_1005),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_935),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1020),
.A2(n_1025),
.B(n_1024),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1047),
.A2(n_1009),
.A3(n_1032),
.B(n_1007),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1034),
.A2(n_1051),
.B(n_1049),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_912),
.B(n_1043),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_949),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1043),
.A2(n_755),
.B1(n_1047),
.B2(n_1030),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_913),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_L g1142 ( 
.A(n_1047),
.B(n_1029),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1034),
.A2(n_1051),
.B(n_1049),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1043),
.A2(n_755),
.B(n_1032),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1043),
.A2(n_755),
.B(n_610),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1043),
.A2(n_755),
.B1(n_1047),
.B2(n_1030),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1033),
.B(n_845),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1043),
.A2(n_755),
.B1(n_1016),
.B2(n_1029),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_895),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_895),
.Y(n_1154)
);

CKINVDCx8_ASAP7_75t_R g1155 ( 
.A(n_932),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_949),
.Y(n_1158)
);

AOI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1015),
.A2(n_1040),
.B(n_1034),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1033),
.B(n_845),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_845),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_1043),
.A2(n_1047),
.B(n_1028),
.C(n_1018),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_1035),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_913),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1047),
.A2(n_1009),
.A3(n_1032),
.B(n_1007),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_944),
.A2(n_896),
.B(n_960),
.Y(n_1171)
);

AOI221x1_ASAP7_75t_L g1172 ( 
.A1(n_1043),
.A2(n_1047),
.B1(n_1032),
.B2(n_1030),
.C(n_1038),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1028),
.A2(n_909),
.B1(n_791),
.B2(n_1043),
.C(n_827),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1047),
.A2(n_1043),
.B(n_1044),
.C(n_1037),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1034),
.A2(n_1051),
.B(n_1049),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1043),
.A2(n_755),
.B1(n_1016),
.B2(n_1029),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1016),
.A2(n_755),
.B1(n_1043),
.B2(n_757),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1034),
.A2(n_1051),
.B(n_1049),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_949),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1028),
.A2(n_909),
.B1(n_791),
.B2(n_1043),
.C(n_827),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1079),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1067),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1075),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1077),
.A2(n_1131),
.B(n_1054),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1143),
.B(n_1160),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1148),
.A2(n_1151),
.B1(n_1176),
.B2(n_1182),
.C(n_1173),
.Y(n_1189)
);

AND2x2_ASAP7_75t_SL g1190 ( 
.A(n_1062),
.B(n_1142),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_1087),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1158),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1167),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1141),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1093),
.A2(n_1078),
.B(n_1165),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1088),
.Y(n_1196)
);

AND2x6_ASAP7_75t_L g1197 ( 
.A(n_1130),
.B(n_1137),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1066),
.B(n_1130),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1066),
.B(n_1137),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1081),
.B(n_1157),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1084),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1112),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1168),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1129),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1088),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1087),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1162),
.B(n_1179),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1155),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1065),
.B(n_1106),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1088),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1156),
.B(n_1181),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1069),
.A2(n_1061),
.B(n_1059),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1177),
.B(n_1065),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1150),
.B(n_1163),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1156),
.B(n_1074),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1074),
.B(n_1073),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1139),
.A2(n_1149),
.B1(n_1146),
.B2(n_1078),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1107),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1135),
.A2(n_1175),
.B(n_1145),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_1107),
.Y(n_1222)
);

INVx8_ASAP7_75t_L g1223 ( 
.A(n_1087),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_SL g1224 ( 
.A(n_1164),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1164),
.B(n_1124),
.Y(n_1225)
);

NAND2x1_ASAP7_75t_L g1226 ( 
.A(n_1096),
.B(n_1153),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1138),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1109),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1124),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1073),
.B(n_1085),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1172),
.B(n_1071),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1080),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1090),
.B(n_1091),
.Y(n_1233)
);

OR2x6_ASAP7_75t_SL g1234 ( 
.A(n_1126),
.B(n_1123),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1083),
.A2(n_1178),
.B(n_1089),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1115),
.Y(n_1236)
);

CKINVDCx8_ASAP7_75t_R g1237 ( 
.A(n_1127),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1123),
.Y(n_1238)
);

OR2x2_ASAP7_75t_SL g1239 ( 
.A(n_1126),
.B(n_1119),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1146),
.B(n_1174),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_SL g1241 ( 
.A1(n_1052),
.A2(n_1094),
.B(n_1093),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1105),
.B(n_1095),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1092),
.B(n_1180),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1153),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1115),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1100),
.B(n_1086),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1111),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1098),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1154),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_SL g1250 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1098),
.C(n_1122),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1154),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1121),
.B(n_1120),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1133),
.B(n_1170),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1122),
.A2(n_1102),
.B(n_1101),
.C(n_1125),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1119),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1133),
.B(n_1170),
.Y(n_1256)
);

NAND2x1p5_ASAP7_75t_L g1257 ( 
.A(n_1110),
.B(n_1113),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1099),
.A2(n_1114),
.B(n_1076),
.C(n_1082),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1118),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1063),
.B(n_1053),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1053),
.A2(n_1064),
.B1(n_1128),
.B2(n_1103),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1063),
.B(n_1070),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1108),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1058),
.Y(n_1264)
);

OR2x6_ASAP7_75t_L g1265 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1070),
.B(n_1104),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1104),
.B(n_1070),
.C(n_1159),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1104),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1072),
.B(n_1097),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1060),
.A2(n_1057),
.B(n_1171),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_L g1271 ( 
.A(n_1132),
.B(n_1152),
.C(n_1134),
.Y(n_1271)
);

OAI221xp5_ASAP7_75t_L g1272 ( 
.A1(n_1144),
.A2(n_1161),
.B1(n_1166),
.B2(n_1169),
.C(n_1068),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_L g1274 ( 
.A(n_1088),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1136),
.A2(n_1148),
.B1(n_1043),
.B2(n_1173),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1079),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1075),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1075),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1157),
.B(n_1162),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1093),
.A2(n_1078),
.B(n_1165),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_1162),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1136),
.A2(n_1043),
.B1(n_1148),
.B2(n_1056),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1084),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1055),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1136),
.A2(n_1043),
.B1(n_1148),
.B2(n_1056),
.Y(n_1288)
);

AOI21xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1136),
.A2(n_1056),
.B(n_1028),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1088),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1136),
.A2(n_755),
.B1(n_1056),
.B2(n_1043),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1107),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1167),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1077),
.A2(n_1131),
.B(n_1054),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1075),
.Y(n_1296)
);

OR2x6_ASAP7_75t_L g1297 ( 
.A(n_1121),
.B(n_802),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1087),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1143),
.B(n_1160),
.Y(n_1299)
);

OAI321xp33_ASAP7_75t_L g1300 ( 
.A1(n_1136),
.A2(n_1148),
.A3(n_1182),
.B1(n_1173),
.B2(n_1056),
.C(n_755),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1136),
.A2(n_1056),
.B(n_1043),
.C(n_1148),
.Y(n_1301)
);

AND2x2_ASAP7_75t_SL g1302 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1067),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1065),
.B(n_1106),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1093),
.A2(n_1078),
.B(n_1165),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1136),
.B(n_1056),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1077),
.A2(n_1131),
.B(n_1054),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1075),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1143),
.B(n_1160),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1270),
.A2(n_1214),
.B(n_1271),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1223),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1236),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1292),
.A2(n_1282),
.B1(n_1310),
.B2(n_1284),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1192),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1285),
.A2(n_1288),
.B1(n_1309),
.B2(n_1273),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1302),
.A2(n_1278),
.B1(n_1189),
.B2(n_1290),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1187),
.A2(n_1307),
.B1(n_1306),
.B2(n_1190),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1215),
.B(n_1252),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1304),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1208),
.B(n_1285),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1245),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1288),
.A2(n_1275),
.B1(n_1230),
.B2(n_1303),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1251),
.Y(n_1327)
);

BUFx10_ASAP7_75t_L g1328 ( 
.A(n_1224),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1196),
.Y(n_1329)
);

INVx11_ASAP7_75t_L g1330 ( 
.A(n_1274),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1301),
.A2(n_1218),
.B1(n_1289),
.B2(n_1219),
.Y(n_1331)
);

OAI21xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1219),
.A2(n_1217),
.B(n_1204),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1268),
.Y(n_1333)
);

BUFx4_ASAP7_75t_SL g1334 ( 
.A(n_1209),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1186),
.A2(n_1295),
.B(n_1311),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1289),
.A2(n_1248),
.B1(n_1239),
.B2(n_1183),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1213),
.B(n_1280),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1253),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1216),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1223),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1252),
.B(n_1225),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1300),
.B(n_1200),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1227),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1287),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1207),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1240),
.A2(n_1308),
.B1(n_1195),
.B2(n_1281),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1183),
.A2(n_1276),
.B1(n_1238),
.B2(n_1283),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1291),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1223),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1247),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1256),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1224),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1201),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1243),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1195),
.A2(n_1281),
.B1(n_1308),
.B2(n_1232),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1185),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1237),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1232),
.A2(n_1199),
.B1(n_1198),
.B2(n_1231),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1276),
.A2(n_1233),
.B1(n_1212),
.B2(n_1234),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1259),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1242),
.A2(n_1255),
.B1(n_1300),
.B2(n_1197),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1246),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1271),
.A2(n_1221),
.B(n_1272),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1207),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1266),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1266),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1262),
.Y(n_1367)
);

CKINVDCx6p67_ASAP7_75t_R g1368 ( 
.A(n_1286),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1203),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1228),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1257),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1205),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1235),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1235),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1202),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1188),
.B(n_1313),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1299),
.B(n_1305),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1226),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1194),
.A2(n_1277),
.B1(n_1296),
.B2(n_1279),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1197),
.B(n_1225),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1193),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1252),
.B(n_1297),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1197),
.B(n_1258),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1294),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1241),
.A2(n_1312),
.B1(n_1305),
.B2(n_1210),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1210),
.A2(n_1264),
.B1(n_1261),
.B2(n_1297),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1267),
.A2(n_1250),
.B(n_1260),
.Y(n_1387)
);

BUFx4f_ASAP7_75t_SL g1388 ( 
.A(n_1211),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1191),
.A2(n_1206),
.B(n_1254),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1229),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1249),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1267),
.A2(n_1220),
.B(n_1293),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1297),
.A2(n_1265),
.B1(n_1263),
.B2(n_1249),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1263),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1249),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1244),
.Y(n_1396)
);

INVx6_ASAP7_75t_L g1397 ( 
.A(n_1298),
.Y(n_1397)
);

OAI21xp33_ASAP7_75t_L g1398 ( 
.A1(n_1265),
.A2(n_1269),
.B(n_1220),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1222),
.A2(n_1244),
.B1(n_1265),
.B2(n_1298),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1263),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1298),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1269),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1269),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1293),
.A2(n_1222),
.B1(n_1244),
.B2(n_1136),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1222),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1251),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1223),
.Y(n_1407)
);

AO21x1_ASAP7_75t_L g1408 ( 
.A1(n_1292),
.A2(n_1078),
.B(n_1056),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1251),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1184),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1188),
.B(n_1299),
.Y(n_1411)
);

CKINVDCx12_ASAP7_75t_R g1412 ( 
.A(n_1216),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1207),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1209),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1302),
.A2(n_1136),
.B1(n_1056),
.B2(n_1278),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1188),
.B(n_1299),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1236),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1302),
.A2(n_1136),
.B1(n_1056),
.B2(n_1278),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1278),
.B(n_1136),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1224),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1285),
.A2(n_1288),
.B1(n_1151),
.B2(n_1176),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1148),
.B2(n_1278),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1218),
.Y(n_1423)
);

BUFx2_ASAP7_75t_R g1424 ( 
.A(n_1237),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1209),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1215),
.B(n_1252),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1209),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1278),
.A2(n_755),
.B(n_1136),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1148),
.B2(n_1278),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1215),
.B(n_1252),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1236),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1251),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1215),
.B(n_1252),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1223),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1148),
.B2(n_1278),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1222),
.B(n_1191),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1223),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1184),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1223),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1222),
.B(n_1191),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1223),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1148),
.B2(n_1278),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1184),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1373),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1338),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1367),
.B(n_1365),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_L g1447 ( 
.A(n_1399),
.B(n_1331),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1316),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1374),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1351),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1333),
.B(n_1366),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1366),
.B(n_1346),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1382),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1422),
.A2(n_1435),
.B(n_1429),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1346),
.B(n_1355),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1316),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1411),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1332),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1341),
.Y(n_1459)
);

BUFx5_ASAP7_75t_L g1460 ( 
.A(n_1382),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1341),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1333),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1337),
.B(n_1317),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1382),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1317),
.B(n_1324),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1402),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1335),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1335),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1402),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1408),
.A2(n_1442),
.B1(n_1435),
.B2(n_1422),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1403),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1403),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1392),
.A2(n_1387),
.B(n_1400),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1363),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1345),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1325),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1355),
.B(n_1322),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1314),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1322),
.B(n_1426),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1383),
.A2(n_1398),
.B(n_1358),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1429),
.A2(n_1442),
.B1(n_1421),
.B2(n_1428),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1421),
.A2(n_1320),
.B1(n_1415),
.B2(n_1418),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1399),
.A2(n_1389),
.B(n_1319),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1358),
.A2(n_1393),
.B(n_1342),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1326),
.A2(n_1321),
.B(n_1319),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1417),
.Y(n_1486)
);

AND2x4_ASAP7_75t_SL g1487 ( 
.A(n_1404),
.B(n_1322),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1426),
.B(n_1430),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1426),
.B(n_1430),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1359),
.B(n_1386),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1347),
.B(n_1431),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1328),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1430),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1356),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1394),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1342),
.A2(n_1380),
.B(n_1360),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1362),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1433),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1318),
.Y(n_1499)
);

AO31x2_ASAP7_75t_L g1500 ( 
.A1(n_1336),
.A2(n_1443),
.A3(n_1323),
.B(n_1410),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1433),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1433),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1361),
.B(n_1376),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1328),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1416),
.B(n_1438),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1361),
.B(n_1344),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1369),
.B(n_1393),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1419),
.A2(n_1354),
.B(n_1385),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1372),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1345),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1343),
.A2(n_1350),
.B(n_1378),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1371),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1436),
.A2(n_1440),
.B(n_1441),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1405),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1396),
.Y(n_1515)
);

NOR2x1_ASAP7_75t_SL g1516 ( 
.A(n_1340),
.B(n_1434),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1379),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1436),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1339),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1379),
.A2(n_1395),
.B(n_1377),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1315),
.A2(n_1441),
.B(n_1349),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1327),
.B(n_1409),
.Y(n_1522)
);

AO21x1_ASAP7_75t_SL g1523 ( 
.A1(n_1401),
.A2(n_1439),
.B(n_1434),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1407),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1381),
.B(n_1406),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1444),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1473),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1413),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1511),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1511),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1413),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1454),
.A2(n_1384),
.B1(n_1375),
.B2(n_1381),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1496),
.B(n_1413),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1511),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1458),
.B(n_1445),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1448),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1525),
.Y(n_1539)
);

NOR2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1465),
.B(n_1368),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1481),
.A2(n_1391),
.B1(n_1424),
.B2(n_1353),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1449),
.B(n_1432),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1454),
.A2(n_1384),
.B1(n_1375),
.B2(n_1370),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1449),
.B(n_1328),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1453),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1449),
.B(n_1352),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1495),
.Y(n_1547)
);

NAND2x1_ASAP7_75t_L g1548 ( 
.A(n_1447),
.B(n_1364),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1482),
.A2(n_1412),
.B1(n_1353),
.B2(n_1370),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1452),
.B(n_1420),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1474),
.B(n_1420),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1474),
.B(n_1420),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1494),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1474),
.B(n_1352),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1446),
.B(n_1397),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1450),
.B(n_1401),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1485),
.A2(n_1414),
.B1(n_1329),
.B2(n_1348),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1478),
.B(n_1348),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1464),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1462),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1477),
.B(n_1391),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1477),
.B(n_1329),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1493),
.B(n_1357),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1466),
.B(n_1427),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1495),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1450),
.B(n_1388),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1466),
.B(n_1414),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1469),
.B(n_1357),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1469),
.B(n_1471),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1451),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1471),
.B(n_1425),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1451),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1456),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1472),
.B(n_1425),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1543),
.B(n_1508),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1540),
.A2(n_1485),
.B(n_1516),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1543),
.B(n_1508),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1476),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1534),
.A2(n_1470),
.B1(n_1447),
.B2(n_1490),
.Y(n_1580)
);

AOI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1541),
.A2(n_1517),
.B1(n_1463),
.B2(n_1457),
.C(n_1455),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1562),
.B(n_1522),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1557),
.A2(n_1490),
.B1(n_1455),
.B2(n_1501),
.Y(n_1583)
);

OAI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1557),
.A2(n_1517),
.B(n_1503),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1486),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1534),
.A2(n_1492),
.B1(n_1504),
.B2(n_1522),
.C(n_1507),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1553),
.B(n_1521),
.C(n_1514),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1538),
.B(n_1486),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1559),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1548),
.B(n_1507),
.C(n_1480),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1549),
.A2(n_1492),
.B1(n_1504),
.B2(n_1503),
.C(n_1526),
.Y(n_1591)
);

OAI21xp33_ASAP7_75t_L g1592 ( 
.A1(n_1549),
.A2(n_1497),
.B(n_1491),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1548),
.B(n_1480),
.C(n_1491),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1573),
.B(n_1520),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1530),
.B(n_1533),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1533),
.B(n_1479),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1533),
.B(n_1479),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1541),
.B(n_1480),
.C(n_1509),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_L g1599 ( 
.A(n_1556),
.B(n_1521),
.C(n_1524),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1520),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1535),
.B(n_1489),
.Y(n_1601)
);

OAI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1562),
.A2(n_1556),
.B1(n_1566),
.B2(n_1567),
.C(n_1537),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1537),
.B(n_1480),
.C(n_1484),
.Y(n_1603)
);

NAND4xp25_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1505),
.C(n_1514),
.D(n_1499),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1535),
.B(n_1575),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1561),
.A2(n_1487),
.B(n_1488),
.Y(n_1606)
);

NAND2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1540),
.B(n_1464),
.Y(n_1607)
);

AOI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1551),
.A2(n_1554),
.B(n_1552),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1460),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1570),
.B(n_1520),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1570),
.B(n_1520),
.Y(n_1611)
);

AND2x2_ASAP7_75t_SL g1612 ( 
.A(n_1559),
.B(n_1487),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1561),
.A2(n_1487),
.B(n_1488),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1571),
.A2(n_1519),
.B1(n_1505),
.B2(n_1506),
.C(n_1502),
.Y(n_1614)
);

NAND3xp33_ASAP7_75t_L g1615 ( 
.A(n_1551),
.B(n_1484),
.C(n_1515),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1572),
.B(n_1500),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1561),
.A2(n_1484),
.B1(n_1483),
.B2(n_1488),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1567),
.B(n_1483),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1575),
.B(n_1460),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1571),
.A2(n_1506),
.B1(n_1498),
.B2(n_1502),
.C(n_1512),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1551),
.A2(n_1554),
.B(n_1552),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1550),
.A2(n_1502),
.B1(n_1498),
.B2(n_1459),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1550),
.B(n_1460),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1550),
.B(n_1544),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1531),
.A2(n_1467),
.B(n_1468),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1528),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1563),
.B(n_1527),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1544),
.B(n_1500),
.Y(n_1628)
);

AND2x2_ASAP7_75t_SL g1629 ( 
.A(n_1559),
.B(n_1484),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1567),
.A2(n_1498),
.B1(n_1461),
.B2(n_1459),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1546),
.B(n_1555),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1552),
.B(n_1515),
.C(n_1518),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1558),
.B(n_1460),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1546),
.B(n_1500),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1558),
.B(n_1554),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1560),
.Y(n_1636)
);

NAND2x1_ASAP7_75t_L g1637 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1626),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1626),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1595),
.B(n_1531),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1625),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1595),
.B(n_1532),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1616),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1610),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1605),
.B(n_1532),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1611),
.B(n_1560),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1629),
.B(n_1536),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1629),
.B(n_1558),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1628),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1596),
.B(n_1529),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1589),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1596),
.B(n_1529),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1634),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1589),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_L g1656 ( 
.A(n_1587),
.B(n_1460),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1593),
.B(n_1590),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1545),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1597),
.B(n_1529),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1612),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1585),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1612),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1588),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1579),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1662),
.B(n_1582),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1640),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1640),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1666),
.B(n_1615),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1659),
.B(n_1609),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1638),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1648),
.B(n_1601),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1644),
.B(n_1601),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1661),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1659),
.B(n_1619),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1659),
.B(n_1619),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1599),
.Y(n_1679)
);

AND2x4_ASAP7_75t_SL g1680 ( 
.A(n_1661),
.B(n_1623),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1639),
.Y(n_1681)
);

NAND4xp25_ASAP7_75t_L g1682 ( 
.A(n_1658),
.B(n_1581),
.C(n_1598),
.D(n_1580),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1659),
.B(n_1651),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1652),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1658),
.A2(n_1578),
.B1(n_1576),
.B2(n_1583),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1641),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1659),
.B(n_1635),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1639),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1641),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.B(n_1633),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1666),
.B(n_1624),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1648),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1650),
.B(n_1617),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1637),
.B(n_1606),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1631),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1654),
.B(n_1547),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1661),
.B(n_1632),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1642),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1547),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1661),
.B(n_1607),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1641),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1643),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1651),
.B(n_1653),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1643),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1646),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1663),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1643),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1653),
.B(n_1623),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1653),
.B(n_1621),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1642),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1645),
.B(n_1565),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1660),
.B(n_1608),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1669),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1668),
.B(n_1686),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1680),
.B(n_1684),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1686),
.B(n_1679),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1669),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1685),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1670),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1670),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1682),
.A2(n_1656),
.B(n_1602),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1679),
.B(n_1682),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1706),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1671),
.B(n_1645),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1671),
.B(n_1662),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1676),
.B(n_1663),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1706),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1693),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1712),
.B(n_1664),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1673),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1660),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1680),
.B(n_1660),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1673),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1692),
.B(n_1636),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1685),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1692),
.B(n_1636),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1712),
.B(n_1664),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1676),
.B(n_1663),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1701),
.A2(n_1586),
.B(n_1618),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1674),
.B(n_1665),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1683),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1683),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1674),
.B(n_1665),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1685),
.Y(n_1745)
);

NAND2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1707),
.B(n_1637),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1707),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1693),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1697),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1697),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1695),
.Y(n_1752)
);

AOI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1694),
.A2(n_1591),
.B(n_1592),
.C(n_1584),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1694),
.Y(n_1754)
);

NAND2x1_ASAP7_75t_SL g1755 ( 
.A(n_1698),
.B(n_1649),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1695),
.A2(n_1657),
.B(n_1618),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1687),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1674),
.B(n_1649),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1696),
.B(n_1649),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1687),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1755),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1729),
.B(n_1700),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1745),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1723),
.B(n_1691),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1725),
.B(n_1726),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1539),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1725),
.B(n_1700),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1717),
.B(n_1691),
.Y(n_1768)
);

INVxp67_ASAP7_75t_SL g1769 ( 
.A(n_1755),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1714),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1675),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1735),
.B(n_1675),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1718),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1745),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1753),
.B(n_1584),
.C(n_1592),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1754),
.B(n_1691),
.Y(n_1776)
);

CKINVDCx16_ASAP7_75t_R g1777 ( 
.A(n_1722),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1747),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1740),
.A2(n_1695),
.B1(n_1746),
.B2(n_1752),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1716),
.B(n_1695),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1719),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1716),
.B(n_1695),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1727),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1720),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1735),
.B(n_1696),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1727),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1751),
.B(n_1713),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1752),
.A2(n_1695),
.B1(n_1698),
.B2(n_1607),
.Y(n_1789)
);

OA21x2_ASAP7_75t_L g1790 ( 
.A1(n_1756),
.A2(n_1681),
.B(n_1667),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1737),
.B(n_1647),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1727),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1721),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1732),
.B(n_1684),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1732),
.B(n_1672),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1733),
.B(n_1672),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1733),
.B(n_1739),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1739),
.B(n_1677),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1737),
.B(n_1647),
.Y(n_1799)
);

AOI222xp33_ASAP7_75t_L g1800 ( 
.A1(n_1775),
.A2(n_1739),
.B1(n_1698),
.B2(n_1724),
.C1(n_1728),
.C2(n_1758),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1770),
.Y(n_1801)
);

NOR2xp67_ASAP7_75t_L g1802 ( 
.A(n_1779),
.B(n_1719),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1770),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1777),
.B(n_1746),
.Y(n_1804)
);

OAI211xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1777),
.A2(n_1734),
.B(n_1742),
.C(n_1731),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1761),
.A2(n_1743),
.B1(n_1738),
.B2(n_1730),
.C(n_1736),
.Y(n_1806)
);

OAI211xp5_ASAP7_75t_SL g1807 ( 
.A1(n_1783),
.A2(n_1736),
.B(n_1759),
.C(n_1744),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1794),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1773),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1778),
.B(n_1741),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1773),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1769),
.A2(n_1698),
.B(n_1657),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1794),
.Y(n_1813)
);

OAI31xp33_ASAP7_75t_L g1814 ( 
.A1(n_1787),
.A2(n_1757),
.A3(n_1760),
.B(n_1614),
.Y(n_1814)
);

NAND2xp33_ASAP7_75t_SL g1815 ( 
.A(n_1768),
.B(n_1710),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1784),
.Y(n_1816)
);

AOI21xp33_ASAP7_75t_L g1817 ( 
.A1(n_1792),
.A2(n_1749),
.B(n_1566),
.Y(n_1817)
);

AOI221x1_ASAP7_75t_L g1818 ( 
.A1(n_1763),
.A2(n_1749),
.B1(n_1604),
.B2(n_1711),
.C(n_1710),
.Y(n_1818)
);

O2A1O1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1764),
.A2(n_1766),
.B(n_1774),
.C(n_1763),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1784),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1789),
.A2(n_1620),
.B1(n_1630),
.B2(n_1677),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1797),
.B(n_1678),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1793),
.Y(n_1823)
);

AOI222xp33_ASAP7_75t_L g1824 ( 
.A1(n_1776),
.A2(n_1574),
.B1(n_1568),
.B2(n_1564),
.C1(n_1690),
.C2(n_1702),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1795),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1780),
.A2(n_1563),
.B1(n_1678),
.B2(n_1704),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1797),
.A2(n_1704),
.B1(n_1690),
.B2(n_1703),
.Y(n_1827)
);

OAI31xp33_ASAP7_75t_L g1828 ( 
.A1(n_1780),
.A2(n_1613),
.A3(n_1574),
.B(n_1652),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1798),
.B(n_1688),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1808),
.B(n_1774),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1825),
.B(n_1765),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1801),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1803),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1804),
.B(n_1782),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1804),
.B(n_1765),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1822),
.B(n_1798),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1822),
.B(n_1782),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1800),
.B(n_1795),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1809),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1825),
.B(n_1796),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1808),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1813),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1829),
.B(n_1813),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1810),
.B(n_1762),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1829),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1811),
.Y(n_1846)
);

NAND2x1_ASAP7_75t_L g1847 ( 
.A(n_1802),
.B(n_1790),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1826),
.B(n_1796),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1816),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1820),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1812),
.B(n_1781),
.Y(n_1851)
);

AND4x1_ASAP7_75t_L g1852 ( 
.A(n_1834),
.B(n_1819),
.C(n_1814),
.D(n_1818),
.Y(n_1852)
);

O2A1O1Ixp33_ASAP7_75t_SL g1853 ( 
.A1(n_1847),
.A2(n_1805),
.B(n_1806),
.C(n_1807),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1838),
.A2(n_1821),
.B1(n_1785),
.B2(n_1788),
.Y(n_1854)
);

NOR3x1_ASAP7_75t_L g1855 ( 
.A(n_1835),
.B(n_1823),
.C(n_1762),
.Y(n_1855)
);

OAI211xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1844),
.A2(n_1828),
.B(n_1824),
.C(n_1817),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1847),
.A2(n_1815),
.B(n_1818),
.C(n_1767),
.Y(n_1857)
);

OAI211xp5_ASAP7_75t_SL g1858 ( 
.A1(n_1844),
.A2(n_1781),
.B(n_1767),
.C(n_1793),
.Y(n_1858)
);

NAND4xp75_ASAP7_75t_L g1859 ( 
.A(n_1842),
.B(n_1790),
.C(n_1815),
.D(n_1334),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_L g1860 ( 
.A(n_1851),
.B(n_1827),
.C(n_1771),
.Y(n_1860)
);

NOR4xp25_ASAP7_75t_L g1861 ( 
.A(n_1839),
.B(n_1771),
.C(n_1786),
.D(n_1772),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1843),
.B(n_1786),
.Y(n_1862)
);

NOR3xp33_ASAP7_75t_SL g1863 ( 
.A(n_1840),
.B(n_1627),
.C(n_1790),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1851),
.A2(n_1772),
.B1(n_1791),
.B2(n_1799),
.C(n_1711),
.Y(n_1864)
);

NAND4xp25_ASAP7_75t_SL g1865 ( 
.A(n_1848),
.B(n_1791),
.C(n_1799),
.D(n_1574),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1837),
.B(n_1688),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1862),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1852),
.B(n_1846),
.C(n_1839),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_1865),
.B(n_1842),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1858),
.Y(n_1870)
);

NOR3x1_ASAP7_75t_L g1871 ( 
.A(n_1859),
.B(n_1833),
.C(n_1832),
.Y(n_1871)
);

NOR3xp33_ASAP7_75t_L g1872 ( 
.A(n_1854),
.B(n_1850),
.C(n_1841),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1855),
.Y(n_1873)
);

NAND2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1866),
.B(n_1831),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1856),
.B(n_1831),
.Y(n_1875)
);

NOR3xp33_ASAP7_75t_L g1876 ( 
.A(n_1853),
.B(n_1860),
.C(n_1857),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1861),
.Y(n_1877)
);

NOR3x1_ASAP7_75t_L g1878 ( 
.A(n_1863),
.B(n_1849),
.C(n_1846),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1864),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1861),
.B(n_1843),
.Y(n_1880)
);

NOR2xp67_ASAP7_75t_L g1881 ( 
.A(n_1865),
.B(n_1845),
.Y(n_1881)
);

OAI211xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1876),
.A2(n_1849),
.B(n_1841),
.C(n_1845),
.Y(n_1882)
);

AOI21xp33_ASAP7_75t_L g1883 ( 
.A1(n_1877),
.A2(n_1830),
.B(n_1848),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1875),
.A2(n_1830),
.B1(n_1837),
.B2(n_1836),
.C(n_1564),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1874),
.A2(n_1836),
.B(n_1830),
.Y(n_1885)
);

NAND4xp75_ASAP7_75t_L g1886 ( 
.A(n_1871),
.B(n_1790),
.C(n_1330),
.D(n_1568),
.Y(n_1886)
);

AOI211xp5_ASAP7_75t_L g1887 ( 
.A1(n_1868),
.A2(n_1568),
.B(n_1564),
.C(n_1566),
.Y(n_1887)
);

OAI211xp5_ASAP7_75t_L g1888 ( 
.A1(n_1880),
.A2(n_1868),
.B(n_1870),
.C(n_1873),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1869),
.A2(n_1881),
.B(n_1872),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1888),
.A2(n_1879),
.B1(n_1867),
.B2(n_1878),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1885),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1882),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1887),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1884),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1886),
.Y(n_1895)
);

AO22x1_ASAP7_75t_L g1896 ( 
.A1(n_1889),
.A2(n_1711),
.B1(n_1667),
.B2(n_1689),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1883),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1891),
.Y(n_1898)
);

OAI21xp33_ASAP7_75t_L g1899 ( 
.A1(n_1890),
.A2(n_1893),
.B(n_1895),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1897),
.Y(n_1900)
);

NOR3xp33_ASAP7_75t_L g1901 ( 
.A(n_1892),
.B(n_1388),
.C(n_1563),
.Y(n_1901)
);

NOR2x1p5_ASAP7_75t_L g1902 ( 
.A(n_1894),
.B(n_1475),
.Y(n_1902)
);

NAND4xp75_ASAP7_75t_L g1903 ( 
.A(n_1896),
.B(n_1681),
.C(n_1689),
.D(n_1667),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1890),
.A2(n_1681),
.B1(n_1699),
.B2(n_1689),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1903),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1898),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1902),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1906),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1908),
.Y(n_1909)
);

OA22x2_ASAP7_75t_L g1910 ( 
.A1(n_1909),
.A2(n_1899),
.B1(n_1900),
.B2(n_1905),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1909),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1910),
.A2(n_1907),
.B(n_1905),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1911),
.Y(n_1913)
);

AOI21xp33_ASAP7_75t_SL g1914 ( 
.A1(n_1912),
.A2(n_1901),
.B(n_1904),
.Y(n_1914)
);

AOI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1913),
.A2(n_1699),
.B1(n_1655),
.B2(n_1708),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1914),
.A2(n_1699),
.B(n_1709),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1915),
.B1(n_1705),
.B2(n_1708),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_R g1918 ( 
.A1(n_1917),
.A2(n_1622),
.B1(n_1523),
.B2(n_1655),
.C(n_1516),
.Y(n_1918)
);

AOI211xp5_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1510),
.B(n_1527),
.C(n_1513),
.Y(n_1919)
);


endmodule