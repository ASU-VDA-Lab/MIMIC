module fake_jpeg_6119_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_22),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_50),
.B1(n_68),
.B2(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_29),
.C(n_28),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_17),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_74),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_78),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_16),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_35),
.B(n_17),
.C(n_34),
.Y(n_95)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_88),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_44),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_44),
.C(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_37),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_31),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_85),
.B(n_89),
.Y(n_132)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_101),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_19),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_64),
.B1(n_46),
.B2(n_41),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_83),
.B1(n_84),
.B2(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_44),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_104),
.Y(n_130)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_46),
.B1(n_60),
.B2(n_32),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_44),
.C(n_39),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_44),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_83),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_107),
.B1(n_94),
.B2(n_92),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_129),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_71),
.B1(n_81),
.B2(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_138),
.B(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_77),
.B1(n_90),
.B2(n_80),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_22),
.B1(n_45),
.B2(n_49),
.Y(n_167)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_104),
.C(n_99),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_93),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_33),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_95),
.B(n_34),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_32),
.B(n_33),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_60),
.B1(n_45),
.B2(n_62),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_130),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_98),
.B(n_111),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_154),
.B(n_159),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_148),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_133),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_158),
.C(n_162),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_15),
.C(n_2),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_108),
.B(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_30),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_97),
.B(n_39),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_105),
.B1(n_19),
.B2(n_25),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_130),
.B(n_122),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_39),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_39),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_168),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_31),
.B(n_39),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_118),
.B1(n_123),
.B2(n_125),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_129),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_22),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_136),
.B1(n_139),
.B2(n_138),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_181),
.B1(n_187),
.B2(n_160),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_136),
.B1(n_140),
.B2(n_118),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_117),
.B1(n_124),
.B2(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_165),
.B(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_22),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_49),
.B1(n_57),
.B2(n_56),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_194),
.C(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_61),
.B1(n_18),
.B2(n_22),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_18),
.B1(n_30),
.B2(n_21),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_193),
.B1(n_176),
.B2(n_179),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_23),
.B1(n_21),
.B2(n_3),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_1),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_168),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_199),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_149),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_204),
.C(n_207),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_163),
.C(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_164),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_216),
.C(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_157),
.B1(n_155),
.B2(n_23),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_23),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_226),
.C(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_208),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

HAxp5_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_189),
.CON(n_225),
.SN(n_225)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_204),
.C(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_180),
.C(n_172),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_230),
.B(n_23),
.Y(n_244)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_232),
.B1(n_214),
.B2(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_181),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_243),
.C(n_245),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_201),
.C(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_247),
.C(n_235),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_241),
.B(n_244),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_242),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_229),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_218),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_23),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_21),
.C(n_2),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_217),
.B(n_220),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_240),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_220),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_255),
.B(n_257),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_228),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_233),
.C(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_266),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_219),
.B1(n_234),
.B2(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_269),
.C(n_21),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_3),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_263),
.B1(n_265),
.B2(n_269),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_21),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_267),
.A2(n_256),
.B1(n_253),
.B2(n_6),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_272),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_4),
.B(n_5),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_7),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_13),
.B(n_6),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_5),
.C(n_6),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_276),
.A2(n_5),
.B(n_7),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_279),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_276),
.B(n_275),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_284),
.A2(n_280),
.B(n_9),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_283),
.B(n_12),
.C(n_13),
.D(n_8),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_285),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_12),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_12),
.C(n_13),
.Y(n_290)
);


endmodule