module fake_netlist_6_4503_n_284 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_44, n_284);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_44;

output n_284;

wire n_52;
wire n_91;
wire n_119;
wire n_146;
wire n_163;
wire n_235;
wire n_256;
wire n_193;
wire n_269;
wire n_147;
wire n_258;
wire n_281;
wire n_154;
wire n_191;
wire n_88;
wire n_209;
wire n_98;
wire n_277;
wire n_260;
wire n_265;
wire n_283;
wire n_113;
wire n_63;
wire n_223;
wire n_278;
wire n_270;
wire n_73;
wire n_279;
wire n_148;
wire n_199;
wire n_226;
wire n_161;
wire n_138;
wire n_208;
wire n_68;
wire n_228;
wire n_252;
wire n_266;
wire n_166;
wire n_184;
wire n_212;
wire n_268;
wire n_271;
wire n_50;
wire n_158;
wire n_210;
wire n_217;
wire n_83;
wire n_206;
wire n_216;
wire n_221;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_227;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_261;
wire n_189;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_130;
wire n_213;
wire n_164;
wire n_257;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_254;
wire n_142;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_62;
wire n_155;
wire n_219;
wire n_75;
wire n_109;
wire n_150;
wire n_233;
wire n_264;
wire n_122;
wire n_263;
wire n_255;
wire n_205;
wire n_140;
wire n_218;
wire n_70;
wire n_120;
wire n_234;
wire n_251;
wire n_214;
wire n_274;
wire n_67;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_237;
wire n_81;
wire n_59;
wire n_244;
wire n_181;
wire n_76;
wire n_182;
wire n_124;
wire n_243;
wire n_238;
wire n_239;
wire n_55;
wire n_126;
wire n_202;
wire n_97;
wire n_94;
wire n_108;
wire n_267;
wire n_282;
wire n_58;
wire n_116;
wire n_280;
wire n_211;
wire n_64;
wire n_220;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_65;
wire n_230;
wire n_93;
wire n_80;
wire n_141;
wire n_240;
wire n_135;
wire n_200;
wire n_196;
wire n_165;
wire n_139;
wire n_134;
wire n_259;
wire n_177;
wire n_176;
wire n_273;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_248;
wire n_107;
wire n_71;
wire n_74;
wire n_229;
wire n_253;
wire n_190;
wire n_123;
wire n_262;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_249;
wire n_173;
wire n_201;
wire n_250;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_272;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_241;
wire n_79;
wire n_275;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_276;
wire n_51;
wire n_56;
wire n_232;

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_25),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_7),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_39),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_15),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_0),
.B(n_1),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_1),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_3),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_56),
.B1(n_58),
.B2(n_69),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_101),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_90),
.B1(n_101),
.B2(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_69),
.C(n_67),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_36),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_31),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_115),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_87),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_119),
.A3(n_117),
.B1(n_114),
.B2(n_112),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_94),
.Y(n_140)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_86),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_96),
.Y(n_147)
);

OR2x6_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_113),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_85),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2x1_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_133),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_122),
.B1(n_129),
.B2(n_88),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_124),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_110),
.B(n_118),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2x1_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_110),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

OR2x6_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_95),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_92),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_143),
.B(n_142),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_143),
.B(n_144),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g176 ( 
.A(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_140),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_165),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_140),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_150),
.B(n_159),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

OA222x2_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_164),
.B1(n_151),
.B2(n_148),
.C1(n_138),
.C2(n_85),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_154),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_153),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_182),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_188),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_180),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_169),
.B(n_170),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_178),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_169),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_178),
.Y(n_215)
);

AOI211x1_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_184),
.B(n_155),
.C(n_176),
.Y(n_216)
);

AO21x2_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_169),
.B(n_181),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_195),
.Y(n_220)
);

AOI33xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_197),
.A3(n_92),
.B1(n_95),
.B2(n_201),
.B3(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_203),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NAND2x1p5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AND2x4_ASAP7_75t_SL g239 ( 
.A(n_220),
.B(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_199),
.Y(n_240)
);

OR2x4_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_93),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_217),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_218),
.Y(n_244)
);

NOR2x1p5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_231),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_199),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_243),
.B(n_221),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_221),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_226),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_239),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_246),
.B1(n_241),
.B2(n_242),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_246),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_253),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_251),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_259),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_263),
.C(n_250),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_249),
.B1(n_257),
.B2(n_265),
.Y(n_271)
);

AOI211xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_257),
.B(n_264),
.C(n_238),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_271),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_181),
.C(n_150),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_4),
.Y(n_275)
);

OAI222xp33_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_181),
.B1(n_150),
.B2(n_185),
.C1(n_205),
.C2(n_23),
.Y(n_276)
);

OAI322xp33_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_10),
.A3(n_12),
.B1(n_18),
.B2(n_21),
.C1(n_26),
.C2(n_27),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

OAI22x1_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_185),
.B1(n_176),
.B2(n_38),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_185),
.B1(n_139),
.B2(n_40),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_163),
.B(n_46),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

AOI221xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_282),
.B1(n_277),
.B2(n_280),
.C(n_48),
.Y(n_284)
);


endmodule