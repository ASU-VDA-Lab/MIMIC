module fake_jpeg_3479_n_63 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_63);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_19),
.B1(n_23),
.B2(n_18),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_22),
.B(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_22),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_20),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_28),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_29),
.B1(n_33),
.B2(n_28),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_38),
.B1(n_21),
.B2(n_20),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_23),
.C(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_36),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_47),
.B(n_13),
.Y(n_55)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_36),
.B1(n_38),
.B2(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_38),
.B1(n_45),
.B2(n_40),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_55),
.B(n_4),
.C(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_48),
.B(n_51),
.Y(n_56)
);

AOI321xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.A3(n_58),
.B1(n_55),
.B2(n_6),
.C(n_7),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_12),
.C(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_5),
.Y(n_60)
);

NOR4xp25_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_9),
.Y(n_63)
);


endmodule