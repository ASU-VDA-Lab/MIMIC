module real_aes_6671_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g427 ( .A(n_0), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_1), .A2(n_125), .B(n_128), .C(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g132 ( .A(n_2), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_3), .A2(n_148), .B(n_526), .Y(n_525) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_4), .A2(n_103), .B1(n_705), .B2(n_708), .C1(n_711), .C2(n_712), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_5), .B(n_160), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_6), .A2(n_148), .B(n_177), .Y(n_176) );
AND2x6_ASAP7_75t_L g125 ( .A(n_7), .B(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_8), .A2(n_230), .B(n_231), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_9), .B(n_40), .Y(n_428) );
INVx1_ASAP7_75t_L g469 ( .A(n_10), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_11), .B(n_136), .Y(n_504) );
INVx1_ASAP7_75t_L g182 ( .A(n_12), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_13), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g117 ( .A(n_14), .Y(n_117) );
INVx1_ASAP7_75t_L g236 ( .A(n_15), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_16), .A2(n_134), .B(n_237), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_17), .B(n_160), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_18), .B(n_153), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_19), .B(n_148), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_20), .B(n_461), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_21), .A2(n_138), .B(n_211), .C(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_22), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_23), .B(n_136), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_24), .A2(n_234), .B(n_235), .C(n_237), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_25), .B(n_136), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_26), .Y(n_516) );
INVx1_ASAP7_75t_L g440 ( .A(n_27), .Y(n_440) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_28), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_29), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_30), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g457 ( .A(n_31), .Y(n_457) );
INVx1_ASAP7_75t_L g171 ( .A(n_32), .Y(n_171) );
INVx2_ASAP7_75t_L g123 ( .A(n_33), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_34), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_35), .A2(n_156), .B(n_211), .C(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g458 ( .A(n_36), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_37), .A2(n_125), .B(n_128), .C(n_195), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_38), .A2(n_128), .B(n_439), .C(n_444), .Y(n_438) );
CKINVDCx14_ASAP7_75t_R g527 ( .A(n_39), .Y(n_527) );
INVx1_ASAP7_75t_L g169 ( .A(n_41), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_42), .A2(n_180), .B(n_199), .C(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_43), .B(n_136), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_44), .A2(n_47), .B1(n_726), .B2(n_727), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_44), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_45), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_46), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_47), .A2(n_101), .B1(n_714), .B2(n_723), .C1(n_733), .C2(n_739), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_47), .Y(n_726) );
INVx1_ASAP7_75t_L g476 ( .A(n_48), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_49), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_50), .B(n_148), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_51), .A2(n_128), .B1(n_138), .B2(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_52), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_53), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_54), .A2(n_156), .B(n_180), .C(n_181), .Y(n_179) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_55), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_56), .Y(n_227) );
INVx1_ASAP7_75t_L g178 ( .A(n_57), .Y(n_178) );
INVx1_ASAP7_75t_L g126 ( .A(n_58), .Y(n_126) );
INVx1_ASAP7_75t_L g116 ( .A(n_59), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_60), .A2(n_89), .B1(n_706), .B2(n_707), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_60), .Y(n_706) );
INVx1_ASAP7_75t_SL g530 ( .A(n_61), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_62), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_63), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_64), .B(n_160), .Y(n_480) );
INVx1_ASAP7_75t_L g519 ( .A(n_65), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_SL g152 ( .A1(n_66), .A2(n_153), .B(n_154), .C(n_156), .Y(n_152) );
INVxp67_ASAP7_75t_L g155 ( .A(n_67), .Y(n_155) );
INVx1_ASAP7_75t_L g718 ( .A(n_68), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_69), .A2(n_148), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_70), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_71), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_72), .A2(n_148), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g220 ( .A(n_73), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_74), .A2(n_230), .B(n_453), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_75), .Y(n_437) );
INVx1_ASAP7_75t_L g486 ( .A(n_76), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_77), .A2(n_125), .B(n_128), .C(n_222), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_78), .A2(n_148), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g489 ( .A(n_79), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_80), .B(n_133), .Y(n_196) );
INVx2_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
INVx1_ASAP7_75t_L g502 ( .A(n_82), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_83), .B(n_153), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g127 ( .A1(n_84), .A2(n_125), .B(n_128), .C(n_131), .Y(n_127) );
INVx2_ASAP7_75t_L g425 ( .A(n_85), .Y(n_425) );
OR2x2_ASAP7_75t_L g704 ( .A(n_85), .B(n_426), .Y(n_704) );
OR2x2_ASAP7_75t_L g722 ( .A(n_85), .B(n_713), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_86), .A2(n_128), .B(n_518), .C(n_521), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_87), .B(n_143), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_88), .Y(n_141) );
CKINVDCx14_ASAP7_75t_R g707 ( .A(n_89), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_90), .A2(n_125), .B(n_128), .C(n_208), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_91), .Y(n_215) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_93), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_94), .B(n_133), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_95), .B(n_146), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_96), .B(n_146), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_97), .A2(n_148), .B(n_149), .Y(n_147) );
INVx2_ASAP7_75t_L g479 ( .A(n_98), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_99), .B(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_422), .B1(n_429), .B2(n_704), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_105), .A2(n_422), .B1(n_430), .B2(n_709), .Y(n_708) );
OR4x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_311), .C(n_371), .D(n_398), .Y(n_105) );
NAND4xp25_ASAP7_75t_SL g106 ( .A(n_107), .B(n_259), .C(n_290), .D(n_307), .Y(n_106) );
O2A1O1Ixp33_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_184), .B(n_186), .C(n_239), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_162), .Y(n_108) );
INVx1_ASAP7_75t_L g301 ( .A(n_109), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_109), .A2(n_342), .B1(n_390), .B2(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_144), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_110), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g252 ( .A(n_110), .B(n_164), .Y(n_252) );
AND2x2_ASAP7_75t_L g294 ( .A(n_110), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_110), .B(n_185), .Y(n_306) );
INVx1_ASAP7_75t_L g346 ( .A(n_110), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_110), .B(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g274 ( .A(n_111), .B(n_164), .Y(n_274) );
INVx3_ASAP7_75t_L g278 ( .A(n_111), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_111), .B(n_336), .Y(n_335) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_118), .B(n_140), .Y(n_111) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_112), .A2(n_165), .B(n_173), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_112), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g201 ( .A(n_112), .Y(n_201) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_113), .Y(n_146) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_114), .B(n_115), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B(n_127), .Y(n_118) );
OAI22xp33_ASAP7_75t_L g165 ( .A1(n_120), .A2(n_158), .B1(n_166), .B2(n_172), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_120), .A2(n_220), .B(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g436 ( .A1(n_120), .A2(n_143), .B(n_437), .C(n_438), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_120), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_120), .A2(n_516), .B(n_517), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_125), .Y(n_120) );
AND2x4_ASAP7_75t_L g148 ( .A(n_121), .B(n_125), .Y(n_148) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g443 ( .A(n_122), .Y(n_443) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g129 ( .A(n_123), .Y(n_129) );
INVx1_ASAP7_75t_L g139 ( .A(n_123), .Y(n_139) );
INVx1_ASAP7_75t_L g130 ( .A(n_124), .Y(n_130) );
INVx3_ASAP7_75t_L g134 ( .A(n_124), .Y(n_134) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_124), .Y(n_136) );
INVx1_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
INVx4_ASAP7_75t_SL g158 ( .A(n_125), .Y(n_158) );
BUFx3_ASAP7_75t_L g444 ( .A(n_125), .Y(n_444) );
INVx5_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
AND2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
BUFx3_ASAP7_75t_L g200 ( .A(n_129), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_135), .C(n_137), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_133), .A2(n_440), .B(n_441), .C(n_442), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_133), .A2(n_234), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_134), .B(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_134), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_134), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
INVx4_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_142), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_142), .B(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_142), .A2(n_498), .B(n_505), .Y(n_497) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_143), .A2(n_229), .B(n_238), .Y(n_228) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_143), .A2(n_464), .B(n_470), .Y(n_463) );
AND2x2_ASAP7_75t_L g365 ( .A(n_144), .B(n_175), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_144), .B(n_278), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_144), .B(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g185 ( .A(n_145), .B(n_164), .Y(n_185) );
INVx1_ASAP7_75t_L g247 ( .A(n_145), .Y(n_247) );
BUFx2_ASAP7_75t_L g251 ( .A(n_145), .Y(n_251) );
AND2x2_ASAP7_75t_L g295 ( .A(n_145), .B(n_163), .Y(n_295) );
OR2x2_ASAP7_75t_L g334 ( .A(n_145), .B(n_163), .Y(n_334) );
AND2x2_ASAP7_75t_L g359 ( .A(n_145), .B(n_175), .Y(n_359) );
AND2x2_ASAP7_75t_L g418 ( .A(n_145), .B(n_248), .Y(n_418) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_159), .Y(n_145) );
INVx4_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_146), .Y(n_473) );
BUFx2_ASAP7_75t_L g230 ( .A(n_148), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_152), .C(n_158), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_150), .A2(n_158), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_150), .A2(n_158), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g453 ( .A1(n_150), .A2(n_158), .B(n_454), .C(n_455), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_150), .A2(n_158), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_150), .A2(n_158), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_150), .A2(n_158), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_150), .A2(n_158), .B(n_527), .C(n_528), .Y(n_526) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
INVx1_ASAP7_75t_L g521 ( .A(n_158), .Y(n_521) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_160), .A2(n_176), .B(n_183), .Y(n_175) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_161), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_161), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_161), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_161), .A2(n_515), .B(n_522), .Y(n_514) );
INVx1_ASAP7_75t_L g393 ( .A(n_162), .Y(n_393) );
OR2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_175), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_163), .B(n_175), .Y(n_279) );
AND2x2_ASAP7_75t_L g289 ( .A(n_163), .B(n_278), .Y(n_289) );
BUFx2_ASAP7_75t_L g300 ( .A(n_163), .Y(n_300) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g322 ( .A(n_164), .B(n_175), .Y(n_322) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_164), .Y(n_377) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_167) );
INVx2_ASAP7_75t_L g170 ( .A(n_168), .Y(n_170) );
INVx4_ASAP7_75t_L g234 ( .A(n_168), .Y(n_234) );
INVx2_ASAP7_75t_L g503 ( .A(n_170), .Y(n_503) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_175), .B(n_185), .Y(n_184) );
INVx1_ASAP7_75t_SL g248 ( .A(n_175), .Y(n_248) );
BUFx2_ASAP7_75t_L g273 ( .A(n_175), .Y(n_273) );
INVx2_ASAP7_75t_L g292 ( .A(n_175), .Y(n_292) );
AND2x2_ASAP7_75t_L g354 ( .A(n_175), .B(n_278), .Y(n_354) );
AOI321xp33_ASAP7_75t_L g373 ( .A1(n_184), .A2(n_374), .A3(n_375), .B1(n_376), .B2(n_378), .C(n_379), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_185), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_185), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g367 ( .A(n_185), .B(n_346), .Y(n_367) );
AND2x2_ASAP7_75t_L g400 ( .A(n_185), .B(n_292), .Y(n_400) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_216), .Y(n_187) );
OR2x2_ASAP7_75t_L g302 ( .A(n_188), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_204), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g254 ( .A(n_191), .Y(n_254) );
AND2x2_ASAP7_75t_L g264 ( .A(n_191), .B(n_218), .Y(n_264) );
AND2x2_ASAP7_75t_L g269 ( .A(n_191), .B(n_244), .Y(n_269) );
INVx1_ASAP7_75t_L g286 ( .A(n_191), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_191), .B(n_267), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_191), .B(n_243), .Y(n_310) );
OR2x2_ASAP7_75t_L g342 ( .A(n_191), .B(n_331), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_191), .B(n_255), .Y(n_381) );
AND2x2_ASAP7_75t_L g415 ( .A(n_191), .B(n_241), .Y(n_415) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
AOI21xp5_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_194), .B(n_201), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_198), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp5_ASAP7_75t_L g501 ( .A1(n_198), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_198), .A2(n_503), .B(n_519), .C(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
INVx1_ASAP7_75t_L g225 ( .A(n_201), .Y(n_225) );
INVx1_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
INVx2_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
AND2x2_ASAP7_75t_L g297 ( .A(n_204), .B(n_268), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_204), .B(n_244), .Y(n_319) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_214), .Y(n_204) );
INVx1_ASAP7_75t_L g461 ( .A(n_205), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_205), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_213), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_212), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_211), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g403 ( .A(n_217), .B(n_254), .Y(n_403) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_228), .Y(n_217) );
INVx2_ASAP7_75t_L g244 ( .A(n_218), .Y(n_244) );
AND2x2_ASAP7_75t_L g397 ( .A(n_218), .B(n_257), .Y(n_397) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_225), .B(n_226), .Y(n_218) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_225), .A2(n_451), .B(n_459), .Y(n_450) );
INVx1_ASAP7_75t_L g549 ( .A(n_225), .Y(n_549) );
AND2x2_ASAP7_75t_L g243 ( .A(n_228), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g258 ( .A(n_228), .Y(n_258) );
INVx1_ASAP7_75t_L g268 ( .A(n_228), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_234), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_234), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_234), .B(n_489), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_245), .B1(n_249), .B2(n_253), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_240), .A2(n_358), .B1(n_395), .B2(n_396), .Y(n_394) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_243), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_244), .B(n_257), .Y(n_331) );
INVx1_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
AND2x2_ASAP7_75t_L g288 ( .A(n_246), .B(n_289), .Y(n_288) );
INVx3_ASAP7_75t_SL g327 ( .A(n_246), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_246), .B(n_252), .Y(n_404) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g413 ( .A(n_249), .Y(n_413) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_250), .B(n_346), .Y(n_388) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_SL g293 ( .A(n_252), .Y(n_293) );
NAND2x1_ASAP7_75t_SL g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g314 ( .A(n_254), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g321 ( .A(n_254), .B(n_258), .Y(n_321) );
AND2x2_ASAP7_75t_L g326 ( .A(n_254), .B(n_267), .Y(n_326) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_254), .Y(n_375) );
OAI311xp33_ASAP7_75t_L g398 ( .A1(n_255), .A2(n_399), .A3(n_401), .B1(n_402), .C1(n_412), .Y(n_398) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g411 ( .A(n_256), .B(n_284), .Y(n_411) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g267 ( .A(n_257), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g315 ( .A(n_257), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g370 ( .A(n_257), .Y(n_370) );
INVx1_ASAP7_75t_L g263 ( .A(n_258), .Y(n_263) );
INVx1_ASAP7_75t_L g283 ( .A(n_258), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_258), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
AOI221xp5_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_262), .B1(n_270), .B2(n_275), .C(n_280), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx4_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
AND2x2_ASAP7_75t_L g378 ( .A(n_264), .B(n_297), .Y(n_378) );
AND2x2_ASAP7_75t_L g385 ( .A(n_264), .B(n_267), .Y(n_385) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_267), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g296 ( .A(n_269), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_272), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g421 ( .A(n_274), .B(n_365), .Y(n_421) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g406 ( .A(n_278), .B(n_334), .Y(n_406) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_279), .A2(n_372), .B(n_373), .C(n_386), .Y(n_371) );
AOI21xp33_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_285), .B(n_287), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp67_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g350 ( .A(n_284), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_285), .A2(n_380), .B1(n_381), .B2(n_382), .C(n_383), .Y(n_379) );
AND2x2_ASAP7_75t_L g356 ( .A(n_286), .B(n_297), .Y(n_356) );
AND2x2_ASAP7_75t_L g409 ( .A(n_286), .B(n_304), .Y(n_409) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_289), .B(n_327), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_294), .B(n_296), .C(n_298), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g337 ( .A(n_292), .B(n_295), .Y(n_337) );
OR2x2_ASAP7_75t_L g380 ( .A(n_292), .B(n_334), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_293), .B(n_359), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_293), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g324 ( .A(n_294), .Y(n_324) );
INVx1_ASAP7_75t_L g390 ( .A(n_297), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_305), .B2(n_306), .Y(n_298) );
INVx1_ASAP7_75t_L g313 ( .A(n_299), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_300), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g376 ( .A(n_301), .B(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g362 ( .A(n_303), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_304), .B(n_390), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_305), .A2(n_364), .B1(n_366), .B2(n_368), .Y(n_363) );
INVx1_ASAP7_75t_L g372 ( .A(n_308), .Y(n_372) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g414 ( .A(n_309), .B(n_409), .Y(n_414) );
AOI222xp33_ASAP7_75t_L g343 ( .A1(n_310), .A2(n_344), .B1(n_347), .B2(n_348), .C1(n_351), .C2(n_352), .Y(n_343) );
NAND4xp25_ASAP7_75t_SL g311 ( .A(n_312), .B(n_332), .C(n_343), .D(n_355), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_317), .B2(n_322), .C(n_323), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_315), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g341 ( .A(n_316), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_317), .A2(n_387), .B1(n_389), .B2(n_391), .C(n_394), .Y(n_386) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g329 ( .A(n_321), .B(n_330), .Y(n_329) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_322), .A2(n_384), .B(n_385), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_327), .B2(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_338), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g374 ( .A(n_345), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_346), .B(n_365), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_346), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_350), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g382 ( .A(n_354), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_360), .B2(n_362), .C(n_363), .Y(n_355) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI222xp33_ASAP7_75t_L g402 ( .A1(n_365), .A2(n_403), .B1(n_404), .B2(n_405), .C1(n_407), .C2(n_410), .Y(n_402) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_369), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g401 ( .A(n_375), .Y(n_401) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp33_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_415), .B2(n_416), .C(n_419), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NOR2x2_ASAP7_75t_L g712 ( .A(n_425), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_426), .Y(n_713) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_430), .B(n_725), .Y(n_724) );
OR5x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_598), .C(n_662), .D(n_678), .E(n_693), .Y(n_430) );
NAND4xp25_ASAP7_75t_L g431 ( .A(n_432), .B(n_532), .C(n_559), .D(n_582), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_481), .B(n_491), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_447), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_SL g511 ( .A(n_435), .Y(n_511) );
AND2x4_ASAP7_75t_L g545 ( .A(n_435), .B(n_534), .Y(n_545) );
OR2x2_ASAP7_75t_L g555 ( .A(n_435), .B(n_513), .Y(n_555) );
OR2x2_ASAP7_75t_L g601 ( .A(n_435), .B(n_450), .Y(n_601) );
AND2x2_ASAP7_75t_L g615 ( .A(n_435), .B(n_512), .Y(n_615) );
AND2x2_ASAP7_75t_L g658 ( .A(n_435), .B(n_548), .Y(n_658) );
AND2x2_ASAP7_75t_L g665 ( .A(n_435), .B(n_524), .Y(n_665) );
AND2x2_ASAP7_75t_L g684 ( .A(n_435), .B(n_574), .Y(n_684) );
AND2x2_ASAP7_75t_L g702 ( .A(n_435), .B(n_544), .Y(n_702) );
OR2x6_ASAP7_75t_L g435 ( .A(n_436), .B(n_445), .Y(n_435) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_443), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g667 ( .A(n_447), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_462), .Y(n_447) );
AND2x2_ASAP7_75t_L g577 ( .A(n_448), .B(n_512), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_448), .B(n_597), .Y(n_596) );
AOI32xp33_ASAP7_75t_L g610 ( .A1(n_448), .A2(n_611), .A3(n_614), .B1(n_616), .B2(n_620), .Y(n_610) );
AND2x2_ASAP7_75t_L g680 ( .A(n_448), .B(n_574), .Y(n_680) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g544 ( .A(n_450), .B(n_513), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_450), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g586 ( .A(n_450), .B(n_533), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_450), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_452), .A2(n_460), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g551 ( .A(n_462), .B(n_495), .Y(n_551) );
AND2x2_ASAP7_75t_L g627 ( .A(n_462), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g699 ( .A(n_462), .Y(n_699) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .Y(n_462) );
OR2x2_ASAP7_75t_L g494 ( .A(n_463), .B(n_472), .Y(n_494) );
AND2x2_ASAP7_75t_L g508 ( .A(n_463), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_463), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g558 ( .A(n_463), .Y(n_558) );
AND2x2_ASAP7_75t_L g585 ( .A(n_463), .B(n_472), .Y(n_585) );
BUFx3_ASAP7_75t_L g588 ( .A(n_463), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_463), .B(n_563), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_463), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g539 ( .A(n_471), .Y(n_539) );
AND2x2_ASAP7_75t_L g557 ( .A(n_471), .B(n_537), .Y(n_557) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g568 ( .A(n_472), .B(n_483), .Y(n_568) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_472), .Y(n_581) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_480), .Y(n_472) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_473), .A2(n_484), .B(n_490), .Y(n_483) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_473), .A2(n_525), .B(n_531), .Y(n_524) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_482), .B(n_588), .Y(n_638) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_SL g509 ( .A(n_483), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_483), .B(n_557), .C(n_558), .Y(n_556) );
OR2x2_ASAP7_75t_L g564 ( .A(n_483), .B(n_537), .Y(n_564) );
AND2x2_ASAP7_75t_L g584 ( .A(n_483), .B(n_537), .Y(n_584) );
AND2x2_ASAP7_75t_L g628 ( .A(n_483), .B(n_497), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_507), .B(n_510), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g703 ( .A(n_493), .B(n_628), .Y(n_703) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_494), .A2(n_601), .B1(n_643), .B2(n_645), .Y(n_642) );
OR2x2_ASAP7_75t_L g649 ( .A(n_494), .B(n_564), .Y(n_649) );
OR2x2_ASAP7_75t_L g673 ( .A(n_494), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_494), .B(n_593), .Y(n_686) );
AND2x2_ASAP7_75t_L g579 ( .A(n_495), .B(n_580), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_495), .A2(n_652), .B(n_667), .Y(n_666) );
AOI32xp33_ASAP7_75t_L g687 ( .A1(n_495), .A2(n_577), .A3(n_688), .B1(n_690), .B2(n_691), .Y(n_687) );
OR2x2_ASAP7_75t_L g698 ( .A(n_495), .B(n_699), .Y(n_698) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g566 ( .A(n_496), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_496), .B(n_580), .Y(n_645) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g537 ( .A(n_497), .Y(n_537) );
AND2x2_ASAP7_75t_L g603 ( .A(n_497), .B(n_568), .Y(n_603) );
AND3x2_ASAP7_75t_L g612 ( .A(n_497), .B(n_508), .C(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g538 ( .A(n_509), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_509), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_509), .B(n_537), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_L g533 ( .A(n_511), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g573 ( .A(n_511), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g591 ( .A(n_511), .B(n_524), .Y(n_591) );
AND2x2_ASAP7_75t_L g609 ( .A(n_511), .B(n_513), .Y(n_609) );
OR2x2_ASAP7_75t_L g623 ( .A(n_511), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g669 ( .A(n_511), .B(n_597), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_512), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
AND2x2_ASAP7_75t_L g570 ( .A(n_513), .B(n_548), .Y(n_570) );
OR2x2_ASAP7_75t_L g624 ( .A(n_513), .B(n_548), .Y(n_624) );
AND2x2_ASAP7_75t_L g677 ( .A(n_513), .B(n_534), .Y(n_677) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g575 ( .A(n_514), .Y(n_575) );
AND2x2_ASAP7_75t_L g597 ( .A(n_514), .B(n_524), .Y(n_597) );
INVx2_ASAP7_75t_L g534 ( .A(n_524), .Y(n_534) );
INVx1_ASAP7_75t_L g554 ( .A(n_524), .Y(n_554) );
AOI211xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B(n_540), .C(n_552), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_533), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g696 ( .A(n_533), .Y(n_696) );
AND2x2_ASAP7_75t_L g574 ( .A(n_534), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_537), .B(n_538), .Y(n_546) );
INVx1_ASAP7_75t_L g631 ( .A(n_537), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_537), .B(n_558), .Y(n_655) );
AND2x2_ASAP7_75t_L g671 ( .A(n_537), .B(n_585), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_538), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g562 ( .A(n_539), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B1(n_547), .B2(n_550), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_543), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_544), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g569 ( .A(n_545), .B(n_570), .Y(n_569) );
AOI221xp5_ASAP7_75t_SL g634 ( .A1(n_545), .A2(n_587), .B1(n_635), .B2(n_640), .C(n_642), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_545), .B(n_608), .Y(n_641) );
INVx1_ASAP7_75t_L g701 ( .A(n_547), .Y(n_701) );
BUFx3_ASAP7_75t_L g608 ( .A(n_548), .Y(n_608) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI21xp33_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_555), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_554), .B(n_608), .Y(n_661) );
INVx1_ASAP7_75t_L g618 ( .A(n_555), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_555), .B(n_608), .Y(n_619) );
INVxp67_ASAP7_75t_L g639 ( .A(n_557), .Y(n_639) );
AND2x2_ASAP7_75t_L g580 ( .A(n_558), .B(n_581), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_565), .B(n_569), .C(n_571), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_SL g594 ( .A(n_562), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_563), .B(n_594), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_563), .B(n_585), .Y(n_636) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_566), .A2(n_572), .B1(n_576), .B2(n_578), .Y(n_571) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g587 ( .A(n_568), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g632 ( .A(n_568), .B(n_633), .Y(n_632) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_570), .A2(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_574), .A2(n_583), .B1(n_586), .B2(n_587), .C(n_589), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_574), .B(n_608), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_574), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g690 ( .A(n_580), .Y(n_690) );
INVxp67_ASAP7_75t_L g613 ( .A(n_581), .Y(n_613) );
INVx1_ASAP7_75t_L g620 ( .A(n_583), .Y(n_620) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g659 ( .A(n_584), .B(n_588), .Y(n_659) );
INVx1_ASAP7_75t_L g633 ( .A(n_588), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_588), .B(n_603), .Y(n_663) );
OAI32xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .A3(n_594), .B1(n_595), .B2(n_596), .Y(n_589) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g602 ( .A(n_597), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_597), .B(n_629), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_597), .B(n_658), .Y(n_689) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_597), .B(n_608), .Y(n_697) );
NAND5xp2_ASAP7_75t_L g598 ( .A(n_599), .B(n_621), .C(n_634), .D(n_646), .E(n_647), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_604), .B2(n_606), .C(n_610), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp33_ASAP7_75t_SL g625 ( .A(n_605), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_608), .B(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_609), .A2(n_622), .B1(n_625), .B2(n_629), .Y(n_621) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_612), .A2(n_617), .B(n_618), .C(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g644 ( .A(n_624), .Y(n_644) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_633), .B(n_682), .Y(n_692) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B1(n_652), .B2(n_656), .C1(n_659), .C2(n_660), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_666), .B2(n_668), .C(n_670), .Y(n_662) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_675), .Y(n_670) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g682 ( .A(n_674), .Y(n_682) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B1(n_683), .B2(n_685), .C(n_687), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .B(n_698), .C(n_700), .Y(n_693) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g710 ( .A(n_704), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_705), .Y(n_711) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_720), .Y(n_715) );
NOR2xp33_ASAP7_75t_SL g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_SL g738 ( .A(n_717), .Y(n_738) );
INVx1_ASAP7_75t_L g737 ( .A(n_719), .Y(n_737) );
OA21x2_ASAP7_75t_L g740 ( .A1(n_719), .A2(n_738), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g728 ( .A(n_720), .Y(n_728) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g732 ( .A(n_722), .Y(n_732) );
BUFx2_ASAP7_75t_L g741 ( .A(n_722), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g723 ( .A1(n_724), .A2(n_728), .B(n_729), .Y(n_723) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
CKINVDCx6p67_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
endmodule