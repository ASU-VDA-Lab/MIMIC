module real_aes_8665_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_0), .A2(n_168), .B(n_171), .C(n_175), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_1), .B(n_159), .Y(n_178) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_2), .B(n_86), .C(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g444 ( .A(n_2), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_3), .B(n_169), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_4), .A2(n_132), .B(n_135), .C(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_5), .A2(n_127), .B(n_542), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_6), .A2(n_127), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_7), .B(n_159), .Y(n_548) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_8), .A2(n_161), .B(n_233), .Y(n_232) );
AND2x6_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_10), .A2(n_132), .B(n_135), .C(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g508 ( .A(n_11), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_12), .B(n_39), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_13), .B(n_174), .Y(n_519) );
INVx1_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_15), .B(n_169), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_16), .A2(n_170), .B(n_528), .C(n_530), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_17), .B(n_159), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_18), .B(n_147), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_19), .A2(n_135), .B(n_138), .C(n_146), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_20), .A2(n_173), .B(n_241), .C(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_21), .B(n_174), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g449 ( .A1(n_22), .A2(n_74), .B1(n_450), .B2(n_739), .C1(n_742), .C2(n_743), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_23), .B(n_174), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_24), .Y(n_489) );
INVx1_ASAP7_75t_L g469 ( .A(n_25), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_26), .A2(n_135), .B(n_146), .C(n_236), .Y(n_235) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_28), .Y(n_515) );
INVx1_ASAP7_75t_L g483 ( .A(n_29), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_30), .A2(n_127), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g130 ( .A(n_31), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_32), .A2(n_185), .B(n_186), .C(n_190), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_33), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_34), .A2(n_173), .B(n_545), .C(n_547), .Y(n_544) );
INVxp67_ASAP7_75t_L g484 ( .A(n_35), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_36), .B(n_238), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_37), .A2(n_135), .B(n_146), .C(n_468), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g543 ( .A(n_38), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_40), .A2(n_175), .B(n_506), .C(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_41), .B(n_126), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_42), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_43), .B(n_169), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_44), .B(n_127), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_45), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_46), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_47), .B(n_446), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_48), .A2(n_185), .B(n_190), .C(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g172 ( .A(n_49), .Y(n_172) );
INVx1_ASAP7_75t_L g216 ( .A(n_50), .Y(n_216) );
INVx1_ASAP7_75t_L g556 ( .A(n_51), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_52), .B(n_127), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_53), .Y(n_155) );
CKINVDCx14_ASAP7_75t_R g504 ( .A(n_54), .Y(n_504) );
INVx1_ASAP7_75t_L g133 ( .A(n_55), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_56), .B(n_127), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_57), .B(n_159), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_58), .A2(n_145), .B(n_201), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g152 ( .A(n_59), .Y(n_152) );
INVx1_ASAP7_75t_SL g546 ( .A(n_60), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_61), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_62), .B(n_169), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_63), .B(n_159), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_64), .B(n_170), .Y(n_251) );
INVx1_ASAP7_75t_L g492 ( .A(n_65), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_66), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_67), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_68), .A2(n_135), .B(n_190), .C(n_199), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_69), .Y(n_225) );
INVx1_ASAP7_75t_L g107 ( .A(n_70), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_71), .A2(n_127), .B(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_72), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_73), .A2(n_127), .B(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_74), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_75), .A2(n_126), .B(n_479), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_76), .Y(n_466) );
INVx1_ASAP7_75t_L g526 ( .A(n_77), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_78), .B(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_79), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_80), .A2(n_127), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g529 ( .A(n_81), .Y(n_529) );
INVx2_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
INVx1_ASAP7_75t_L g518 ( .A(n_83), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_84), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_85), .B(n_174), .Y(n_252) );
OR2x2_ASAP7_75t_L g441 ( .A(n_86), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g453 ( .A(n_86), .B(n_443), .Y(n_453) );
INVx2_ASAP7_75t_L g458 ( .A(n_86), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_87), .A2(n_135), .B(n_190), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_88), .B(n_127), .Y(n_183) );
INVx1_ASAP7_75t_L g187 ( .A(n_89), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_90), .A2(n_100), .B1(n_108), .B2(n_747), .Y(n_99) );
INVxp67_ASAP7_75t_L g228 ( .A(n_91), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_92), .A2(n_115), .B1(n_437), .B2(n_438), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_92), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_93), .B(n_161), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_94), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g200 ( .A(n_95), .Y(n_200) );
INVx1_ASAP7_75t_L g247 ( .A(n_96), .Y(n_247) );
INVx2_ASAP7_75t_L g559 ( .A(n_97), .Y(n_559) );
AND2x2_ASAP7_75t_L g218 ( .A(n_98), .B(n_149), .Y(n_218) );
BUFx4f_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
CKINVDCx6p67_ASAP7_75t_R g747 ( .A(n_101), .Y(n_747) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
AND2x2_ASAP7_75t_L g443 ( .A(n_102), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AO21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_113), .B(n_448), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g746 ( .A(n_110), .Y(n_746) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI21xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_439), .B(n_445), .Y(n_113) );
INVx1_ASAP7_75t_L g438 ( .A(n_115), .Y(n_438) );
INVx2_ASAP7_75t_L g454 ( .A(n_115), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_115), .A2(n_451), .B1(n_740), .B2(n_741), .Y(n_739) );
AND2x2_ASAP7_75t_SL g115 ( .A(n_116), .B(n_392), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_327), .Y(n_116) );
NAND4xp25_ASAP7_75t_SL g117 ( .A(n_118), .B(n_272), .C(n_296), .D(n_319), .Y(n_117) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_209), .B1(n_243), .B2(n_256), .C(n_259), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_179), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_121), .A2(n_157), .B1(n_210), .B2(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_121), .B(n_180), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_121), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_121), .B(n_333), .Y(n_419) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_157), .Y(n_121) );
AND2x2_ASAP7_75t_L g287 ( .A(n_122), .B(n_180), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_122), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_122), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_122), .B(n_158), .Y(n_315) );
INVx2_ASAP7_75t_L g347 ( .A(n_122), .Y(n_347) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_122), .Y(n_391) );
AND2x2_ASAP7_75t_L g408 ( .A(n_122), .B(n_285), .Y(n_408) );
INVx5_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g326 ( .A(n_123), .B(n_285), .Y(n_326) );
AND2x4_ASAP7_75t_L g340 ( .A(n_123), .B(n_157), .Y(n_340) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_123), .Y(n_344) );
AND2x2_ASAP7_75t_L g364 ( .A(n_123), .B(n_279), .Y(n_364) );
AND2x2_ASAP7_75t_L g414 ( .A(n_123), .B(n_181), .Y(n_414) );
AND2x2_ASAP7_75t_L g424 ( .A(n_123), .B(n_158), .Y(n_424) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_154), .Y(n_123) );
AOI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_134), .B(n_147), .Y(n_124) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g248 ( .A(n_128), .B(n_132), .Y(n_248) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g242 ( .A(n_130), .Y(n_242) );
INVx1_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_131), .Y(n_141) );
INVx3_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
INVx1_ASAP7_75t_L g238 ( .A(n_131), .Y(n_238) );
BUFx3_ASAP7_75t_L g146 ( .A(n_132), .Y(n_146) );
INVx4_ASAP7_75t_SL g177 ( .A(n_132), .Y(n_177) );
INVx5_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx3_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_136), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_142), .B(n_144), .Y(n_138) );
INVx2_ASAP7_75t_L g143 ( .A(n_140), .Y(n_143) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_143), .A2(n_187), .B(n_188), .C(n_189), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_143), .A2(n_189), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_143), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g517 ( .A1(n_143), .A2(n_494), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_144), .A2(n_169), .B(n_469), .C(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_145), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_148), .B(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_149), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_149), .A2(n_213), .B(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_149), .A2(n_248), .B(n_466), .C(n_467), .Y(n_465) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_149), .A2(n_502), .B(n_509), .Y(n_501) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_L g162 ( .A(n_150), .B(n_151), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_156), .A2(n_514), .B(n_520), .Y(n_513) );
AND2x2_ASAP7_75t_L g280 ( .A(n_157), .B(n_180), .Y(n_280) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_157), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_157), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g370 ( .A(n_157), .Y(n_370) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g258 ( .A(n_158), .B(n_195), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_158), .B(n_196), .Y(n_285) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_163), .B(n_178), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_160), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_160), .A2(n_197), .B(n_207), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_160), .B(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_160), .A2(n_246), .B(n_253), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_160), .B(n_472), .Y(n_471) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_160), .A2(n_488), .B(n_495), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_160), .B(n_521), .Y(n_520) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_161), .A2(n_234), .B(n_235), .Y(n_233) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g255 ( .A(n_162), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_177), .Y(n_164) );
INVx2_ASAP7_75t_L g185 ( .A(n_166), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_166), .A2(n_177), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_166), .A2(n_177), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_166), .A2(n_177), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_166), .A2(n_177), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_166), .A2(n_177), .B(n_543), .C(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_166), .A2(n_177), .B(n_556), .C(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_169), .B(n_228), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_169), .A2(n_202), .B1(n_483), .B2(n_484), .Y(n_482) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_170), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_173), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g506 ( .A(n_174), .Y(n_506) );
INVx2_ASAP7_75t_L g494 ( .A(n_175), .Y(n_494) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_176), .Y(n_189) );
INVx1_ASAP7_75t_L g530 ( .A(n_176), .Y(n_530) );
INVx1_ASAP7_75t_L g190 ( .A(n_177), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_179), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_193), .Y(n_179) );
OR2x2_ASAP7_75t_L g311 ( .A(n_180), .B(n_194), .Y(n_311) );
AND2x2_ASAP7_75t_L g348 ( .A(n_180), .B(n_258), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_180), .B(n_279), .Y(n_359) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_180), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_180), .B(n_315), .Y(n_432) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx2_ASAP7_75t_L g257 ( .A(n_181), .Y(n_257) );
AND2x2_ASAP7_75t_L g266 ( .A(n_181), .B(n_194), .Y(n_266) );
AND2x2_ASAP7_75t_L g382 ( .A(n_181), .B(n_277), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_181), .B(n_315), .Y(n_404) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_194), .Y(n_350) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_195), .Y(n_302) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g279 ( .A(n_196), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_206), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_203), .C(n_204), .Y(n_199) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_202), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_202), .B(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g547 ( .A(n_205), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_219), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_210), .B(n_292), .Y(n_411) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_211), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g263 ( .A(n_211), .B(n_264), .Y(n_263) );
INVx5_ASAP7_75t_SL g271 ( .A(n_211), .Y(n_271) );
OR2x2_ASAP7_75t_L g294 ( .A(n_211), .B(n_264), .Y(n_294) );
OR2x2_ASAP7_75t_L g304 ( .A(n_211), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g367 ( .A(n_211), .B(n_221), .Y(n_367) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_211), .B(n_220), .Y(n_405) );
NOR4xp25_ASAP7_75t_L g426 ( .A(n_211), .B(n_347), .C(n_427), .D(n_428), .Y(n_426) );
AND2x2_ASAP7_75t_L g436 ( .A(n_211), .B(n_268), .Y(n_436) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_218), .Y(n_211) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g261 ( .A(n_220), .B(n_257), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_220), .B(n_263), .Y(n_430) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
OR2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_221), .B(n_245), .Y(n_289) );
INVxp67_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_221), .B(n_264), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_221), .B(n_231), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_221), .B(n_268), .Y(n_373) );
OR2x2_ASAP7_75t_L g402 ( .A(n_221), .B(n_231), .Y(n_402) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_221) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_222), .A2(n_524), .B(n_531), .Y(n_523) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_222), .A2(n_541), .B(n_548), .Y(n_540) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_222), .A2(n_554), .B(n_560), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_230), .B(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_230), .B(n_271), .Y(n_410) );
OR2x2_ASAP7_75t_L g431 ( .A(n_230), .B(n_308), .Y(n_431) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g244 ( .A(n_231), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g268 ( .A(n_231), .B(n_264), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_231), .B(n_245), .Y(n_283) );
AND2x2_ASAP7_75t_L g353 ( .A(n_231), .B(n_277), .Y(n_353) );
AND2x2_ASAP7_75t_L g387 ( .A(n_231), .B(n_271), .Y(n_387) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_232), .B(n_271), .Y(n_290) );
AND2x2_ASAP7_75t_L g318 ( .A(n_232), .B(n_245), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_240), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_240), .A2(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_243), .B(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_244), .A2(n_333), .B1(n_369), .B2(n_386), .C(n_388), .Y(n_385) );
INVx5_ASAP7_75t_SL g264 ( .A(n_245), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_249), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_248), .A2(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_248), .A2(n_515), .B(n_516), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g477 ( .A(n_255), .Y(n_477) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI33xp33_ASAP7_75t_L g284 ( .A1(n_257), .A2(n_285), .A3(n_286), .B1(n_288), .B2(n_291), .B3(n_295), .Y(n_284) );
OR2x2_ASAP7_75t_L g300 ( .A(n_257), .B(n_301), .Y(n_300) );
AOI322xp5_ASAP7_75t_L g409 ( .A1(n_257), .A2(n_326), .A3(n_333), .B1(n_410), .B2(n_411), .C1(n_412), .C2(n_415), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_257), .B(n_285), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_SL g433 ( .A1(n_257), .A2(n_285), .B(n_434), .C(n_436), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_258), .A2(n_273), .B1(n_278), .B2(n_281), .C(n_284), .Y(n_272) );
INVx1_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_258), .B(n_414), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B1(n_265), .B2(n_267), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g342 ( .A(n_263), .B(n_277), .Y(n_342) );
AND2x2_ASAP7_75t_L g400 ( .A(n_263), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g308 ( .A(n_264), .B(n_271), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_264), .B(n_277), .Y(n_336) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_266), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_266), .B(n_344), .Y(n_398) );
OAI321xp33_ASAP7_75t_L g417 ( .A1(n_266), .A2(n_339), .A3(n_418), .B1(n_419), .B2(n_420), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g384 ( .A(n_267), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_268), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g323 ( .A(n_268), .B(n_271), .Y(n_323) );
AOI321xp33_ASAP7_75t_L g381 ( .A1(n_268), .A2(n_285), .A3(n_382), .B1(n_383), .B2(n_384), .C(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g298 ( .A(n_270), .B(n_283), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_271), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_271), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_271), .B(n_357), .Y(n_394) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g317 ( .A(n_275), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g282 ( .A(n_276), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g390 ( .A(n_277), .Y(n_390) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_280), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_287), .B(n_322), .Y(n_371) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OR2x2_ASAP7_75t_L g335 ( .A(n_290), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g380 ( .A(n_290), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_291), .A2(n_338), .B1(n_341), .B2(n_343), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g435 ( .A(n_294), .B(n_358), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .B1(n_303), .B2(n_309), .C(n_312), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g379 ( .A(n_305), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_307), .B(n_357), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_307), .A2(n_375), .B(n_377), .Y(n_374) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g420 ( .A(n_308), .B(n_402), .Y(n_420) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_SL g322 ( .A(n_311), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g366 ( .A(n_318), .B(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g428 ( .A(n_318), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_322), .B(n_340), .Y(n_376) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
NAND5xp2_ASAP7_75t_L g327 ( .A(n_328), .B(n_345), .C(n_354), .D(n_374), .E(n_381), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B(n_334), .C(n_337), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_341), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_349), .B(n_351), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_346), .A2(n_400), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_399) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AOI321xp33_ASAP7_75t_L g354 ( .A1(n_347), .A2(n_355), .A3(n_359), .B1(n_360), .B2(n_366), .C(n_368), .Y(n_354) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g425 ( .A(n_359), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g377 ( .A(n_362), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NOR2xp67_ASAP7_75t_SL g389 ( .A(n_363), .B(n_370), .Y(n_389) );
AOI321xp33_ASAP7_75t_SL g421 ( .A1(n_366), .A2(n_422), .A3(n_423), .B1(n_424), .B2(n_425), .C(n_426), .Y(n_421) );
O2A1O1Ixp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_371), .C(n_372), .Y(n_368) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_379), .B(n_387), .Y(n_416) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .C(n_391), .Y(n_388) );
NOR3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_417), .C(n_429), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_395), .B(n_399), .C(n_409), .Y(n_393) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_398), .A2(n_430), .B1(n_431), .B2(n_432), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g422 ( .A(n_420), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
CKINVDCx14_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_441), .Y(n_447) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_442), .B(n_458), .Y(n_745) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g457 ( .A(n_443), .B(n_458), .Y(n_457) );
AOI21xp33_ASAP7_75t_L g448 ( .A1(n_445), .A2(n_449), .B(n_746), .Y(n_448) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B1(n_455), .B2(n_459), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g741 ( .A(n_456), .Y(n_741) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g740 ( .A(n_459), .Y(n_740) );
OR4x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_629), .C(n_676), .D(n_716), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_575), .C(n_604), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_497), .B(n_532), .C(n_568), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_462), .A2(n_588), .B(n_605), .C(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_473), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_464), .B(n_567), .Y(n_566) );
INVx3_ASAP7_75t_SL g571 ( .A(n_464), .Y(n_571) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_464), .Y(n_583) );
AND2x4_ASAP7_75t_L g587 ( .A(n_464), .B(n_539), .Y(n_587) );
AND2x2_ASAP7_75t_L g598 ( .A(n_464), .B(n_487), .Y(n_598) );
OR2x2_ASAP7_75t_L g622 ( .A(n_464), .B(n_535), .Y(n_622) );
AND2x2_ASAP7_75t_L g635 ( .A(n_464), .B(n_540), .Y(n_635) );
AND2x2_ASAP7_75t_L g675 ( .A(n_464), .B(n_661), .Y(n_675) );
AND2x2_ASAP7_75t_L g682 ( .A(n_464), .B(n_645), .Y(n_682) );
AND2x2_ASAP7_75t_L g712 ( .A(n_464), .B(n_474), .Y(n_712) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_471), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_473), .B(n_639), .Y(n_651) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_474), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g589 ( .A(n_474), .B(n_486), .Y(n_589) );
BUFx3_ASAP7_75t_L g597 ( .A(n_474), .Y(n_597) );
OR2x2_ASAP7_75t_L g618 ( .A(n_474), .B(n_500), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_474), .B(n_639), .Y(n_729) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_478), .B(n_485), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_476), .A2(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g536 ( .A(n_478), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_485), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_486), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
AND2x2_ASAP7_75t_L g645 ( .A(n_486), .B(n_540), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_486), .A2(n_648), .B1(n_650), .B2(n_652), .C(n_653), .Y(n_647) );
AND2x2_ASAP7_75t_L g661 ( .A(n_486), .B(n_535), .Y(n_661) );
AND2x2_ASAP7_75t_L g687 ( .A(n_486), .B(n_571), .Y(n_687) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g567 ( .A(n_487), .B(n_540), .Y(n_567) );
BUFx2_ASAP7_75t_L g701 ( .A(n_487), .Y(n_701) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI32xp33_ASAP7_75t_L g667 ( .A1(n_498), .A2(n_628), .A3(n_642), .B1(n_668), .B2(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
AND2x2_ASAP7_75t_L g608 ( .A(n_499), .B(n_552), .Y(n_608) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g590 ( .A(n_500), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_500), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g662 ( .A(n_500), .B(n_552), .Y(n_662) );
AND2x2_ASAP7_75t_L g673 ( .A(n_500), .B(n_565), .Y(n_673) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g574 ( .A(n_501), .B(n_553), .Y(n_574) );
AND2x2_ASAP7_75t_L g578 ( .A(n_501), .B(n_553), .Y(n_578) );
AND2x2_ASAP7_75t_L g613 ( .A(n_501), .B(n_564), .Y(n_613) );
AND2x2_ASAP7_75t_L g620 ( .A(n_501), .B(n_522), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_501), .A2(n_571), .B(n_582), .C(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g679 ( .A(n_501), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_501), .B(n_512), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_510), .B(n_562), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_510), .B(n_578), .Y(n_668) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g573 ( .A(n_511), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
AND2x2_ASAP7_75t_L g565 ( .A(n_512), .B(n_523), .Y(n_565) );
OR2x2_ASAP7_75t_L g580 ( .A(n_512), .B(n_523), .Y(n_580) );
AND2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_564), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_512), .Y(n_607) );
AND2x2_ASAP7_75t_L g626 ( .A(n_512), .B(n_563), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_512), .A2(n_591), .B1(n_637), .B2(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_512), .B(n_679), .Y(n_703) );
AND2x2_ASAP7_75t_L g718 ( .A(n_512), .B(n_578), .Y(n_718) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g550 ( .A(n_513), .Y(n_550) );
AND2x2_ASAP7_75t_L g592 ( .A(n_513), .B(n_523), .Y(n_592) );
AND2x2_ASAP7_75t_L g594 ( .A(n_513), .B(n_552), .Y(n_594) );
AND3x2_ASAP7_75t_L g656 ( .A(n_513), .B(n_620), .C(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g691 ( .A(n_522), .B(n_563), .Y(n_691) );
INVx1_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g552 ( .A(n_523), .B(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_523), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_523), .B(n_562), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_523), .B(n_603), .C(n_679), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_549), .B1(n_561), .B2(n_566), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_535), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g643 ( .A(n_535), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g659 ( .A1(n_538), .A2(n_660), .A3(n_661), .B(n_662), .Y(n_659) );
AND2x2_ASAP7_75t_L g684 ( .A(n_538), .B(n_571), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_538), .B(n_597), .Y(n_730) );
AND2x2_ASAP7_75t_L g639 ( .A(n_539), .B(n_571), .Y(n_639) );
AND2x2_ASAP7_75t_L g700 ( .A(n_539), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g570 ( .A(n_540), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g628 ( .A(n_540), .Y(n_628) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
CKINVDCx16_ASAP7_75t_R g649 ( .A(n_550), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_551), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AOI221x1_ASAP7_75t_SL g616 ( .A1(n_552), .A2(n_617), .B1(n_619), .B2(n_621), .C(n_623), .Y(n_616) );
INVx2_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_553), .Y(n_658) );
INVx1_ASAP7_75t_L g646 ( .A(n_561), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_562), .B(n_579), .Y(n_671) );
INVx1_ASAP7_75t_SL g734 ( .A(n_562), .Y(n_734) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g652 ( .A(n_565), .B(n_578), .Y(n_652) );
INVx1_ASAP7_75t_L g720 ( .A(n_566), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_566), .B(n_649), .Y(n_733) );
INVx2_ASAP7_75t_SL g572 ( .A(n_567), .Y(n_572) );
AND2x2_ASAP7_75t_L g615 ( .A(n_567), .B(n_571), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_567), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_567), .B(n_642), .Y(n_669) );
AOI21xp33_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_572), .B(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_570), .B(n_642), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_570), .B(n_597), .Y(n_738) );
OR2x2_ASAP7_75t_L g610 ( .A(n_571), .B(n_589), .Y(n_610) );
AND2x2_ASAP7_75t_L g709 ( .A(n_571), .B(n_700), .Y(n_709) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_572), .A2(n_585), .B1(n_590), .B2(n_593), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_572), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g632 ( .A(n_574), .B(n_580), .Y(n_632) );
INVx1_ASAP7_75t_L g696 ( .A(n_574), .Y(n_696) );
AOI311xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_581), .A3(n_583), .B(n_584), .C(n_595), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_579), .A2(n_711), .B1(n_723), .B2(n_726), .C(n_728), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_579), .B(n_734), .Y(n_736) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g633 ( .A(n_581), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_582), .A2(n_624), .B(n_625), .C(n_627), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
O2A1O1Ixp33_ASAP7_75t_SL g692 ( .A1(n_586), .A2(n_588), .B(n_693), .C(n_694), .Y(n_692) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_587), .B(n_661), .Y(n_727) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_590), .A2(n_610), .B1(n_611), .B2(n_614), .C(n_616), .Y(n_609) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g612 ( .A(n_592), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g695 ( .A(n_592), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_596), .A2(n_654), .B(n_655), .C(n_659), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_597), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_597), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g619 ( .A(n_603), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_607), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g721 ( .A(n_610), .Y(n_721) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_613), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g648 ( .A(n_613), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g725 ( .A(n_613), .Y(n_725) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g666 ( .A(n_615), .B(n_642), .Y(n_666) );
INVx1_ASAP7_75t_SL g660 ( .A(n_622), .Y(n_660) );
INVx1_ASAP7_75t_L g637 ( .A(n_628), .Y(n_637) );
NAND3xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_647), .C(n_663), .Y(n_629) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .A3(n_634), .B1(n_636), .B2(n_640), .C1(n_644), .C2(n_646), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g683 ( .A1(n_631), .A2(n_684), .B(n_685), .C(n_692), .Y(n_683) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_634), .A2(n_655), .B1(n_686), .B2(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g644 ( .A(n_642), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g681 ( .A(n_642), .B(n_682), .Y(n_681) );
AOI32xp33_ASAP7_75t_L g732 ( .A1(n_642), .A2(n_733), .A3(n_734), .B1(n_735), .B2(n_737), .Y(n_732) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g654 ( .A(n_645), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_645), .A2(n_698), .B1(n_702), .B2(n_704), .C(n_707), .Y(n_697) );
AND2x2_ASAP7_75t_L g711 ( .A(n_645), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g714 ( .A(n_649), .B(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g724 ( .A(n_649), .B(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g715 ( .A(n_658), .B(n_679), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_667), .C(n_670), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_674), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_680), .B(n_683), .C(n_697), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_691), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g706 ( .A(n_703), .Y(n_706) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_713), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI211xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_719), .B(n_722), .C(n_732), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI21xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
endmodule