module fake_jpeg_2300_n_543 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_543);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_72),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_9),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_27),
.B(n_7),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_81),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_7),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_91),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_93),
.Y(n_115)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_6),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_27),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_38),
.Y(n_99)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_15),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_105),
.B(n_131),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_50),
.B1(n_26),
.B2(n_30),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_107),
.A2(n_46),
.B1(n_84),
.B2(n_88),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_116),
.B(n_104),
.Y(n_211)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_73),
.B(n_94),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_56),
.Y(n_187)
);

BUFx4f_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_63),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_145),
.Y(n_170)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_142),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_68),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_67),
.B(n_50),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_158),
.Y(n_168)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_149),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_71),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_151),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_78),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_55),
.B(n_26),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_87),
.B(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_74),
.B(n_23),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_46),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_15),
.Y(n_223)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_167),
.Y(n_266)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_58),
.B1(n_40),
.B2(n_75),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_172),
.A2(n_193),
.B1(n_0),
.B2(n_2),
.Y(n_268)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_174),
.Y(n_256)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_176),
.B(n_189),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_178),
.Y(n_235)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_179),
.Y(n_253)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_183),
.Y(n_271)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_187),
.B(n_209),
.Y(n_234)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_126),
.B(n_46),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_116),
.A2(n_82),
.B1(n_79),
.B2(n_85),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_190),
.A2(n_197),
.B1(n_141),
.B2(n_128),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_127),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_204),
.B1(n_112),
.B2(n_164),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_135),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_40),
.B1(n_46),
.B2(n_30),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_135),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_198),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_140),
.B(n_102),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_111),
.A2(n_21),
.B(n_29),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_200),
.A2(n_17),
.B(n_18),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_29),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_202),
.B(n_205),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_113),
.A2(n_21),
.B(n_69),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_139),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_56),
.B1(n_51),
.B2(n_42),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_108),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_132),
.B(n_16),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_223),
.Y(n_265)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_16),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_215),
.Y(n_269)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_217),
.Y(n_240)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_222),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_221),
.Y(n_275)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_121),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_224),
.Y(n_251)
);

INVx6_ASAP7_75t_SL g225 ( 
.A(n_157),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_225),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_108),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_133),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_229),
.B(n_246),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_187),
.A2(n_160),
.B1(n_106),
.B2(n_110),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_230),
.A2(n_273),
.B1(n_182),
.B2(n_220),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_233),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_155),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_242),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_170),
.B(n_155),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_168),
.A2(n_153),
.B1(n_133),
.B2(n_125),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_247),
.B(n_254),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_191),
.A2(n_153),
.B1(n_125),
.B2(n_128),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_249),
.A2(n_255),
.B1(n_257),
.B2(n_260),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_200),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_274),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_141),
.B1(n_109),
.B2(n_51),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_217),
.A2(n_109),
.B1(n_42),
.B2(n_19),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_209),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_277),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_193),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_210),
.B(n_0),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_177),
.B(n_0),
.C(n_3),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

CKINVDCx10_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_280),
.Y(n_330)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_313),
.Y(n_362)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_245),
.B(n_173),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_291),
.B(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_171),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_298),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_265),
.B(n_236),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_304),
.B(n_307),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_171),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_278),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_300),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_242),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_306),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_229),
.A2(n_172),
.B1(n_212),
.B2(n_185),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_303),
.A2(n_282),
.B1(n_325),
.B2(n_314),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_220),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_186),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_265),
.B(n_216),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_252),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_240),
.A2(n_219),
.B1(n_195),
.B2(n_208),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_309),
.A2(n_319),
.B1(n_183),
.B2(n_271),
.Y(n_363)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_310),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_266),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_311),
.Y(n_366)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_316),
.Y(n_345)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_277),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_321),
.Y(n_349)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_228),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_323),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_230),
.B(n_169),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_326),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_266),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_250),
.C(n_243),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_331),
.B(n_332),
.C(n_353),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_234),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_335),
.B1(n_312),
.B2(n_283),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_290),
.A2(n_255),
.B1(n_247),
.B2(n_260),
.Y(n_335)
);

AOI32xp33_ASAP7_75t_L g337 ( 
.A1(n_302),
.A2(n_243),
.A3(n_250),
.B1(n_264),
.B2(n_237),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_290),
.A2(n_264),
.B(n_237),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_288),
.B(n_323),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_268),
.B1(n_227),
.B2(n_259),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_344),
.B1(n_352),
.B2(n_326),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_279),
.A2(n_253),
.B(n_238),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_343),
.A2(n_367),
.B(n_188),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_276),
.B1(n_259),
.B2(n_258),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_280),
.A2(n_271),
.B(n_253),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_361),
.B(n_285),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_314),
.A2(n_276),
.B1(n_258),
.B2(n_201),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_231),
.C(n_216),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_305),
.B(n_182),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_368),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_282),
.A2(n_296),
.B(n_303),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_296),
.A2(n_231),
.B(n_167),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_224),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_355),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_378),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_362),
.A2(n_281),
.B(n_294),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_370),
.B(n_382),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_284),
.Y(n_372)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_324),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_373),
.B(n_381),
.Y(n_411)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_377),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_355),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_287),
.Y(n_379)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_334),
.A2(n_286),
.B1(n_315),
.B2(n_321),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_380),
.A2(n_388),
.B1(n_374),
.B2(n_378),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_316),
.Y(n_381)
);

INVx13_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_385),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_319),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_387),
.A2(n_351),
.B1(n_350),
.B2(n_333),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_361),
.A2(n_328),
.B1(n_340),
.B2(n_362),
.Y(n_388)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_390),
.Y(n_420)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_289),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_391),
.A2(n_400),
.B1(n_364),
.B2(n_358),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_292),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_392),
.B(n_345),
.Y(n_424)
);

INVx6_ASAP7_75t_SL g393 ( 
.A(n_362),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_394),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_328),
.B(n_318),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_367),
.A2(n_310),
.B(n_313),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_404),
.B(n_342),
.Y(n_425)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_399),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_317),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_403),
.C(n_206),
.Y(n_428)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_301),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_354),
.A2(n_352),
.B1(n_349),
.B2(n_344),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_401),
.A2(n_390),
.B1(n_384),
.B2(n_388),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_224),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_387),
.A2(n_343),
.B1(n_335),
.B2(n_333),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_405),
.A2(n_414),
.B1(n_429),
.B2(n_396),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_353),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_406),
.B(n_413),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_386),
.B(n_360),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_408),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_368),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_357),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_370),
.B(n_357),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_417),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_331),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_419),
.B(n_397),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_422),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_345),
.B(n_356),
.C(n_342),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_431),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_425),
.A2(n_389),
.B(n_385),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_402),
.C(n_386),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_369),
.A2(n_218),
.B1(n_3),
.B2(n_5),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_371),
.A2(n_3),
.B(n_5),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_432),
.A2(n_434),
.B1(n_375),
.B2(n_399),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_401),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_436),
.B(n_441),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_394),
.Y(n_440)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_391),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_443),
.B(n_446),
.C(n_447),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_445),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_398),
.C(n_403),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_380),
.C(n_404),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_449),
.A2(n_454),
.B1(n_425),
.B2(n_405),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_395),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_375),
.C(n_389),
.Y(n_452)
);

XNOR2x1_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_431),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_434),
.A2(n_376),
.B1(n_382),
.B2(n_377),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_412),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_460),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_376),
.Y(n_457)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_377),
.C(n_382),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_422),
.Y(n_461)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_461),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_416),
.B(n_432),
.C(n_420),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_416),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_435),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_470),
.Y(n_498)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_449),
.A2(n_415),
.B1(n_433),
.B2(n_430),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_474),
.A2(n_476),
.B1(n_439),
.B2(n_473),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_456),
.A2(n_415),
.B1(n_433),
.B2(n_430),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_482),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_442),
.B(n_426),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_480),
.B(n_484),
.Y(n_499)
);

XOR2x1_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_422),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_422),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_440),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_485),
.A2(n_490),
.B1(n_492),
.B2(n_495),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_486),
.A2(n_467),
.B1(n_468),
.B2(n_472),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_443),
.C(n_470),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_489),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_452),
.C(n_447),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_453),
.B(n_439),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_494),
.Y(n_513)
);

INVx13_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_482),
.B(n_462),
.CI(n_438),
.CON(n_493),
.SN(n_493)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_497),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_477),
.Y(n_494)
);

INVx13_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_464),
.Y(n_497)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_500),
.A2(n_418),
.B1(n_459),
.B2(n_454),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_474),
.A2(n_451),
.B(n_457),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_501),
.B(n_483),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_455),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_507),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_463),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_514),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_505),
.A2(n_509),
.B1(n_500),
.B2(n_497),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_465),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_489),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_499),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_458),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_484),
.C(n_480),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_510),
.A2(n_478),
.B(n_487),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_SL g516 ( 
.A(n_511),
.B(n_501),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_518),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_490),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_519),
.B(n_521),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_524),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_486),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_513),
.A2(n_448),
.B1(n_437),
.B2(n_445),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_460),
.C(n_487),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_512),
.C(n_514),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_529),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_517),
.A2(n_512),
.B(n_510),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_528),
.A2(n_504),
.B(n_493),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_525),
.B1(n_444),
.B2(n_523),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_532),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_516),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_533),
.A2(n_535),
.B(n_527),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_526),
.B(n_527),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_534),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_539),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_540),
.A2(n_536),
.B1(n_495),
.B2(n_437),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_523),
.B(n_493),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_542),
.A2(n_492),
.B(n_429),
.Y(n_543)
);


endmodule