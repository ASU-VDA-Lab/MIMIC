module fake_aes_5551_n_806 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_806);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_806;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_396;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_8), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_91), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_10), .Y(n_230) );
BUFx10_ASAP7_75t_L g231 ( .A(n_167), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_203), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_122), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_31), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_49), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_190), .B(n_102), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
CKINVDCx14_ASAP7_75t_R g238 ( .A(n_157), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_64), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_106), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_216), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_19), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_73), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_40), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_117), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_159), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_89), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_210), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_134), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_208), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_198), .B(n_109), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_20), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_82), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_87), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_155), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
BUFx5_ASAP7_75t_L g258 ( .A(n_196), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g259 ( .A(n_16), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_211), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_62), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_128), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_71), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_179), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_219), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_24), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_207), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_171), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_103), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_197), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_202), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_214), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_191), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_72), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_215), .Y(n_275) );
CKINVDCx14_ASAP7_75t_R g276 ( .A(n_172), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_114), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_124), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_186), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_131), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_153), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_116), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_100), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_65), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_36), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_93), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_218), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_95), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_213), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_199), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_204), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_59), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_101), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_32), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_193), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_121), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_94), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_205), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_180), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_209), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_57), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_147), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_139), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_75), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_108), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_92), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_34), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_145), .Y(n_308) );
BUFx5_ASAP7_75t_L g309 ( .A(n_201), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_126), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_137), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_136), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_10), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_169), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_52), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_206), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_135), .Y(n_317) );
BUFx10_ASAP7_75t_L g318 ( .A(n_18), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_88), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_144), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_99), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_38), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_110), .Y(n_323) );
BUFx2_ASAP7_75t_SL g324 ( .A(n_195), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_181), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_189), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_113), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_220), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_200), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_188), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_192), .Y(n_331) );
XNOR2xp5_ASAP7_75t_L g332 ( .A(n_77), .B(n_212), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_26), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_83), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_178), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_14), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_96), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_187), .Y(n_338) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_129), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_168), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_7), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_184), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_265), .B(n_0), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_228), .B(n_0), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_237), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_231), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_230), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_258), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_227), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_237), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_286), .B(n_1), .Y(n_351) );
BUFx8_ASAP7_75t_L g352 ( .A(n_258), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_258), .Y(n_354) );
OA21x2_ASAP7_75t_L g355 ( .A1(n_229), .A2(n_12), .B(n_11), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_234), .Y(n_356) );
BUFx8_ASAP7_75t_L g357 ( .A(n_258), .Y(n_357) );
BUFx8_ASAP7_75t_SL g358 ( .A(n_313), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_243), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_237), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_288), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_344), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_359), .B(n_339), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_348), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_351), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_354), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_351), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_344), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_345), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_349), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_349), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_356), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_353), .B(n_232), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_356), .Y(n_376) );
NOR2x1p5_ASAP7_75t_L g377 ( .A(n_346), .B(n_250), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_343), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_247), .B(n_245), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_372), .B(n_352), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_373), .B(n_357), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_376), .B(n_238), .Y(n_382) );
OR2x6_ASAP7_75t_L g383 ( .A(n_375), .B(n_361), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_371), .B(n_259), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_377), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_365), .A2(n_276), .B1(n_324), .B2(n_255), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_371), .B(n_233), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_364), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_375), .B(n_235), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_367), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_367), .B(n_239), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_362), .B(n_240), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_368), .B(n_241), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_378), .B(n_246), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_374), .B(n_248), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_366), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_379), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_369), .B(n_256), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_370), .B(n_261), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_363), .B(n_263), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_384), .A2(n_355), .B(n_257), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_382), .A2(n_355), .B(n_260), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_385), .B(n_332), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_398), .A2(n_262), .B(n_254), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_391), .A2(n_267), .B(n_268), .C(n_264), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_383), .B(n_341), .Y(n_407) );
BUFx4f_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_271), .B(n_275), .C(n_274), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_387), .A2(n_285), .B(n_277), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g411 ( .A(n_389), .B(n_251), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_392), .A2(n_291), .B(n_290), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_380), .A2(n_270), .B(n_249), .Y(n_413) );
AO21x1_ASAP7_75t_L g414 ( .A1(n_397), .A2(n_297), .B(n_294), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_381), .A2(n_300), .B(n_301), .C(n_298), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_401), .A2(n_303), .B(n_306), .C(n_302), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_316), .B(n_308), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_394), .A2(n_320), .B(n_327), .C(n_319), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_388), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_386), .B(n_273), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
BUFx4f_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_400), .A2(n_299), .B1(n_305), .B2(n_293), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_399), .Y(n_425) );
AO22x2_ASAP7_75t_L g426 ( .A1(n_407), .A2(n_358), .B1(n_329), .B2(n_334), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_411), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_424), .Y(n_428) );
AO32x2_ASAP7_75t_L g429 ( .A1(n_414), .A2(n_309), .A3(n_258), .B1(n_360), .B2(n_350), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_418), .A2(n_335), .B(n_336), .C(n_328), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_408), .B(n_317), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_409), .B(n_323), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_415), .B(n_242), .C(n_236), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_416), .B(n_266), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_419), .Y(n_435) );
OAI21x1_ASAP7_75t_SL g436 ( .A1(n_405), .A2(n_253), .B(n_244), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_413), .B(n_2), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_421), .B(n_3), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_419), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_404), .B(n_4), .Y(n_440) );
OAI21x1_ASAP7_75t_L g441 ( .A1(n_402), .A2(n_281), .B(n_278), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_403), .A2(n_410), .B(n_417), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_420), .B(n_5), .Y(n_443) );
AO31x2_ASAP7_75t_L g444 ( .A1(n_406), .A2(n_311), .A3(n_325), .B(n_307), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_422), .B(n_269), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_412), .A2(n_252), .B(n_292), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_425), .Y(n_447) );
OAI21x1_ASAP7_75t_L g448 ( .A1(n_423), .A2(n_309), .B(n_242), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_409), .B(n_272), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_424), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
BUFx10_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_409), .B(n_279), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_402), .A2(n_331), .B(n_304), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_430), .A2(n_283), .B(n_282), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_429), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_429), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_428), .A2(n_296), .B1(n_315), .B2(n_280), .Y(n_459) );
AOI21x1_ASAP7_75t_L g460 ( .A1(n_455), .A2(n_309), .B(n_350), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_452), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_426), .A2(n_342), .B1(n_333), .B2(n_287), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_443), .Y(n_463) );
OAI21x1_ASAP7_75t_L g464 ( .A1(n_448), .A2(n_15), .B(n_13), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_431), .B(n_6), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
AO221x2_ASAP7_75t_L g468 ( .A1(n_432), .A2(n_6), .B1(n_7), .B2(n_8), .C(n_9), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_435), .B(n_9), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_437), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_442), .B(n_360), .C(n_289), .Y(n_471) );
OAI21x1_ASAP7_75t_L g472 ( .A1(n_436), .A2(n_17), .B(n_21), .Y(n_472) );
BUFx8_ASAP7_75t_L g473 ( .A(n_447), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_433), .A2(n_434), .B(n_446), .Y(n_474) );
OAI21x1_ASAP7_75t_L g475 ( .A1(n_439), .A2(n_22), .B(n_23), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_440), .B(n_25), .Y(n_476) );
OAI21x1_ASAP7_75t_L g477 ( .A1(n_445), .A2(n_27), .B(n_28), .Y(n_477) );
AO31x2_ASAP7_75t_L g478 ( .A1(n_444), .A2(n_33), .A3(n_29), .B(n_30), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_444), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_454), .A2(n_295), .B(n_284), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_453), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_426), .A2(n_312), .B1(n_314), .B2(n_310), .Y(n_482) );
OAI21x1_ASAP7_75t_L g483 ( .A1(n_449), .A2(n_35), .B(n_37), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_428), .A2(n_322), .B1(n_326), .B2(n_321), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_429), .Y(n_486) );
CKINVDCx6p67_ASAP7_75t_R g487 ( .A(n_450), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_451), .B(n_330), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_455), .B(n_338), .C(n_337), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_450), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_451), .B(n_340), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_430), .A2(n_39), .B(n_41), .Y(n_492) );
OAI21x1_ASAP7_75t_L g493 ( .A1(n_441), .A2(n_42), .B(n_43), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_450), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_428), .A2(n_44), .B1(n_45), .B2(n_46), .C(n_47), .Y(n_495) );
NOR2xp67_ASAP7_75t_L g496 ( .A(n_427), .B(n_48), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_451), .B(n_50), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_470), .B(n_51), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_462), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_479), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_469), .B(n_56), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_466), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_463), .B(n_226), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_494), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_469), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_481), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_496), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_473), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_465), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_468), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_488), .B(n_58), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_468), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_491), .B(n_60), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_458), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_482), .B(n_61), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_486), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_484), .B(n_225), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_476), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_475), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_472), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_456), .B(n_63), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_460), .Y(n_528) );
INVx4_ASAP7_75t_L g529 ( .A(n_495), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_497), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_459), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_477), .B(n_66), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_483), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_493), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_471), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_492), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_480), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_461), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_476), .B(n_67), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_490), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_490), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_470), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
INVx4_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_470), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_476), .B(n_68), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_470), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_490), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_470), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_461), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_487), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_470), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_487), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_461), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_461), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_461), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_461), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_548), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_503), .B(n_69), .Y(n_564) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_512), .B(n_70), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_512), .B(n_224), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_507), .B(n_74), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_542), .B(n_76), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_542), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_505), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_500), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_510), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_552), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_541), .Y(n_574) );
BUFx3_ASAP7_75t_L g575 ( .A(n_558), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_546), .B(n_78), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_549), .B(n_79), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_548), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_551), .B(n_80), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_554), .B(n_81), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_557), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_502), .B(n_84), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_544), .B(n_85), .Y(n_583) );
INVxp67_ASAP7_75t_R g584 ( .A(n_501), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_545), .B(n_86), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_517), .Y(n_586) );
BUFx3_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_547), .B(n_223), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_520), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_543), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_553), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_555), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_513), .B(n_90), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_515), .B(n_222), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_521), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_523), .Y(n_597) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_550), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_559), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_556), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_506), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_560), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_561), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_562), .B(n_97), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_532), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_556), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_525), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_508), .B(n_98), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_518), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_531), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_530), .B(n_104), .Y(n_612) );
INVx6_ASAP7_75t_L g613 ( .A(n_519), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_538), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_509), .B(n_105), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_526), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_527), .B(n_107), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_498), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_540), .B(n_221), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_504), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_537), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_511), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_535), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_529), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_524), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_514), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_516), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_534), .Y(n_628) );
BUFx3_ASAP7_75t_L g629 ( .A(n_522), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_533), .Y(n_630) );
OR2x6_ASAP7_75t_L g631 ( .A(n_499), .B(n_111), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_539), .B(n_112), .Y(n_632) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_536), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_528), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_503), .B(n_115), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_500), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_500), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_603), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_596), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_606), .B(n_118), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_604), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_570), .B(n_119), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_624), .B(n_120), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_591), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_578), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_624), .B(n_123), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_614), .B(n_125), .Y(n_649) );
INVx4_ASAP7_75t_L g650 ( .A(n_573), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_592), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_596), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_602), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_602), .Y(n_654) );
NAND2x1_ASAP7_75t_L g655 ( .A(n_569), .B(n_127), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_571), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_611), .B(n_130), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_621), .B(n_132), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_571), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_599), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_636), .Y(n_661) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_598), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_600), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_597), .B(n_133), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_584), .B(n_138), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_637), .B(n_140), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_637), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_601), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_575), .Y(n_669) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_634), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_610), .B(n_141), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_572), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_622), .B(n_142), .Y(n_673) );
AND2x4_ASAP7_75t_SL g674 ( .A(n_563), .B(n_143), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_607), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_572), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_586), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_569), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_566), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_586), .B(n_589), .Y(n_680) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_623), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_595), .Y(n_682) );
INVx1_ASAP7_75t_SL g683 ( .A(n_587), .Y(n_683) );
AND2x4_ASAP7_75t_SL g684 ( .A(n_568), .B(n_146), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_595), .B(n_149), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_564), .B(n_150), .Y(n_686) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_627), .A2(n_151), .B1(n_152), .B2(n_154), .C1(n_156), .C2(n_158), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_588), .B(n_160), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_618), .B(n_161), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_590), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_635), .B(n_162), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_608), .Y(n_692) );
NAND2x1_ASAP7_75t_L g693 ( .A(n_565), .B(n_163), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_620), .B(n_164), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_626), .B(n_165), .Y(n_695) );
NAND2x1_ASAP7_75t_L g696 ( .A(n_568), .B(n_166), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_638), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_670), .B(n_616), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_645), .B(n_613), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_668), .B(n_613), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_682), .B(n_629), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_680), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_640), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_663), .B(n_582), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_681), .B(n_628), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_678), .B(n_630), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_675), .B(n_583), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_662), .B(n_625), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_652), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_653), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_656), .B(n_593), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_654), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_659), .B(n_594), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_661), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_667), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_672), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_679), .B(n_585), .Y(n_717) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_647), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_676), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_646), .B(n_609), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_677), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_692), .B(n_633), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_639), .B(n_615), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_642), .B(n_615), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_651), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_660), .B(n_576), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_683), .B(n_612), .Y(n_727) );
INVx3_ASAP7_75t_L g728 ( .A(n_690), .Y(n_728) );
BUFx3_ASAP7_75t_L g729 ( .A(n_650), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_690), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_690), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_666), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_649), .B(n_577), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_703), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_698), .B(n_669), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g736 ( .A(n_729), .B(n_696), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_697), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_714), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_715), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_699), .B(n_643), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_702), .B(n_641), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_719), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_718), .B(n_664), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_705), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_705), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_722), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_700), .B(n_687), .C(n_665), .D(n_673), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_701), .A2(n_696), .B(n_693), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_722), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_720), .B(n_686), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_708), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_721), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_708), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_709), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_711), .B(n_657), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_710), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_713), .B(n_666), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_712), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_746), .B(n_704), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_736), .A2(n_732), .B1(n_727), .B2(n_728), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_734), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_735), .Y(n_762) );
NOR2x1_ASAP7_75t_L g763 ( .A(n_748), .B(n_728), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_747), .A2(n_717), .B1(n_707), .B2(n_706), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_758), .Y(n_765) );
AOI222xp33_ASAP7_75t_L g766 ( .A1(n_755), .A2(n_726), .B1(n_723), .B2(n_724), .C1(n_706), .C2(n_733), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_737), .Y(n_767) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_743), .B(n_731), .C(n_730), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_738), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_749), .A2(n_648), .B1(n_644), .B2(n_684), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g771 ( .A(n_744), .B(n_644), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_761), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_764), .B(n_739), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_762), .A2(n_756), .B1(n_754), .B2(n_742), .C(n_752), .Y(n_774) );
NAND2xp33_ASAP7_75t_R g775 ( .A(n_759), .B(n_648), .Y(n_775) );
CKINVDCx14_ASAP7_75t_R g776 ( .A(n_770), .Y(n_776) );
OAI221xp5_ASAP7_75t_L g777 ( .A1(n_763), .A2(n_750), .B1(n_757), .B2(n_745), .C(n_753), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_765), .Y(n_778) );
AOI22xp5_ASAP7_75t_SL g779 ( .A1(n_771), .A2(n_740), .B1(n_751), .B2(n_691), .Y(n_779) );
AOI31xp33_ASAP7_75t_L g780 ( .A1(n_760), .A2(n_688), .A3(n_617), .B(n_741), .Y(n_780) );
AOI211xp5_ASAP7_75t_L g781 ( .A1(n_777), .A2(n_768), .B(n_769), .C(n_767), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_776), .A2(n_766), .B1(n_617), .B2(n_631), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_775), .A2(n_631), .B1(n_725), .B2(n_716), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_780), .A2(n_655), .B(n_674), .Y(n_784) );
O2A1O1Ixp33_ASAP7_75t_L g785 ( .A1(n_773), .A2(n_695), .B(n_694), .C(n_689), .Y(n_785) );
NAND2xp33_ASAP7_75t_SL g786 ( .A(n_779), .B(n_685), .Y(n_786) );
NOR3xp33_ASAP7_75t_L g787 ( .A(n_786), .B(n_774), .C(n_671), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_781), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_782), .B(n_772), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_783), .B(n_778), .Y(n_790) );
NOR4xp25_ASAP7_75t_L g791 ( .A(n_788), .B(n_785), .C(n_579), .D(n_658), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_789), .B(n_784), .Y(n_792) );
NOR2xp67_ASAP7_75t_L g793 ( .A(n_792), .B(n_790), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_791), .B(n_787), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_793), .B(n_580), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_794), .B(n_619), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_795), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_796), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_798), .Y(n_799) );
XOR2x1_ASAP7_75t_L g800 ( .A(n_797), .B(n_567), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_799), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_801), .A2(n_800), .B(n_605), .Y(n_802) );
OR2x6_ASAP7_75t_L g803 ( .A(n_802), .B(n_632), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_803), .B(n_170), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_804), .A2(n_173), .B1(n_174), .B2(n_176), .C(n_177), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_805), .A2(n_182), .B1(n_183), .B2(n_185), .Y(n_806) );
endmodule