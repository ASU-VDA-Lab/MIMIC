module fake_jpeg_28943_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_45),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_29),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_9),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_43),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_26),
.B1(n_23),
.B2(n_18),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_21),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_24),
.B1(n_17),
.B2(n_19),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_34),
.A2(n_29),
.B1(n_19),
.B2(n_3),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_29),
.C(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_47),
.B1(n_66),
.B2(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_29),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_3),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_90),
.Y(n_108)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_91),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_99),
.B1(n_102),
.B2(n_109),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_75),
.B(n_90),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_66),
.B1(n_69),
.B2(n_54),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_48),
.C(n_5),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_83),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_54),
.B1(n_61),
.B2(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_61),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_122),
.B(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_71),
.C(n_70),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_124),
.C(n_77),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_80),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_70),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_92),
.B(n_91),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_106),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_124),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_104),
.C(n_76),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_128),
.C(n_127),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_75),
.B(n_95),
.C(n_99),
.D(n_109),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_103),
.B(n_96),
.C(n_4),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_139),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_118),
.C(n_110),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_78),
.C(n_86),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_116),
.B1(n_87),
.B2(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_116),
.B1(n_84),
.B2(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_130),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_126),
.B(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_153),
.C(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_139),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_145),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_147),
.B1(n_145),
.B2(n_6),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_158),
.Y(n_163)
);

OAI31xp33_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_145),
.A3(n_11),
.B(n_14),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_164),
.B(n_162),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_160),
.C(n_164),
.Y(n_167)
);


endmodule