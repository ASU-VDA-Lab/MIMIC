module fake_jpeg_222_n_672 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_672);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_672;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_59),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_60),
.B(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_62),
.Y(n_218)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_26),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g144 ( 
.A(n_67),
.Y(n_144)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_73),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_1),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_76),
.A2(n_46),
.B(n_27),
.C(n_56),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_81),
.B(n_124),
.Y(n_154)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_93),
.Y(n_143)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_87),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

CKINVDCx9p33_ASAP7_75t_R g91 ( 
.A(n_23),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g173 ( 
.A(n_91),
.Y(n_173)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_3),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_94),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_98),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_105),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_31),
.B(n_3),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_119),
.Y(n_147)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_109),
.Y(n_215)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_111),
.Y(n_198)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_117),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_28),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_31),
.B(n_3),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_126),
.Y(n_230)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_41),
.B(n_46),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_32),
.Y(n_164)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_76),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_133),
.B(n_149),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_78),
.A2(n_22),
.B1(n_27),
.B2(n_56),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_134),
.A2(n_155),
.B1(n_162),
.B2(n_174),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_142),
.B(n_150),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_77),
.B(n_22),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_67),
.B(n_22),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_151),
.B(n_164),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_103),
.A2(n_32),
.B1(n_36),
.B2(n_56),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_28),
.B(n_57),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_158),
.B(n_15),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_107),
.A2(n_54),
.B1(n_36),
.B2(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_59),
.B(n_36),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_171),
.B(n_185),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_61),
.A2(n_54),
.B1(n_57),
.B2(n_55),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_114),
.B(n_54),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_179),
.B(n_18),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_59),
.A2(n_40),
.B1(n_57),
.B2(n_55),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_183),
.A2(n_192),
.B1(n_193),
.B2(n_228),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_62),
.B(n_55),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_62),
.B(n_51),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_191),
.B(n_195),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_86),
.A2(n_28),
.B1(n_51),
.B2(n_45),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_86),
.A2(n_40),
.B1(n_51),
.B2(n_45),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_64),
.B(n_45),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_70),
.A2(n_43),
.B1(n_40),
.B2(n_34),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_199),
.A2(n_202),
.B1(n_216),
.B2(n_217),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_72),
.A2(n_43),
.B1(n_34),
.B2(n_39),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_82),
.Y(n_211)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_74),
.A2(n_43),
.B1(n_34),
.B2(n_39),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_214),
.A2(n_223),
.B1(n_18),
.B2(n_11),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_75),
.A2(n_58),
.B1(n_39),
.B2(n_35),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_83),
.A2(n_58),
.B1(n_39),
.B2(n_35),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_87),
.B(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_219),
.B(n_229),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_88),
.A2(n_102),
.B1(n_121),
.B2(n_113),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_221),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_94),
.A2(n_58),
.B1(n_39),
.B2(n_35),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_122),
.A2(n_58),
.B1(n_39),
.B2(n_35),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_95),
.B(n_4),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_231),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_109),
.B(n_108),
.C(n_101),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_232),
.A2(n_280),
.B(n_231),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_234),
.B(n_237),
.Y(n_330)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_157),
.Y(n_235)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_235),
.Y(n_346)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_230),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_238),
.Y(n_337)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_239),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_240),
.Y(n_349)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_241),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_243),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_244),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_141),
.B(n_99),
.C(n_58),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_315),
.C(n_217),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_175),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_247),
.B(n_290),
.Y(n_358)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_197),
.A2(n_35),
.B1(n_30),
.B2(n_6),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_250),
.A2(n_253),
.B1(n_254),
.B2(n_276),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_251),
.B(n_277),
.Y(n_339)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_143),
.A2(n_35),
.B1(n_30),
.B2(n_6),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_147),
.A2(n_30),
.B1(n_5),
.B2(n_6),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_136),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_259),
.Y(n_353)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_260),
.Y(n_355)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_261),
.Y(n_359)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_166),
.Y(n_262)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_262),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_188),
.B(n_189),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_263),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_132),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_265),
.B(n_284),
.Y(n_344)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_266),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_267),
.A2(n_194),
.B1(n_177),
.B2(n_181),
.Y(n_329)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_176),
.Y(n_268)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_269),
.Y(n_371)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_270),
.Y(n_374)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_184),
.Y(n_272)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_275),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_212),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_278),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_140),
.B(n_8),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_279),
.B(n_281),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_162),
.A2(n_8),
.B(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_137),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_294),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_189),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_139),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_285),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_223),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_145),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_289),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_154),
.B(n_11),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_138),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_296),
.Y(n_375)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

CKINVDCx12_ASAP7_75t_R g325 ( 
.A(n_293),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_146),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g297 ( 
.A(n_153),
.B(n_16),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_297),
.A2(n_298),
.B(n_238),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_226),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_300),
.Y(n_316)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_301),
.A2(n_310),
.B1(n_311),
.B2(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_305),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_148),
.B(n_152),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_303),
.A2(n_306),
.B1(n_312),
.B2(n_153),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_156),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_180),
.B(n_165),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_168),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_309),
.Y(n_360)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_200),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_174),
.B(n_169),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_159),
.B(n_169),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_159),
.B(n_177),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_221),
.A2(n_213),
.B1(n_190),
.B2(n_135),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_314),
.A2(n_298),
.B1(n_249),
.B2(n_270),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_SL g315 ( 
.A(n_132),
.B(n_209),
.C(n_228),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_134),
.B(n_192),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_320),
.B(n_323),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_324),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_304),
.A2(n_135),
.B1(n_215),
.B2(n_207),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_326),
.A2(n_327),
.B1(n_329),
.B2(n_364),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_207),
.B1(n_215),
.B2(n_178),
.Y(n_327)
);

AOI22x1_ASAP7_75t_SL g328 ( 
.A1(n_295),
.A2(n_183),
.B1(n_193),
.B2(n_178),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_328),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_296),
.A2(n_165),
.B(n_220),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_331),
.A2(n_342),
.B(n_324),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_282),
.A2(n_216),
.B1(n_227),
.B2(n_194),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_338),
.A2(n_340),
.B1(n_354),
.B2(n_305),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_246),
.A2(n_227),
.B1(n_181),
.B2(n_182),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_288),
.A2(n_182),
.B(n_220),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_280),
.A2(n_308),
.B1(n_301),
.B2(n_274),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_292),
.B(n_245),
.C(n_242),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_334),
.C(n_344),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_232),
.A2(n_236),
.B1(n_275),
.B2(n_309),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_373),
.B1(n_241),
.B2(n_244),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_312),
.A2(n_255),
.B1(n_252),
.B2(n_269),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_366),
.A2(n_368),
.B1(n_247),
.B2(n_260),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_256),
.A2(n_262),
.B1(n_273),
.B2(n_271),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_356),
.Y(n_378)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_320),
.A2(n_297),
.B(n_263),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_379),
.A2(n_390),
.B(n_422),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_375),
.B(n_257),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_380),
.B(n_382),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_354),
.B(n_263),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_381),
.B(n_372),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_233),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_264),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_383),
.Y(n_436)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_248),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_385),
.B(n_396),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_386),
.A2(n_394),
.B1(n_395),
.B2(n_401),
.Y(n_430)
);

AO21x2_ASAP7_75t_L g387 ( 
.A1(n_340),
.A2(n_259),
.B(n_285),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_387),
.A2(n_406),
.B1(n_409),
.B2(n_346),
.Y(n_447)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

AOI21xp33_ASAP7_75t_L g390 ( 
.A1(n_369),
.A2(n_342),
.B(n_365),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_290),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_408),
.C(n_421),
.Y(n_439)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_327),
.A2(n_243),
.B1(n_300),
.B2(n_235),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_326),
.A2(n_266),
.B1(n_261),
.B2(n_239),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_316),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_397),
.B(n_318),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_316),
.B(n_251),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_403),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_330),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_416),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_320),
.A2(n_307),
.B1(n_278),
.B2(n_293),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_334),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_404),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_338),
.A2(n_343),
.B1(n_336),
.B2(n_328),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_407),
.B(n_419),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_363),
.A2(n_347),
.B1(n_370),
.B2(n_319),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_370),
.B(n_339),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_417),
.Y(n_453)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_411),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_337),
.A2(n_358),
.B(n_317),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_361),
.B(n_367),
.Y(n_429)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_349),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_332),
.B(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_420),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_351),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_350),
.B(n_371),
.C(n_374),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_317),
.A2(n_325),
.B(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_424),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_348),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_353),
.A2(n_348),
.B1(n_367),
.B2(n_361),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_426),
.A2(n_353),
.B1(n_341),
.B2(n_335),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_390),
.A2(n_355),
.B(n_359),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_427),
.A2(n_429),
.B(n_442),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_434),
.A2(n_445),
.B1(n_461),
.B2(n_465),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_392),
.B(n_341),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_438),
.B(n_441),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_382),
.B(n_335),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_438),
.C(n_439),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_385),
.B(n_380),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_405),
.A2(n_362),
.B(n_376),
.Y(n_442)
);

XOR2x2_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_376),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_444),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_401),
.A2(n_346),
.B1(n_353),
.B2(n_318),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_410),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_454),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_447),
.A2(n_415),
.B1(n_394),
.B2(n_384),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_383),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_457),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_389),
.B(n_372),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_460),
.B(n_398),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_321),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_416),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_391),
.A2(n_321),
.B(n_322),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_463),
.A2(n_422),
.B(n_413),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_388),
.A2(n_322),
.B1(n_403),
.B2(n_399),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_406),
.A2(n_386),
.B1(n_387),
.B2(n_378),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_466),
.A2(n_387),
.B1(n_415),
.B2(n_422),
.Y(n_498)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_443),
.Y(n_474)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_475),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_437),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_476),
.B(n_479),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_477),
.A2(n_496),
.B1(n_498),
.B2(n_506),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_412),
.C(n_408),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_478),
.B(n_483),
.C(n_490),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_437),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_455),
.A2(n_412),
.B1(n_387),
.B2(n_379),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_480),
.A2(n_488),
.B1(n_505),
.B2(n_463),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_449),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_482),
.B(n_493),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_435),
.C(n_444),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_381),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_484),
.B(n_453),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_485),
.Y(n_542)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_486),
.Y(n_525)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_455),
.A2(n_387),
.B1(n_396),
.B2(n_409),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_464),
.Y(n_489)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_435),
.B(n_404),
.C(n_421),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_492),
.A2(n_428),
.B(n_427),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_449),
.Y(n_493)
);

CKINVDCx14_ASAP7_75t_R g509 ( 
.A(n_494),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_444),
.B(n_411),
.C(n_417),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_495),
.B(n_502),
.C(n_442),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_466),
.A2(n_447),
.B1(n_452),
.B2(n_451),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

AND2x4_ASAP7_75t_SL g499 ( 
.A(n_460),
.B(n_418),
.Y(n_499)
);

CKINVDCx14_ASAP7_75t_R g532 ( 
.A(n_499),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_420),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_414),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_504),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_450),
.B(n_423),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_425),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_430),
.A2(n_387),
.B1(n_395),
.B2(n_393),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_451),
.A2(n_426),
.B1(n_452),
.B2(n_431),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_507),
.A2(n_520),
.B1(n_524),
.B2(n_534),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_501),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_510),
.B(n_511),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_468),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_468),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_512),
.B(n_513),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_499),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_441),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_527),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_486),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_515),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_429),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_518),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_480),
.A2(n_432),
.B1(n_428),
.B2(n_433),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_523),
.B(n_469),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_496),
.A2(n_431),
.B1(n_433),
.B2(n_430),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_477),
.A2(n_465),
.B1(n_448),
.B2(n_461),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_526),
.A2(n_497),
.B1(n_505),
.B2(n_487),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_448),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_530),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_490),
.B(n_453),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_488),
.A2(n_461),
.B1(n_462),
.B2(n_427),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_470),
.B(n_467),
.C(n_464),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_535),
.B(n_543),
.C(n_495),
.Y(n_548)
);

AOI22x1_ASAP7_75t_L g540 ( 
.A1(n_491),
.A2(n_436),
.B1(n_467),
.B2(n_456),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_540),
.A2(n_506),
.B1(n_499),
.B2(n_472),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_470),
.B(n_483),
.Y(n_543)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_508),
.Y(n_545)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_545),
.Y(n_575)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_548),
.B(n_526),
.Y(n_591)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_517),
.Y(n_550)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_550),
.Y(n_579)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_533),
.Y(n_551)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_551),
.Y(n_584)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_534),
.A2(n_491),
.B(n_481),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_552),
.A2(n_554),
.B(n_523),
.Y(n_583)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_553),
.Y(n_587)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_525),
.Y(n_555)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_555),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_522),
.B(n_471),
.C(n_474),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_556),
.B(n_563),
.C(n_564),
.Y(n_574)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_525),
.Y(n_557)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_557),
.Y(n_597)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_560),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_562),
.A2(n_539),
.B1(n_537),
.B2(n_542),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_522),
.B(n_502),
.C(n_500),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_514),
.C(n_543),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_519),
.B(n_504),
.C(n_472),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_565),
.B(n_572),
.C(n_527),
.Y(n_581)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_541),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_566),
.B(n_568),
.Y(n_576)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_569),
.B(n_573),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_570),
.A2(n_507),
.B1(n_524),
.B2(n_518),
.Y(n_580)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_536),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_571),
.B(n_489),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_528),
.B(n_469),
.C(n_475),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_577),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_580),
.A2(n_590),
.B1(n_595),
.B2(n_573),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_591),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_554),
.A2(n_540),
.B(n_516),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_582),
.A2(n_583),
.B(n_594),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_567),
.B(n_509),
.Y(n_585)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_585),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_549),
.B(n_530),
.C(n_535),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_589),
.C(n_593),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_549),
.B(n_540),
.C(n_521),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_570),
.A2(n_532),
.B1(n_516),
.B2(n_539),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_592),
.A2(n_544),
.B1(n_551),
.B2(n_560),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_564),
.B(n_503),
.C(n_529),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_544),
.A2(n_552),
.B(n_547),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_545),
.A2(n_546),
.B1(n_557),
.B2(n_555),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_585),
.B(n_559),
.Y(n_599)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_576),
.A2(n_561),
.B1(n_552),
.B2(n_550),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_602),
.A2(n_595),
.B1(n_597),
.B2(n_588),
.Y(n_625)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_577),
.Y(n_604)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_604),
.Y(n_632)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_606),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_576),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_607),
.B(n_611),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_594),
.A2(n_544),
.B(n_572),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_616),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_609),
.A2(n_575),
.B1(n_578),
.B2(n_588),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_563),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_612),
.Y(n_629)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_596),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_582),
.A2(n_565),
.B(n_556),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_558),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_614),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_583),
.A2(n_569),
.B(n_558),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_581),
.B(n_591),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_593),
.B(n_548),
.C(n_553),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_617),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_574),
.B(n_586),
.C(n_580),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_618),
.B(n_590),
.C(n_592),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_619),
.B(n_623),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_621),
.A2(n_625),
.B1(n_606),
.B2(n_603),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_617),
.B(n_575),
.C(n_578),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_618),
.B(n_616),
.C(n_605),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_624),
.B(n_626),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_601),
.B(n_587),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_600),
.Y(n_628)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_628),
.Y(n_641)
);

NOR2x1_ASAP7_75t_L g633 ( 
.A(n_614),
.B(n_597),
.Y(n_633)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_633),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_605),
.B(n_587),
.C(n_596),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_635),
.B(n_598),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_636),
.B(n_638),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_633),
.A2(n_603),
.B(n_612),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_637),
.A2(n_645),
.B(n_622),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_635),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_630),
.B(n_615),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_643),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_632),
.A2(n_599),
.B1(n_598),
.B2(n_609),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_622),
.A2(n_615),
.B(n_608),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_624),
.B(n_613),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_646),
.B(n_647),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_620),
.B(n_610),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_648),
.B(n_623),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_644),
.A2(n_628),
.B(n_631),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_649),
.A2(n_656),
.B(n_657),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_638),
.B(n_627),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_651),
.B(n_640),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_653),
.Y(n_661)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_655),
.A2(n_641),
.B(n_639),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_SL g656 ( 
.A1(n_642),
.A2(n_630),
.B(n_634),
.Y(n_656)
);

OAI21xp33_ASAP7_75t_L g657 ( 
.A1(n_637),
.A2(n_619),
.B(n_629),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g664 ( 
.A(n_659),
.B(n_660),
.C(n_662),
.Y(n_664)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_654),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_650),
.A2(n_629),
.B(n_636),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_663),
.A2(n_650),
.B(n_652),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_665),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_658),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_666),
.A2(n_661),
.B(n_579),
.Y(n_668)
);

BUFx24_ASAP7_75t_SL g669 ( 
.A(n_668),
.Y(n_669)
);

NAND2x1_ASAP7_75t_L g670 ( 
.A(n_669),
.B(n_664),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_670),
.A2(n_667),
.B(n_579),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_671),
.A2(n_584),
.B(n_668),
.Y(n_672)
);


endmodule