module fake_jpeg_26321_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_15;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_67;
wire n_66;

BUFx12_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_22),
.Y(n_33)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_14),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_22),
.B(n_25),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_17),
.B1(n_18),
.B2(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_10),
.B1(n_13),
.B2(n_11),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_38),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_24),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_11),
.B1(n_10),
.B2(n_16),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_6),
.C(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_47),
.B(n_14),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_14),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_41),
.B1(n_30),
.B2(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

AOI22x1_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_54)
);

XOR2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_31),
.B1(n_36),
.B2(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_44),
.C(n_48),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_46),
.C(n_54),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.C(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_51),
.C(n_21),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_21),
.C(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_3),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_69),
.Y(n_73)
);


endmodule