module fake_jpeg_3004_n_59 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_59);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx9p33_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_22),
.Y(n_24)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_19),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_21),
.B1(n_19),
.B2(n_8),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_1),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_21),
.C(n_33),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_39),
.B(n_2),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_31),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_26),
.B1(n_27),
.B2(n_4),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_3),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_7),
.C(n_12),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_50),
.B(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_5),
.C(n_6),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_49),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);


endmodule