module fake_jpeg_6589_n_103 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_1),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_62),
.B1(n_55),
.B2(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_75),
.B1(n_51),
.B2(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_51),
.B1(n_50),
.B2(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_77),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_57),
.B1(n_43),
.B2(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_58),
.B1(n_59),
.B2(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_5),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_38),
.B1(n_12),
.B2(n_13),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_41),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.C(n_90),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_11),
.B(n_19),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_88),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_91),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_20),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_26),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_27),
.C(n_28),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_35),
.Y(n_103)
);


endmodule