module fake_jpeg_3771_n_213 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_213);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_36),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_14),
.B(n_24),
.Y(n_34)
);

OR2x4_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_41),
.Y(n_78)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_40),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_28),
.B1(n_15),
.B2(n_17),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_72),
.B1(n_12),
.B2(n_11),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_27),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_1),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_70),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_21),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_75),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_20),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_22),
.B1(n_18),
.B2(n_12),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_78),
.B1(n_54),
.B2(n_65),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_107),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_26),
.B(n_24),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_59),
.B(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_88),
.B(n_89),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_104),
.B1(n_65),
.B2(n_73),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_3),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_80),
.C(n_76),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_114),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_112),
.Y(n_138)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_50),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_80),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_121),
.B1(n_133),
.B2(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_R g119 ( 
.A(n_93),
.B(n_100),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_48),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_55),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_91),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_121),
.C(n_125),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_89),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_123),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_149),
.B(n_153),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_92),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_99),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_54),
.B1(n_47),
.B2(n_52),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_103),
.B(n_55),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_135),
.C(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_123),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_146),
.B(n_123),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_142),
.B(n_145),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_181),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_134),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_153),
.B1(n_149),
.B2(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_157),
.C(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_160),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_182),
.C(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_186),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_178),
.B(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_139),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_170),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_192),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_173),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_183),
.B(n_181),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_188),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_203),
.B(n_193),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_143),
.B(n_187),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_144),
.C(n_150),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_198),
.B(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_153),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_195),
.A3(n_167),
.B1(n_187),
.B2(n_153),
.C1(n_162),
.C2(n_171),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_109),
.C(n_140),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_210),
.B1(n_90),
.B2(n_6),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_206),
.C(n_58),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_212),
.Y(n_213)
);


endmodule