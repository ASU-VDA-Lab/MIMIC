module fake_netlist_6_3165_n_779 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_779);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_779;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_683;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_44),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_46),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_20),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_29),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_5),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_51),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_45),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_49),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_66),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_97),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_94),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_34),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_69),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_106),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_18),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_65),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_89),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_103),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_96),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_11),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_113),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_5),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_42),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_0),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_100),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_8),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_73),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_81),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_78),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_139),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_114),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_0),
.Y(n_209)
);

AND2x4_ASAP7_75t_SL g210 ( 
.A(n_161),
.B(n_23),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_24),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_1),
.Y(n_212)
);

CKINVDCx6p67_ASAP7_75t_R g213 ( 
.A(n_158),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_1),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_2),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_151),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_149),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_164),
.B(n_165),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_162),
.B(n_2),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_3),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_3),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_4),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_169),
.B(n_6),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_6),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_150),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_185),
.B1(n_161),
.B2(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_172),
.B1(n_197),
.B2(n_152),
.Y(n_247)
);

AO22x2_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_208),
.B1(n_211),
.B2(n_238),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_152),
.B1(n_200),
.B2(n_198),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_200),
.B1(n_201),
.B2(n_193),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_206),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_209),
.A2(n_190),
.B1(n_188),
.B2(n_184),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_7),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_180),
.B1(n_179),
.B2(n_178),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_182),
.B1(n_177),
.B2(n_174),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_213),
.A2(n_173),
.B1(n_10),
.B2(n_11),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_214),
.B1(n_239),
.B2(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_25),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_208),
.B(n_26),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_235),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_27),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_211),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_31),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_32),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_16),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_236),
.A2(n_218),
.B1(n_210),
.B2(n_211),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_R g278 ( 
.A(n_223),
.B(n_145),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g280 ( 
.A1(n_205),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_19),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_210),
.A2(n_205),
.B1(n_222),
.B2(n_223),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_33),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_232),
.A2(n_207),
.B1(n_216),
.B2(n_21),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_207),
.B(n_21),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_216),
.A2(n_22),
.B1(n_35),
.B2(n_37),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_243),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_216),
.B(n_22),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_224),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_224),
.A2(n_41),
.B1(n_43),
.B2(n_47),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_48),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_224),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

BUFx6f_ASAP7_75t_SL g299 ( 
.A(n_264),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_50),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_52),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_225),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_248),
.B(n_225),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_221),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_53),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_271),
.B(n_221),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_247),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_277),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_225),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_250),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_225),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_251),
.B(n_225),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_250),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_221),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_260),
.B(n_221),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_L g338 ( 
.A(n_249),
.B(n_221),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_270),
.Y(n_340)
);

XNOR2x2_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_54),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_251),
.B(n_55),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_261),
.B(n_228),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_259),
.B(n_258),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_259),
.Y(n_347)
);

XNOR2x2_ASAP7_75t_L g348 ( 
.A(n_272),
.B(n_56),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_253),
.A2(n_230),
.B(n_228),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_292),
.B(n_228),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_227),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_269),
.B(n_227),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_255),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_237),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_296),
.B(n_237),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_230),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_310),
.B(n_57),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_230),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_298),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_58),
.Y(n_372)
);

BUFx4f_ASAP7_75t_SL g373 ( 
.A(n_322),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_345),
.A2(n_328),
.B(n_336),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_359),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_318),
.B(n_230),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_356),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_59),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_60),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_237),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_324),
.B(n_332),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_294),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_328),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_337),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_237),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_326),
.B(n_237),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_326),
.B(n_230),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_327),
.B(n_227),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_359),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_347),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_359),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_312),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_305),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_306),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_302),
.Y(n_411)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g413 ( 
.A(n_346),
.B(n_227),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_61),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_314),
.B(n_345),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_343),
.B(n_233),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_334),
.B(n_62),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_343),
.B(n_227),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_314),
.B(n_230),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_351),
.A2(n_231),
.B(n_228),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_316),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_314),
.B(n_228),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_346),
.B(n_233),
.Y(n_424)
);

AND2x2_ASAP7_75t_SL g425 ( 
.A(n_352),
.B(n_233),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_63),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_314),
.B(n_231),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_314),
.B(n_231),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_314),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_366),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_394),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_373),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_361),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_393),
.B(n_330),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_344),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_386),
.B(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_385),
.B(n_317),
.Y(n_446)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_413),
.B(n_317),
.Y(n_447)
);

NAND2x1p5_ASAP7_75t_L g448 ( 
.A(n_365),
.B(n_333),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_353),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_398),
.B(n_333),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_374),
.B(n_314),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_354),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_367),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_323),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_390),
.B(n_320),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_391),
.B(n_323),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_365),
.B(n_349),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g465 ( 
.A(n_365),
.B(n_355),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_322),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_365),
.B(n_202),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_381),
.B(n_342),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_403),
.B(n_335),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_395),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_395),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_300),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_388),
.B(n_424),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_410),
.B(n_411),
.Y(n_480)
);

OR2x6_ASAP7_75t_SL g481 ( 
.A(n_411),
.B(n_348),
.Y(n_481)
);

NAND2x1p5_ASAP7_75t_L g482 ( 
.A(n_372),
.B(n_202),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_382),
.B(n_202),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_414),
.B(n_299),
.Y(n_484)
);

AO21x2_ASAP7_75t_L g485 ( 
.A1(n_416),
.A2(n_319),
.B(n_303),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_417),
.B(n_229),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_429),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_480),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_443),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_437),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_439),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_441),
.B(n_417),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_413),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_419),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_444),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_436),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_466),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_452),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_457),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_437),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_468),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_382),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

BUFx8_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_478),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_458),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

CKINVDCx8_ASAP7_75t_R g519 ( 
.A(n_433),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_382),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_455),
.Y(n_521)
);

CKINVDCx11_ASAP7_75t_R g522 ( 
.A(n_481),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_438),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_447),
.A2(n_413),
.B1(n_383),
.B2(n_382),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

CKINVDCx11_ASAP7_75t_R g527 ( 
.A(n_442),
.Y(n_527)
);

BUFx16f_ASAP7_75t_R g528 ( 
.A(n_442),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_474),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_419),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_459),
.B(n_447),
.Y(n_533)
);

BUFx2_ASAP7_75t_SL g534 ( 
.A(n_440),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_518),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_499),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_488),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_517),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_518),
.Y(n_539)
);

CKINVDCx11_ASAP7_75t_R g540 ( 
.A(n_508),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_505),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g545 ( 
.A1(n_533),
.A2(n_461),
.B1(n_475),
.B2(n_459),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_516),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_525),
.A2(n_475),
.B1(n_461),
.B2(n_472),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_496),
.B(n_446),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_498),
.A2(n_470),
.B1(n_485),
.B2(n_348),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_505),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_521),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_491),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_497),
.A2(n_460),
.B1(n_464),
.B2(n_470),
.Y(n_553)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_506),
.B(n_477),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_527),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_515),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_510),
.A2(n_485),
.B1(n_457),
.B2(n_383),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_510),
.A2(n_457),
.B1(n_383),
.B2(n_450),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_508),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_510),
.A2(n_464),
.B1(n_448),
.B2(n_520),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_530),
.A2(n_457),
.B1(n_425),
.B2(n_464),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_517),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_487),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_489),
.A2(n_460),
.B1(n_463),
.B2(n_444),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_522),
.A2(n_457),
.B1(n_425),
.B2(n_414),
.Y(n_565)
);

OAI22xp33_ASAP7_75t_L g566 ( 
.A1(n_510),
.A2(n_463),
.B1(n_471),
.B2(n_473),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_493),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_522),
.A2(n_425),
.B1(n_414),
.B2(n_426),
.Y(n_568)
);

BUFx4f_ASAP7_75t_SL g569 ( 
.A(n_524),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_506),
.B(n_477),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_L g571 ( 
.A1(n_531),
.A2(n_454),
.B(n_448),
.Y(n_571)
);

INVx6_ASAP7_75t_L g572 ( 
.A(n_513),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_454),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_492),
.A2(n_418),
.B1(n_426),
.B2(n_384),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_520),
.A2(n_465),
.B1(n_483),
.B2(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_495),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_549),
.A2(n_545),
.B1(n_548),
.B2(n_568),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_551),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_572),
.A2(n_503),
.B1(n_501),
.B2(n_513),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_542),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_568),
.A2(n_519),
.B1(n_509),
.B2(n_465),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_540),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_536),
.B(n_534),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_552),
.Y(n_585)
);

BUFx4f_ASAP7_75t_SL g586 ( 
.A(n_559),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_550),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_545),
.A2(n_553),
.B1(n_565),
.B2(n_547),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_565),
.A2(n_519),
.B1(n_509),
.B2(n_504),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_567),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_553),
.A2(n_501),
.B1(n_503),
.B2(n_507),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_556),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_535),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_564),
.A2(n_504),
.B1(n_493),
.B2(n_557),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

OAI211xp5_ASAP7_75t_SL g597 ( 
.A1(n_564),
.A2(n_527),
.B(n_421),
.C(n_370),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_561),
.A2(n_576),
.B1(n_574),
.B2(n_536),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_561),
.A2(n_370),
.B1(n_368),
.B2(n_426),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_537),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_539),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_574),
.A2(n_368),
.B1(n_418),
.B2(n_426),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_572),
.A2(n_418),
.B1(n_513),
.B2(n_384),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_563),
.B(n_523),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_418),
.B1(n_484),
.B2(n_412),
.Y(n_605)
);

BUFx4f_ASAP7_75t_SL g606 ( 
.A(n_555),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_538),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_544),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_500),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_571),
.A2(n_484),
.B1(n_412),
.B2(n_456),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_562),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_558),
.A2(n_299),
.B1(n_529),
.B2(n_506),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_566),
.A2(n_484),
.B1(n_412),
.B2(n_456),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_569),
.A2(n_506),
.B1(n_484),
.B2(n_299),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_569),
.A2(n_506),
.B1(n_484),
.B2(n_528),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_562),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_566),
.Y(n_620)
);

INVx6_ASAP7_75t_L g621 ( 
.A(n_550),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_575),
.A2(n_430),
.B(n_486),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_560),
.A2(n_412),
.B1(n_402),
.B2(n_400),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_543),
.A2(n_412),
.B1(n_402),
.B2(n_400),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_543),
.A2(n_412),
.B1(n_401),
.B2(n_430),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_550),
.A2(n_467),
.B1(n_482),
.B2(n_483),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_383),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_588),
.A2(n_412),
.B1(n_401),
.B2(n_363),
.Y(n_630)
);

AOI21xp33_ASAP7_75t_SL g631 ( 
.A1(n_589),
.A2(n_570),
.B(n_554),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_588),
.A2(n_467),
.B1(n_500),
.B2(n_550),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_577),
.A2(n_412),
.B1(n_363),
.B2(n_360),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_577),
.A2(n_592),
.B1(n_595),
.B2(n_597),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_580),
.B(n_532),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_578),
.B(n_360),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_581),
.A2(n_614),
.B1(n_586),
.B2(n_611),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_593),
.B(n_583),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_592),
.A2(n_396),
.B1(n_375),
.B2(n_378),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_598),
.A2(n_396),
.B1(n_375),
.B2(n_378),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_584),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_598),
.A2(n_490),
.B1(n_494),
.B2(n_502),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_599),
.A2(n_490),
.B1(n_494),
.B2(n_502),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_604),
.B(n_490),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_582),
.A2(n_415),
.B1(n_494),
.B2(n_502),
.Y(n_645)
);

AO22x1_ASAP7_75t_L g646 ( 
.A1(n_587),
.A2(n_532),
.B1(n_517),
.B2(n_415),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_618),
.A2(n_603),
.B1(n_602),
.B2(n_599),
.Y(n_647)
);

OAI221xp5_ASAP7_75t_L g648 ( 
.A1(n_603),
.A2(n_486),
.B1(n_422),
.B2(n_377),
.C(n_409),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_602),
.A2(n_409),
.B1(n_408),
.B2(n_404),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_585),
.B(n_532),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_594),
.B(n_517),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_579),
.A2(n_570),
.B1(n_554),
.B2(n_526),
.Y(n_652)
);

OAI21xp33_ASAP7_75t_L g653 ( 
.A1(n_623),
.A2(n_409),
.B(n_408),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_623),
.A2(n_404),
.B1(n_367),
.B2(n_369),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_621),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_621),
.A2(n_606),
.B1(n_600),
.B2(n_587),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_612),
.A2(n_364),
.B1(n_397),
.B2(n_233),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_616),
.A2(n_526),
.B1(n_512),
.B2(n_511),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_612),
.A2(n_233),
.B1(n_229),
.B2(n_462),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_621),
.A2(n_512),
.B1(n_511),
.B2(n_505),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_616),
.A2(n_229),
.B1(n_462),
.B2(n_431),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_601),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_613),
.B(n_229),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_615),
.B(n_67),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_627),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_625),
.A2(n_229),
.B1(n_462),
.B2(n_431),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_641),
.B(n_607),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_638),
.B(n_608),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_644),
.B(n_609),
.Y(n_669)
);

AOI221xp5_ASAP7_75t_L g670 ( 
.A1(n_634),
.A2(n_600),
.B1(n_610),
.B2(n_628),
.C(n_622),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_645),
.C(n_639),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_641),
.B(n_619),
.Y(n_672)
);

OAI221xp5_ASAP7_75t_SL g673 ( 
.A1(n_633),
.A2(n_605),
.B1(n_625),
.B2(n_624),
.C(n_617),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_640),
.B(n_624),
.C(n_605),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_665),
.B(n_619),
.Y(n_675)
);

AOI221xp5_ASAP7_75t_L g676 ( 
.A1(n_647),
.A2(n_590),
.B1(n_626),
.B2(n_591),
.C(n_596),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_596),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_662),
.B(n_596),
.Y(n_678)
);

AND4x1_ASAP7_75t_L g679 ( 
.A(n_630),
.B(n_661),
.C(n_666),
.D(n_642),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_665),
.B(n_596),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_635),
.B(n_591),
.Y(n_681)
);

NAND4xp25_ASAP7_75t_L g682 ( 
.A(n_656),
.B(n_526),
.C(n_512),
.D(n_511),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_635),
.B(n_591),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_650),
.B(n_591),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_650),
.B(n_68),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_655),
.B(n_431),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_629),
.B(n_70),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_629),
.B(n_72),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_649),
.A2(n_376),
.B1(n_407),
.B2(n_405),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_SL g690 ( 
.A1(n_631),
.A2(n_74),
.B(n_75),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_651),
.B(n_76),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_636),
.B(n_664),
.Y(n_692)
);

NOR2x1_ASAP7_75t_L g693 ( 
.A(n_680),
.B(n_655),
.Y(n_693)
);

NAND3x1_ASAP7_75t_SL g694 ( 
.A(n_670),
.B(n_664),
.C(n_646),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_667),
.Y(n_695)
);

OAI211xp5_ASAP7_75t_L g696 ( 
.A1(n_690),
.A2(n_631),
.B(n_659),
.C(n_653),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_667),
.Y(n_697)
);

NAND4xp75_ASAP7_75t_L g698 ( 
.A(n_676),
.B(n_663),
.C(n_655),
.D(n_646),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_671),
.B(n_632),
.C(n_643),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_685),
.B(n_652),
.C(n_657),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_683),
.B(n_660),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_686),
.B(n_658),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_683),
.B(n_654),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_692),
.B(n_648),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_673),
.B(n_687),
.C(n_691),
.Y(n_705)
);

OAI211xp5_ASAP7_75t_SL g706 ( 
.A1(n_669),
.A2(n_420),
.B(n_427),
.C(n_423),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_691),
.B(n_231),
.C(n_389),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_675),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_695),
.B(n_672),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_693),
.B(n_675),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_708),
.Y(n_711)
);

NAND4xp75_ASAP7_75t_L g712 ( 
.A(n_704),
.B(n_686),
.C(n_688),
.D(n_672),
.Y(n_712)
);

XNOR2xp5_ASAP7_75t_L g713 ( 
.A(n_705),
.B(n_694),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_697),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_701),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_703),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_702),
.B(n_681),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_714),
.Y(n_718)
);

XNOR2x1_ASAP7_75t_L g719 ( 
.A(n_713),
.B(n_698),
.Y(n_719)
);

XNOR2x1_ASAP7_75t_L g720 ( 
.A(n_712),
.B(n_699),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_715),
.A2(n_702),
.B1(n_700),
.B2(n_696),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_714),
.Y(n_722)
);

XNOR2x1_ASAP7_75t_L g723 ( 
.A(n_719),
.B(n_717),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_718),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_722),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_725),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_725),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_724),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_728),
.A2(n_721),
.B(n_715),
.C(n_723),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_729),
.A2(n_720),
.B1(n_715),
.B2(n_716),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_730),
.A2(n_727),
.B1(n_715),
.B2(n_716),
.Y(n_732)
);

AO22x2_ASAP7_75t_L g733 ( 
.A1(n_730),
.A2(n_717),
.B1(n_710),
.B2(n_707),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_731),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_732),
.Y(n_735)
);

AOI221xp5_ASAP7_75t_L g736 ( 
.A1(n_733),
.A2(n_696),
.B1(n_710),
.B2(n_711),
.C(n_674),
.Y(n_736)
);

AOI221xp5_ASAP7_75t_L g737 ( 
.A1(n_731),
.A2(n_710),
.B1(n_711),
.B2(n_668),
.C(n_709),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_731),
.A2(n_684),
.B1(n_706),
.B2(n_682),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_731),
.A2(n_678),
.B1(n_677),
.B2(n_679),
.Y(n_739)
);

AOI221xp5_ASAP7_75t_L g740 ( 
.A1(n_731),
.A2(n_689),
.B1(n_231),
.B2(n_82),
.C(n_83),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_739),
.B(n_77),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_734),
.A2(n_204),
.B1(n_203),
.B2(n_202),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_738),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_736),
.B(n_79),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_737),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_741),
.B(n_742),
.Y(n_747)
);

NAND4xp75_ASAP7_75t_L g748 ( 
.A(n_744),
.B(n_740),
.C(n_86),
.D(n_87),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_746),
.A2(n_204),
.B1(n_203),
.B2(n_202),
.Y(n_749)
);

OAI211xp5_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_204),
.B(n_203),
.C(n_91),
.Y(n_750)
);

NOR4xp25_ASAP7_75t_L g751 ( 
.A(n_743),
.B(n_85),
.C(n_88),
.D(n_92),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_747),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_749),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_748),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_751),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_750),
.B(n_98),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_747),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_747),
.B(n_99),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_747),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_759),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_757),
.A2(n_204),
.B1(n_203),
.B2(n_428),
.Y(n_761)
);

OA22x2_ASAP7_75t_L g762 ( 
.A1(n_752),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_762)
);

AO22x2_ASAP7_75t_L g763 ( 
.A1(n_755),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_763)
);

OAI22x1_ASAP7_75t_L g764 ( 
.A1(n_754),
.A2(n_204),
.B1(n_203),
.B2(n_112),
.Y(n_764)
);

AOI211xp5_ASAP7_75t_L g765 ( 
.A1(n_758),
.A2(n_110),
.B(n_111),
.C(n_115),
.Y(n_765)
);

OAI22x1_ASAP7_75t_L g766 ( 
.A1(n_753),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_756),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_760),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_763),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_767),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_762),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_766),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_768),
.A2(n_756),
.B1(n_764),
.B2(n_765),
.Y(n_773)
);

AO22x1_ASAP7_75t_L g774 ( 
.A1(n_769),
.A2(n_761),
.B1(n_127),
.B2(n_128),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_773),
.B(n_770),
.Y(n_775)
);

OA22x2_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_771),
.B1(n_772),
.B2(n_774),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_776),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_777),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.C(n_131),
.Y(n_778)
);

AOI211xp5_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_132),
.B(n_134),
.C(n_136),
.Y(n_779)
);


endmodule