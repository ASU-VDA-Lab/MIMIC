module fake_jpeg_27102_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVxp67_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx2_ASAP7_75t_SL g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_3),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_19),
.B1(n_22),
.B2(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.C(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_4),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_6),
.B1(n_10),
.B2(n_7),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_10),
.B1(n_7),
.B2(n_14),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_28),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_18),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_25),
.B1(n_33),
.B2(n_24),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_33),
.B1(n_37),
.B2(n_26),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_34),
.C(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI221xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_13),
.B1(n_42),
.B2(n_48),
.C(n_40),
.Y(n_50)
);


endmodule