module fake_netlist_6_4254_n_2999 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2999);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2999;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2510;
wire n_1954;
wire n_1735;
wire n_2044;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_405;
wire n_2660;
wire n_538;
wire n_2981;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_494;
wire n_539;
wire n_493;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_2714;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2749;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_835;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_2932;
wire n_595;
wire n_1767;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_417;
wire n_2857;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_623;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_811;
wire n_527;
wire n_1207;
wire n_683;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2357;
wire n_2025;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_2990;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_497;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_401;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_664;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_392;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_466;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2904;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_579;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_411;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_482;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_523;
wire n_707;
wire n_2986;
wire n_1900;
wire n_1548;
wire n_799;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_2834;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_414;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_393;
wire n_984;
wire n_2600;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_2899;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_18),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_244),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_370),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_286),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_201),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_6),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_192),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_7),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_26),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_6),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_155),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_303),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_77),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_190),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_44),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_386),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_169),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_216),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_291),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_42),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_302),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_213),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_351),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_128),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_177),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g421 ( 
.A(n_9),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_199),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_250),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_292),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_245),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_164),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_307),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_387),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_262),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_377),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_290),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_34),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_33),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_115),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_96),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_164),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_71),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_191),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_308),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_220),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_106),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_246),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_91),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_122),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_17),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_210),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_181),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_258),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_312),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_102),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_57),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_59),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_268),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_2),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_1),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_128),
.Y(n_461)
);

BUFx5_ASAP7_75t_L g462 ( 
.A(n_167),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_371),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_373),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_173),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_157),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_110),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_243),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_330),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_18),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_161),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_54),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_182),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_318),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_234),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_338),
.Y(n_476)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_241),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_322),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_67),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_41),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_127),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_339),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_255),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_112),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_73),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_257),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_13),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_360),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_211),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_199),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_357),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_169),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_40),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_7),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_55),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_313),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_113),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_375),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_310),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_192),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_305),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_103),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_190),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_48),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_229),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_260),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_270),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_368),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_125),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_343),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_382),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_232),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_158),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_84),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_297),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_16),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_28),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_389),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_300),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_218),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_224),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_149),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_76),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_89),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_222),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_58),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_70),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_84),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_81),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_273),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_271),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_127),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_71),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_205),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_4),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_321),
.Y(n_537)
);

BUFx8_ASAP7_75t_SL g538 ( 
.A(n_242),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_80),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_105),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_381),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_252),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_105),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_385),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_337),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_142),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_155),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_228),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_5),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_185),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_201),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_196),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_209),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_31),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_144),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_315),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_236),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_92),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_137),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_196),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_186),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_46),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_259),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_135),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_29),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_284),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_99),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_309),
.Y(n_568)
);

BUFx2_ASAP7_75t_SL g569 ( 
.A(n_277),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_227),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_326),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_295),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_346),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_341),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_323),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_361),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_266),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_30),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_43),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_175),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_33),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_274),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_200),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_5),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_153),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_233),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_152),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_251),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_122),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_391),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_8),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_121),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_21),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_366),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_109),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_294),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_64),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_353),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_363),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_157),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_193),
.Y(n_601)
);

INVxp33_ASAP7_75t_SL g602 ( 
.A(n_75),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_345),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_3),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_219),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_20),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_207),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_72),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_289),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_86),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_108),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_336),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_187),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_335),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_70),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_31),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_247),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_73),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_203),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_40),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_81),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_39),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_129),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_130),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_374),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_110),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_87),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_19),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_180),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_364),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_11),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_29),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_379),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_185),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_202),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_314),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_269),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_206),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_350),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_37),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_46),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_21),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_261),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_153),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_119),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_32),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_275),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_388),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_263),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_137),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_156),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_26),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_11),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_282),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_23),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_87),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_235),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_4),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_184),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_352),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_204),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_129),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_96),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_8),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_281),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_113),
.Y(n_666)
);

INVx4_ASAP7_75t_R g667 ( 
.A(n_53),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_288),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_141),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_47),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_22),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_16),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_280),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_176),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_166),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_93),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_151),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_240),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_170),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_367),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_1),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_249),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_100),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_187),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_134),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_150),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_369),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_93),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_193),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_114),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_47),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_24),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_163),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_34),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_184),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_145),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_38),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_145),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_474),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_521),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_541),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_421),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_393),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_421),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_506),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_421),
.Y(n_706)
);

CKINVDCx14_ASAP7_75t_R g707 ( 
.A(n_473),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_421),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_396),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_487),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_421),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_611),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_421),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_421),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_421),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_462),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_459),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_462),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_612),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_465),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_462),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_462),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_469),
.Y(n_723)
);

CKINVDCx16_ASAP7_75t_R g724 ( 
.A(n_661),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_466),
.Y(n_725)
);

INVxp33_ASAP7_75t_SL g726 ( 
.A(n_501),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_462),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_462),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_477),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_462),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_418),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_462),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_595),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_467),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_430),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_467),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_576),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_467),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_467),
.Y(n_739)
);

INVxp33_ASAP7_75t_SL g740 ( 
.A(n_644),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_467),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_552),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_536),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_481),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_536),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_536),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_454),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_536),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_536),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_483),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_392),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_552),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_552),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_454),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_593),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_593),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_500),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_593),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_487),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_540),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_540),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_670),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_581),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_670),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_484),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_485),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_581),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_454),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_601),
.Y(n_772)
);

CKINVDCx16_ASAP7_75t_R g773 ( 
.A(n_653),
.Y(n_773)
);

INVxp33_ASAP7_75t_SL g774 ( 
.A(n_392),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_601),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_601),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_601),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_601),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_645),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_645),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_645),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_645),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_491),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_645),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_495),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_398),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_399),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_498),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_496),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_496),
.Y(n_790)
);

INVxp33_ASAP7_75t_SL g791 ( 
.A(n_397),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_400),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_526),
.Y(n_793)
);

CKINVDCx14_ASAP7_75t_R g794 ( 
.A(n_653),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_504),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_504),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_614),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_653),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_564),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_564),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_591),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_521),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_591),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_503),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_407),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_586),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_669),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_586),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_419),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_680),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_598),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_422),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_432),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_434),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_505),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_669),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_438),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_439),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_598),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_672),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_448),
.Y(n_821)
);

INVxp33_ASAP7_75t_L g822 ( 
.A(n_445),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_672),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_689),
.Y(n_824)
);

INVxp33_ASAP7_75t_SL g825 ( 
.A(n_397),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_510),
.Y(n_826)
);

CKINVDCx16_ASAP7_75t_R g827 ( 
.A(n_404),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_447),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_689),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_451),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_456),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_460),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_461),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_470),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_472),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_479),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_494),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_401),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_734),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_734),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_723),
.B(n_519),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_736),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_701),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_726),
.A2(n_401),
.B1(n_409),
.B2(n_402),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_712),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_736),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_802),
.B(n_519),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_712),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_700),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_806),
.B(n_412),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_763),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_700),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_701),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_763),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_811),
.B(n_412),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_769),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_738),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_701),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_808),
.B(n_480),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_701),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_808),
.B(n_480),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_738),
.Y(n_863)
);

XOR2xp5_ASAP7_75t_L g864 ( 
.A(n_827),
.B(n_435),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_819),
.B(n_493),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_739),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_769),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_739),
.Y(n_868)
);

BUFx8_ASAP7_75t_SL g869 ( 
.A(n_703),
.Y(n_869)
);

BUFx8_ASAP7_75t_SL g870 ( 
.A(n_709),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_741),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_742),
.B(n_415),
.Y(n_873)
);

INVx6_ASAP7_75t_L g874 ( 
.A(n_819),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_743),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_743),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_699),
.B(n_602),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_745),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_745),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_746),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_715),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_746),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_748),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_748),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_707),
.Y(n_885)
);

CKINVDCx8_ASAP7_75t_R g886 ( 
.A(n_719),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_731),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_749),
.Y(n_889)
);

NOR2x1_ASAP7_75t_L g890 ( 
.A(n_749),
.B(n_569),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_765),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_821),
.B(n_415),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_768),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_705),
.B(n_416),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_770),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_772),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_724),
.B(n_538),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_729),
.B(n_416),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_742),
.B(n_431),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_737),
.B(n_431),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_759),
.B(n_488),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_775),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_760),
.B(n_493),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_776),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_710),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_721),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_777),
.Y(n_907)
);

CKINVDCx8_ASAP7_75t_R g908 ( 
.A(n_773),
.Y(n_908)
);

OA21x2_ASAP7_75t_L g909 ( 
.A1(n_711),
.A2(n_509),
.B(n_488),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_778),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_SL g911 ( 
.A1(n_726),
.A2(n_471),
.B1(n_524),
.B2(n_436),
.Y(n_911)
);

INVx6_ASAP7_75t_L g912 ( 
.A(n_798),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_779),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_761),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_780),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_721),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_762),
.B(n_509),
.Y(n_917)
);

AOI22x1_ASAP7_75t_SL g918 ( 
.A1(n_735),
.A2(n_589),
.B1(n_613),
.B2(n_585),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_789),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_764),
.B(n_635),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_781),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_717),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_789),
.Y(n_923)
);

OA21x2_ASAP7_75t_L g924 ( 
.A1(n_711),
.A2(n_638),
.B(n_635),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_782),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_784),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_752),
.B(n_638),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_753),
.B(n_395),
.Y(n_928)
);

OA21x2_ASAP7_75t_L g929 ( 
.A1(n_713),
.A2(n_408),
.B(n_403),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_790),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_790),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_702),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_803),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_755),
.B(n_425),
.Y(n_934)
);

OAI22x1_ASAP7_75t_R g935 ( 
.A1(n_750),
.A2(n_624),
.B1(n_652),
.B2(n_615),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_717),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_756),
.B(n_427),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_704),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_803),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_758),
.B(n_437),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_710),
.B(n_441),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_807),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_807),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_706),
.B(n_449),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_708),
.B(n_450),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_713),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_816),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_714),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_816),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_714),
.Y(n_950)
);

INVx6_ASAP7_75t_L g951 ( 
.A(n_813),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_716),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_716),
.B(n_458),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_718),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_718),
.B(n_463),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_720),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_722),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_722),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_727),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_727),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_728),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_728),
.B(n_541),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_730),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_869),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_922),
.B(n_720),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_870),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_952),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_888),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_905),
.B(n_877),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_888),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_885),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_952),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_963),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_886),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_963),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_885),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_932),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_886),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_932),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_938),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_874),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_R g982 ( 
.A(n_908),
.B(n_757),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_908),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_938),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_850),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_847),
.B(n_730),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_852),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_852),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_849),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_855),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_912),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_914),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_849),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_914),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_936),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_912),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_912),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_850),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_897),
.B(n_793),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_855),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_857),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_946),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_936),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_R g1004 ( 
.A(n_905),
.B(n_797),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_956),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_946),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_864),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_857),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_848),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_912),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_948),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_848),
.Y(n_1012)
);

NOR2xp67_ASAP7_75t_L g1013 ( 
.A(n_845),
.B(n_725),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_853),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_853),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_867),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_918),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_850),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_918),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_874),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_874),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_867),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_874),
.Y(n_1023)
);

NOR2xp67_ASAP7_75t_L g1024 ( 
.A(n_898),
.B(n_725),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_864),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_847),
.B(n_795),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_948),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_957),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_935),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_951),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_911),
.Y(n_1031)
);

AND3x2_ASAP7_75t_L g1032 ( 
.A(n_841),
.B(n_548),
.C(n_747),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_900),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_957),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_951),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_958),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_951),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_872),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_892),
.B(n_810),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_951),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_958),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_941),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_844),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_860),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_856),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_L g1046 ( 
.A(n_919),
.B(n_744),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_856),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_856),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_872),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_847),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_850),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_860),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_862),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_960),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_862),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_875),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_865),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_865),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_894),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_851),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_960),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_903),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_903),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_953),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_953),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_944),
.B(n_744),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_928),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_R g1068 ( 
.A(n_929),
.B(n_766),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_961),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_850),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_953),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_955),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_955),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_934),
.Y(n_1074)
);

NAND2xp33_ASAP7_75t_R g1075 ( 
.A(n_929),
.B(n_766),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_934),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_934),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_937),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_955),
.B(n_767),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_937),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_937),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_919),
.B(n_732),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_940),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_961),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_945),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_950),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_901),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_950),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_950),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_917),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_SL g1091 ( 
.A(n_927),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_927),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_920),
.B(n_774),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_875),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_884),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_927),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_962),
.B(n_767),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_873),
.B(n_899),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_R g1099 ( 
.A(n_929),
.B(n_783),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_950),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_919),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_890),
.B(n_783),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_931),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_931),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_884),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_854),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_931),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_950),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_873),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_873),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_929),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_942),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_909),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_942),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_899),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_899),
.B(n_785),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_942),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_895),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_942),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_895),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_930),
.B(n_795),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_942),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_962),
.B(n_785),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_854),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_909),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_943),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_896),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_896),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_954),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_854),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_904),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_904),
.B(n_774),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_954),
.B(n_732),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_907),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_987),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1098),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1098),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1052),
.B(n_794),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1052),
.B(n_788),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_1051),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1085),
.B(n_1087),
.Y(n_1141)
);

CKINVDCx6p67_ASAP7_75t_R g1142 ( 
.A(n_974),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1115),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_987),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_1025),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1112),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1059),
.B(n_791),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1092),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1053),
.B(n_788),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_988),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_988),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_990),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1121),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_1051),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_981),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1121),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1132),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1053),
.B(n_804),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_990),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1004),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1062),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_981),
.B(n_468),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1051),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1050),
.B(n_1059),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_994),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1030),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1055),
.B(n_804),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1090),
.B(n_954),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1051),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_989),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1055),
.B(n_815),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_967),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_972),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1051),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_964),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_973),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1000),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1070),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1026),
.B(n_475),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_975),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1000),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1044),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1104),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1026),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1045),
.Y(n_1186)
);

NOR2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1050),
.B(n_1035),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1060),
.B(n_954),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1070),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1001),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1047),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1063),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_982),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1048),
.Y(n_1194)
);

INVx5_ASAP7_75t_L g1195 ( 
.A(n_1070),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_SL g1196 ( 
.A(n_971),
.B(n_791),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1112),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1109),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1057),
.B(n_815),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1109),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1060),
.B(n_954),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_964),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_986),
.B(n_959),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1114),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1057),
.B(n_959),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1110),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1001),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1093),
.B(n_959),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1008),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1008),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1070),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1007),
.B(n_969),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1016),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1125),
.B(n_909),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_1070),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1106),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1125),
.B(n_959),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1058),
.B(n_959),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1106),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1111),
.A2(n_909),
.B1(n_924),
.B2(n_740),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1110),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1058),
.B(n_825),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1020),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1106),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1118),
.B(n_1127),
.C(n_1120),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1106),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1009),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_977),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1016),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_979),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_980),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_984),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1118),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1120),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1127),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1106),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1022),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1130),
.Y(n_1238)
);

AND2x6_ASAP7_75t_L g1239 ( 
.A(n_1114),
.B(n_541),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1021),
.Y(n_1240)
);

AND2x6_ASAP7_75t_L g1241 ( 
.A(n_1117),
.B(n_541),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1130),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1101),
.B(n_881),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1128),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1022),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1128),
.Y(n_1246)
);

NAND3x1_ASAP7_75t_L g1247 ( 
.A(n_1031),
.B(n_525),
.C(n_518),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1103),
.B(n_881),
.Y(n_1248)
);

NOR2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1037),
.B(n_826),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1131),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_966),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1038),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1064),
.B(n_541),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1064),
.B(n_633),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1131),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1134),
.B(n_825),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1134),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_968),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1023),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1038),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1113),
.A2(n_625),
.B1(n_648),
.B2(n_596),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1049),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1133),
.A2(n_924),
.B(n_887),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1049),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1096),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1056),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1107),
.B(n_1046),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1065),
.B(n_633),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_991),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1012),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1013),
.B(n_754),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1056),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1065),
.B(n_881),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1071),
.B(n_633),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1094),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1094),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1095),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_993),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1040),
.B(n_826),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1095),
.Y(n_1280)
);

CKINVDCx14_ASAP7_75t_R g1281 ( 
.A(n_999),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1116),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1130),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1071),
.B(n_476),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_SL g1285 ( 
.A(n_971),
.B(n_656),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1072),
.B(n_1073),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1024),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1033),
.Y(n_1288)
);

AND2x6_ASAP7_75t_L g1289 ( 
.A(n_1117),
.B(n_633),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_996),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1105),
.Y(n_1291)
);

AND2x2_ASAP7_75t_SL g1292 ( 
.A(n_1082),
.B(n_633),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1105),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1079),
.B(n_838),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_997),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1067),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1010),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1072),
.B(n_489),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1068),
.B(n_1099),
.C(n_1075),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1083),
.B(n_740),
.Y(n_1300)
);

AND3x1_ASAP7_75t_L g1301 ( 
.A(n_1043),
.B(n_751),
.C(n_733),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1002),
.Y(n_1302)
);

BUFx10_ASAP7_75t_L g1303 ( 
.A(n_976),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1073),
.B(n_502),
.Y(n_1304)
);

AND2x2_ASAP7_75t_SL g1305 ( 
.A(n_1119),
.B(n_639),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1130),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1006),
.B(n_1011),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_995),
.B(n_838),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1042),
.B(n_406),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_965),
.B(n_836),
.C(n_828),
.Y(n_1310)
);

OR2x6_ASAP7_75t_L g1311 ( 
.A(n_1102),
.B(n_771),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1066),
.B(n_822),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1027),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1014),
.B(n_671),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1130),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_985),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1028),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1034),
.B(n_887),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_985),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1036),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1003),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_985),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1097),
.B(n_639),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1119),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1015),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1041),
.B(n_887),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1054),
.B(n_906),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_998),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1074),
.B(n_507),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_978),
.B(n_517),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_SL g1331 ( 
.A(n_1303),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1136),
.B(n_1076),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1157),
.B(n_1005),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1137),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1299),
.A2(n_1078),
.B1(n_1080),
.B2(n_1077),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1135),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1141),
.B(n_1081),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1312),
.B(n_1169),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1208),
.B(n_1061),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_SL g1340 ( 
.A(n_1176),
.B(n_968),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1173),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1147),
.B(n_976),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1220),
.B(n_1069),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1220),
.B(n_1084),
.Y(n_1344)
);

AND2x4_ASAP7_75t_SL g1345 ( 
.A(n_1303),
.B(n_983),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1147),
.B(n_1039),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1135),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1256),
.B(n_1091),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1174),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1153),
.B(n_1086),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1177),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1225),
.B(n_1123),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1314),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1156),
.B(n_1088),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1233),
.A2(n_970),
.B1(n_516),
.B2(n_532),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1256),
.B(n_1091),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1314),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1193),
.Y(n_1358)
);

NAND2xp33_ASAP7_75t_L g1359 ( 
.A(n_1267),
.B(n_970),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1185),
.B(n_1122),
.Y(n_1360)
);

NAND2xp33_ASAP7_75t_L g1361 ( 
.A(n_1155),
.B(n_1122),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1292),
.A2(n_517),
.B1(n_554),
.B2(n_539),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1188),
.B(n_1089),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_SL g1364 ( 
.A(n_1223),
.B(n_639),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1292),
.A2(n_554),
.B1(n_677),
.B2(n_539),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1167),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1144),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1234),
.A2(n_544),
.B1(n_553),
.B2(n_508),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1301),
.A2(n_411),
.B1(n_414),
.B2(n_409),
.C(n_402),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1222),
.B(n_1165),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1180),
.A2(n_684),
.B1(n_677),
.B2(n_924),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1181),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1139),
.B(n_1032),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1262),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1264),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1188),
.B(n_1100),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1222),
.B(n_1091),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1180),
.A2(n_684),
.B1(n_924),
.B2(n_534),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1235),
.B(n_394),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1165),
.B(n_1108),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1201),
.B(n_1129),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1266),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1275),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1201),
.B(n_1261),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1243),
.B(n_1248),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1144),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1309),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1244),
.B(n_676),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1276),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1150),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1180),
.B(n_1126),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1307),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1252),
.A2(n_543),
.B1(n_555),
.B2(n_529),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1273),
.B(n_1126),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1217),
.B(n_998),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1203),
.A2(n_916),
.B(n_906),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1302),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1302),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1246),
.B(n_681),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1150),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1205),
.B(n_1124),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1205),
.B(n_1124),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1218),
.B(n_1320),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1151),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1151),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1313),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1313),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1317),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1152),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1152),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1317),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1218),
.B(n_1124),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1282),
.A2(n_1018),
.B1(n_998),
.B2(n_563),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1228),
.B(n_1230),
.Y(n_1414)
);

INVxp67_ASAP7_75t_SL g1415 ( 
.A(n_1155),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1252),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1231),
.B(n_1018),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1250),
.B(n_394),
.Y(n_1418)
);

NAND2xp33_ASAP7_75t_L g1419 ( 
.A(n_1155),
.B(n_1164),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1214),
.A2(n_571),
.B1(n_582),
.B2(n_557),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1155),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1260),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1255),
.B(n_405),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1257),
.B(n_685),
.Y(n_1424)
);

INVx4_ASAP7_75t_L g1425 ( 
.A(n_1167),
.Y(n_1425)
);

NOR2xp67_ASAP7_75t_L g1426 ( 
.A(n_1287),
.B(n_1017),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1260),
.A2(n_561),
.B1(n_567),
.B2(n_560),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1272),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1232),
.B(n_1214),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1272),
.Y(n_1430)
);

OAI22x1_ASAP7_75t_SL g1431 ( 
.A1(n_1145),
.A2(n_1029),
.B1(n_1019),
.B2(n_696),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1305),
.B(n_1018),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1160),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1305),
.B(n_1159),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1166),
.B(n_594),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1160),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1277),
.B(n_599),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1277),
.B(n_603),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1280),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_SL g1440 ( 
.A(n_1223),
.B(n_639),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1280),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1291),
.A2(n_580),
.B1(n_583),
.B2(n_578),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1291),
.B(n_605),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1293),
.B(n_609),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1293),
.B(n_619),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1178),
.B(n_654),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1178),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1182),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1182),
.B(n_657),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1171),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1164),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1190),
.B(n_660),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1281),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1263),
.A2(n_916),
.B(n_906),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1190),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1145),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1207),
.B(n_668),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1294),
.B(n_514),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1207),
.B(n_839),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1196),
.A2(n_410),
.B1(n_413),
.B2(n_405),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1209),
.B(n_839),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1253),
.A2(n_608),
.B(n_628),
.C(n_600),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1209),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1210),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1210),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1325),
.B(n_410),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1213),
.B(n_840),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1213),
.B(n_1229),
.Y(n_1468)
);

O2A1O1Ixp5_ASAP7_75t_L g1469 ( 
.A1(n_1323),
.A2(n_842),
.B(n_846),
.C(n_840),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1229),
.B(n_842),
.Y(n_1470)
);

INVx8_ASAP7_75t_L g1471 ( 
.A(n_1284),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1237),
.B(n_846),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1309),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1212),
.B(n_1183),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1149),
.B(n_1158),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1168),
.B(n_413),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1172),
.B(n_417),
.Y(n_1477)
);

INVxp33_ASAP7_75t_L g1478 ( 
.A(n_1308),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1198),
.A2(n_423),
.B1(n_424),
.B2(n_417),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1237),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1199),
.B(n_423),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1245),
.B(n_858),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1392),
.B(n_1279),
.Y(n_1483)
);

NOR3xp33_ASAP7_75t_L g1484 ( 
.A(n_1346),
.B(n_1300),
.C(n_1286),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1366),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1385),
.B(n_1200),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1451),
.A2(n_1154),
.B(n_1140),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1451),
.A2(n_1154),
.B(n_1140),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1353),
.B(n_1206),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1451),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1336),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1357),
.B(n_1338),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1341),
.Y(n_1493)
);

NOR2xp67_ASAP7_75t_L g1494 ( 
.A(n_1453),
.B(n_1310),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1451),
.A2(n_1154),
.B(n_1140),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1419),
.A2(n_1175),
.B(n_1170),
.Y(n_1496)
);

BUFx8_ASAP7_75t_L g1497 ( 
.A(n_1331),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1349),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1333),
.B(n_1300),
.C(n_1285),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1387),
.B(n_1473),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1336),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1370),
.A2(n_1221),
.B(n_1298),
.C(n_1284),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1370),
.B(n_1240),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1450),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1351),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_L g1506 ( 
.A(n_1425),
.B(n_1240),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1372),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1454),
.A2(n_1175),
.B(n_1170),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1366),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1384),
.B(n_1337),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1339),
.A2(n_1175),
.B(n_1170),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1337),
.B(n_1148),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1395),
.A2(n_1211),
.B(n_1189),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1342),
.B(n_1161),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1380),
.B(n_1143),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1333),
.B(n_1321),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1458),
.B(n_1227),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1429),
.A2(n_1211),
.B(n_1189),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1343),
.A2(n_1245),
.B(n_1323),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1474),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1391),
.A2(n_1211),
.B(n_1189),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1380),
.B(n_1259),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1416),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1425),
.B(n_1259),
.Y(n_1524)
);

OAI321xp33_ASAP7_75t_L g1525 ( 
.A1(n_1369),
.A2(n_1311),
.A3(n_1271),
.B1(n_1253),
.B2(n_1274),
.C(n_1268),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1471),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1471),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1362),
.A2(n_1298),
.B(n_1304),
.C(n_1284),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1347),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1334),
.B(n_1298),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1475),
.B(n_1162),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1403),
.B(n_1186),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1347),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1421),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1394),
.A2(n_1315),
.B(n_1236),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1422),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1377),
.B(n_1191),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1458),
.B(n_1304),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1332),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1344),
.A2(n_1268),
.B(n_1254),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1414),
.B(n_1304),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1342),
.B(n_1281),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1362),
.B(n_1254),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1361),
.A2(n_1315),
.B(n_1236),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1426),
.B(n_1184),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1421),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1474),
.B(n_1388),
.Y(n_1547)
);

AOI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1401),
.A2(n_1274),
.B(n_1318),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1365),
.B(n_1278),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1415),
.A2(n_1315),
.B(n_1236),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1402),
.A2(n_1215),
.B(n_1195),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1428),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1430),
.Y(n_1553)
);

AO21x1_ASAP7_75t_L g1554 ( 
.A1(n_1420),
.A2(n_1327),
.B(n_1326),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1377),
.B(n_1348),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1386),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1412),
.A2(n_1215),
.B(n_1195),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1388),
.B(n_1399),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1332),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1386),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1335),
.B(n_1187),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1468),
.A2(n_1215),
.B(n_1195),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1363),
.A2(n_1381),
.B(n_1376),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1434),
.A2(n_1194),
.B1(n_1286),
.B2(n_1319),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1365),
.B(n_1329),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1456),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1432),
.A2(n_1197),
.B(n_1146),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1399),
.B(n_1184),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1378),
.A2(n_1215),
.B(n_1195),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1368),
.A2(n_1311),
.B(n_1271),
.C(n_1329),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1547),
.B(n_1348),
.Y(n_1571)
);

AND2x4_ASAP7_75t_SL g1572 ( 
.A(n_1526),
.B(n_1303),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1558),
.B(n_1424),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1485),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1508),
.A2(n_1396),
.B(n_1197),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1547),
.A2(n_1397),
.B1(n_1406),
.B2(n_1398),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1493),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1513),
.A2(n_1521),
.B(n_1518),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1496),
.A2(n_1179),
.B(n_1164),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1510),
.A2(n_1356),
.B(n_1424),
.C(n_1352),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_SL g1581 ( 
.A1(n_1484),
.A2(n_1356),
.B(n_1440),
.C(n_1364),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1498),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1514),
.B(n_1478),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1485),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1538),
.A2(n_1355),
.B(n_1477),
.C(n_1476),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1510),
.A2(n_1469),
.B(n_1354),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1486),
.B(n_1471),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1544),
.A2(n_1179),
.B(n_1164),
.Y(n_1588)
);

AOI22x1_ASAP7_75t_L g1589 ( 
.A1(n_1540),
.A2(n_1408),
.B1(n_1411),
.B2(n_1407),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1566),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1522),
.A2(n_1378),
.B1(n_1371),
.B2(n_1413),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1511),
.A2(n_1216),
.B(n_1179),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1505),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1559),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1490),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1514),
.A2(n_1481),
.B(n_1418),
.C(n_1423),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1534),
.Y(n_1597)
);

NAND2x1p5_ASAP7_75t_L g1598 ( 
.A(n_1526),
.B(n_1439),
.Y(n_1598)
);

BUFx8_ASAP7_75t_SL g1599 ( 
.A(n_1561),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1502),
.A2(n_1359),
.B(n_1435),
.C(n_1379),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1535),
.A2(n_1216),
.B(n_1179),
.Y(n_1601)
);

INVx6_ASAP7_75t_L g1602 ( 
.A(n_1526),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1502),
.A2(n_1350),
.B(n_1373),
.C(n_1329),
.Y(n_1603)
);

AO22x1_ASAP7_75t_L g1604 ( 
.A1(n_1542),
.A2(n_1258),
.B1(n_1176),
.B2(n_1202),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_SL g1605 ( 
.A(n_1499),
.B(n_1258),
.C(n_1340),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1515),
.B(n_1265),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1541),
.A2(n_1371),
.B1(n_1375),
.B2(n_1374),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1525),
.A2(n_1383),
.B(n_1389),
.C(n_1382),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1503),
.A2(n_1270),
.B1(n_1417),
.B2(n_1311),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1556),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1483),
.B(n_1393),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1569),
.A2(n_1219),
.B(n_1216),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1542),
.B(n_1345),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1520),
.B(n_1296),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1526),
.B(n_1269),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1519),
.A2(n_1219),
.B(n_1216),
.Y(n_1616)
);

OAI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1512),
.A2(n_1543),
.B1(n_1565),
.B2(n_1492),
.Y(n_1617)
);

NOR3xp33_ASAP7_75t_SL g1618 ( 
.A(n_1555),
.B(n_1358),
.C(n_1460),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1503),
.B(n_1441),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1550),
.A2(n_1224),
.B(n_1219),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1555),
.A2(n_1271),
.B(n_1466),
.C(n_1462),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1537),
.A2(n_1479),
.B(n_1330),
.C(n_1288),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1507),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1516),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1610),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1575),
.A2(n_1548),
.B(n_1567),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1571),
.B(n_1564),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_SL g1628 ( 
.A(n_1580),
.B(n_1570),
.C(n_1517),
.Y(n_1628)
);

O2A1O1Ixp5_ASAP7_75t_L g1629 ( 
.A1(n_1581),
.A2(n_1537),
.B(n_1554),
.C(n_1568),
.Y(n_1629)
);

INVx8_ASAP7_75t_L g1630 ( 
.A(n_1595),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1615),
.B(n_1527),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1578),
.A2(n_1557),
.B(n_1551),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1577),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1603),
.A2(n_1528),
.B(n_1568),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1582),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1593),
.Y(n_1636)
);

NAND3x1_ASAP7_75t_L g1637 ( 
.A(n_1583),
.B(n_1545),
.C(n_1524),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1623),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1601),
.A2(n_1563),
.B(n_1562),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1606),
.B(n_1500),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1600),
.A2(n_1528),
.B(n_1532),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1592),
.A2(n_1488),
.B(n_1487),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1597),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1576),
.B(n_1523),
.Y(n_1644)
);

AO31x2_ASAP7_75t_L g1645 ( 
.A1(n_1616),
.A2(n_1438),
.A3(n_1443),
.B(n_1437),
.Y(n_1645)
);

AOI221x1_ASAP7_75t_L g1646 ( 
.A1(n_1609),
.A2(n_1500),
.B1(n_1549),
.B2(n_1561),
.C(n_1489),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1589),
.A2(n_1495),
.B(n_1445),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1619),
.A2(n_1446),
.B(n_1444),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1588),
.A2(n_1452),
.B(n_1449),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1579),
.A2(n_1457),
.B(n_1459),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1605),
.B(n_1504),
.Y(n_1651)
);

AOI221x1_ASAP7_75t_L g1652 ( 
.A1(n_1608),
.A2(n_1552),
.B1(n_1553),
.B2(n_1536),
.C(n_1530),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1585),
.A2(n_1532),
.B(n_1506),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1617),
.A2(n_1531),
.B(n_1467),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1583),
.A2(n_1192),
.B1(n_1494),
.B2(n_1138),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1617),
.B(n_1559),
.Y(n_1656)
);

AOI221x1_ASAP7_75t_L g1657 ( 
.A1(n_1586),
.A2(n_641),
.B1(n_655),
.B2(n_632),
.C(n_629),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1595),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1597),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1612),
.A2(n_1470),
.B(n_1461),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1581),
.A2(n_1591),
.B(n_1620),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1614),
.B(n_1202),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1619),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1587),
.A2(n_1490),
.B(n_1224),
.Y(n_1664)
);

AOI31xp67_ASAP7_75t_L g1665 ( 
.A1(n_1611),
.A2(n_1560),
.A3(n_1556),
.B(n_1501),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1576),
.B(n_1618),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1598),
.A2(n_1482),
.B(n_1472),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1594),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1598),
.A2(n_1560),
.B(n_1400),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1621),
.A2(n_1400),
.B(n_1390),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1596),
.A2(n_1247),
.B(n_1163),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_SL g1672 ( 
.A1(n_1607),
.A2(n_1622),
.B(n_1546),
.C(n_1534),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1614),
.B(n_1539),
.Y(n_1673)
);

INVx3_ASAP7_75t_SL g1674 ( 
.A(n_1630),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1665),
.Y(n_1675)
);

AO21x2_ASAP7_75t_L g1676 ( 
.A1(n_1661),
.A2(n_1618),
.B(n_1464),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1663),
.B(n_1666),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1665),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1633),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1640),
.A2(n_1613),
.B1(n_1615),
.B2(n_1331),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1657),
.A2(n_1480),
.B(n_1447),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1642),
.A2(n_1404),
.B(n_1390),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1624),
.B(n_1613),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1662),
.A2(n_1615),
.B1(n_1574),
.B2(n_1345),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1625),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1643),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1642),
.A2(n_1405),
.B(n_1404),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1639),
.A2(n_1410),
.B(n_1405),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1625),
.Y(n_1689)
);

BUFx10_ASAP7_75t_L g1690 ( 
.A(n_1631),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1634),
.B(n_1604),
.C(n_1427),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1639),
.A2(n_1433),
.B(n_1410),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1659),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1628),
.A2(n_1590),
.B1(n_1599),
.B2(n_1269),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1635),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1666),
.A2(n_1290),
.B1(n_1297),
.B2(n_1295),
.Y(n_1697)
);

AO21x2_ASAP7_75t_L g1698 ( 
.A1(n_1632),
.A2(n_1546),
.B(n_1529),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1629),
.A2(n_1247),
.B(n_1163),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1630),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1636),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1632),
.A2(n_1436),
.B(n_1433),
.Y(n_1702)
);

CKINVDCx6p67_ASAP7_75t_R g1703 ( 
.A(n_1631),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1644),
.B(n_1491),
.Y(n_1704)
);

NAND2x1_ASAP7_75t_L g1705 ( 
.A(n_1641),
.B(n_1490),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1647),
.A2(n_1448),
.B(n_1436),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1657),
.A2(n_913),
.B(n_907),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1673),
.B(n_1142),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1638),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1670),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1670),
.Y(n_1713)
);

AO21x2_ASAP7_75t_L g1714 ( 
.A1(n_1626),
.A2(n_1533),
.B(n_1163),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1668),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1647),
.A2(n_1455),
.B(n_1448),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1656),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1671),
.A2(n_1295),
.B1(n_1297),
.B2(n_1290),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1626),
.A2(n_1463),
.B(n_1455),
.Y(n_1719)
);

AO21x1_ASAP7_75t_L g1720 ( 
.A1(n_1627),
.A2(n_690),
.B(n_663),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1649),
.A2(n_1465),
.B(n_1463),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1645),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1653),
.A2(n_1572),
.B(n_1393),
.C(n_1442),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1627),
.A2(n_1490),
.B(n_1224),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1658),
.B(n_1527),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1644),
.B(n_639),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1655),
.B(n_1142),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1649),
.A2(n_1465),
.B(n_1197),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1651),
.A2(n_1330),
.B1(n_1249),
.B2(n_1497),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1658),
.B(n_1527),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1646),
.B(n_1654),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1664),
.B(n_1251),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1630),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1637),
.A2(n_1667),
.B(n_1660),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1650),
.A2(n_1204),
.B(n_1146),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1672),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1650),
.A2(n_1204),
.B(n_1146),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1645),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1630),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1637),
.B(n_1584),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1652),
.A2(n_1672),
.B(n_1667),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1645),
.B(n_647),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1648),
.A2(n_691),
.B(n_695),
.C(n_694),
.Y(n_1743)
);

OAI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1660),
.A2(n_1324),
.B(n_1204),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1648),
.A2(n_1442),
.B(n_1427),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1658),
.B(n_1527),
.Y(n_1746)
);

AO31x2_ASAP7_75t_L g1747 ( 
.A1(n_1645),
.A2(n_1409),
.A3(n_1367),
.B(n_1322),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1669),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1669),
.A2(n_1324),
.B(n_1316),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1645),
.A2(n_1324),
.B(n_1316),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1630),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_1659),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1634),
.A2(n_1224),
.B(n_1219),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1656),
.B(n_1509),
.Y(n_1754)
);

OAI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1642),
.A2(n_893),
.B(n_891),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1634),
.A2(n_428),
.B(n_429),
.C(n_424),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1663),
.Y(n_1757)
);

O2A1O1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1628),
.A2(n_1330),
.B(n_786),
.C(n_792),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1643),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1715),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1677),
.B(n_515),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1715),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1677),
.B(n_523),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1679),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1752),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1757),
.B(n_647),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1679),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1757),
.B(n_647),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1701),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1717),
.B(n_527),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1723),
.A2(n_1322),
.B(n_1319),
.Y(n_1771)
);

AO21x2_ASAP7_75t_L g1772 ( 
.A1(n_1741),
.A2(n_831),
.B(n_830),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1701),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1711),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1711),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1752),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1692),
.B(n_1251),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1740),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1731),
.A2(n_1322),
.B(n_1319),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1757),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1696),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1755),
.A2(n_925),
.B(n_913),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1691),
.Y(n_1783)
);

AO21x2_ASAP7_75t_L g1784 ( 
.A1(n_1734),
.A2(n_831),
.B(n_830),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1685),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1694),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1748),
.B(n_930),
.Y(n_1787)
);

OAI21x1_ASAP7_75t_SL g1788 ( 
.A1(n_1720),
.A2(n_832),
.B(n_805),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1703),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1703),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1686),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1717),
.B(n_1759),
.Y(n_1792)
);

BUFx4f_ASAP7_75t_SL g1793 ( 
.A(n_1674),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1685),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1742),
.B(n_647),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1756),
.A2(n_1743),
.B(n_1758),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1754),
.B(n_1704),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1689),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1689),
.Y(n_1799)
);

OAI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1755),
.A2(n_926),
.B(n_925),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1736),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1742),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1748),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1754),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1726),
.B(n_647),
.Y(n_1806)
);

AO21x2_ASAP7_75t_L g1807 ( 
.A1(n_1678),
.A2(n_832),
.B(n_809),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1675),
.Y(n_1808)
);

OAI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1735),
.A2(n_926),
.B(n_893),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1708),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1753),
.A2(n_1328),
.B(n_1242),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1704),
.B(n_528),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1738),
.Y(n_1813)
);

AOI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1732),
.A2(n_812),
.B(n_787),
.Y(n_1814)
);

OA21x2_ASAP7_75t_L g1815 ( 
.A1(n_1678),
.A2(n_799),
.B(n_796),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1726),
.Y(n_1816)
);

NAND2x1p5_ASAP7_75t_L g1817 ( 
.A(n_1705),
.B(n_1238),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1675),
.Y(n_1818)
);

OAI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1680),
.A2(n_414),
.B1(n_420),
.B2(n_411),
.Y(n_1819)
);

OAI21x1_ASAP7_75t_L g1820 ( 
.A1(n_1735),
.A2(n_902),
.B(n_891),
.Y(n_1820)
);

AO21x2_ASAP7_75t_L g1821 ( 
.A1(n_1712),
.A2(n_1750),
.B(n_1713),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_SL g1822 ( 
.A1(n_1727),
.A2(n_1497),
.B1(n_426),
.B2(n_440),
.Y(n_1822)
);

AO21x1_ASAP7_75t_L g1823 ( 
.A1(n_1699),
.A2(n_817),
.B(n_814),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1722),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1695),
.A2(n_833),
.B(n_818),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1722),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1690),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1683),
.B(n_530),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1712),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1713),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1676),
.B(n_533),
.Y(n_1831)
);

OA21x2_ASAP7_75t_L g1832 ( 
.A1(n_1750),
.A2(n_799),
.B(n_796),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1747),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1676),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1698),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1747),
.B(n_834),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1745),
.A2(n_1328),
.B(n_1242),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1698),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1724),
.A2(n_1328),
.B(n_1242),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1747),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1690),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1720),
.B(n_1251),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1747),
.B(n_800),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1676),
.B(n_546),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1674),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1747),
.B(n_800),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1737),
.A2(n_1744),
.B(n_1728),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1698),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1719),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1719),
.Y(n_1850)
);

AO21x1_ASAP7_75t_L g1851 ( 
.A1(n_1705),
.A2(n_837),
.B(n_835),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1681),
.A2(n_1242),
.B(n_1238),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1681),
.A2(n_1283),
.B(n_1238),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1681),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1718),
.A2(n_1602),
.B1(n_426),
.B2(n_440),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1714),
.B(n_801),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1706),
.Y(n_1857)
);

OA21x2_ASAP7_75t_L g1858 ( 
.A1(n_1737),
.A2(n_820),
.B(n_801),
.Y(n_1858)
);

AO21x2_ASAP7_75t_L g1859 ( 
.A1(n_1744),
.A2(n_823),
.B(n_820),
.Y(n_1859)
);

NAND2x1p5_ASAP7_75t_L g1860 ( 
.A(n_1708),
.B(n_1238),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1707),
.A2(n_1306),
.B(n_1283),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1708),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1710),
.B(n_547),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_1688),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1739),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1728),
.A2(n_902),
.B(n_863),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1714),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1709),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1684),
.A2(n_428),
.B(n_433),
.C(n_429),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1690),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1714),
.B(n_823),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1709),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1697),
.A2(n_1729),
.B(n_1707),
.Y(n_1873)
);

OAI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1707),
.A2(n_478),
.B(n_464),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1688),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1709),
.A2(n_1306),
.B(n_1283),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1721),
.B(n_824),
.Y(n_1877)
);

OAI21x1_ASAP7_75t_L g1878 ( 
.A1(n_1706),
.A2(n_863),
.B(n_858),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1716),
.A2(n_871),
.B(n_866),
.Y(n_1879)
);

CKINVDCx14_ASAP7_75t_R g1880 ( 
.A(n_1739),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1733),
.Y(n_1881)
);

AO21x2_ASAP7_75t_L g1882 ( 
.A1(n_1749),
.A2(n_829),
.B(n_824),
.Y(n_1882)
);

OAI21x1_ASAP7_75t_L g1883 ( 
.A1(n_1716),
.A2(n_871),
.B(n_866),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1725),
.A2(n_443),
.B1(n_446),
.B2(n_420),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1693),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1693),
.Y(n_1886)
);

BUFx2_ASAP7_75t_L g1887 ( 
.A(n_1733),
.Y(n_1887)
);

INVx5_ASAP7_75t_L g1888 ( 
.A(n_1725),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1682),
.Y(n_1889)
);

NOR2xp67_ASAP7_75t_L g1890 ( 
.A(n_1700),
.B(n_829),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1721),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1682),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1687),
.Y(n_1893)
);

OAI21x1_ASAP7_75t_L g1894 ( 
.A1(n_1749),
.A2(n_878),
.B(n_876),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1725),
.B(n_549),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1687),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1702),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1702),
.Y(n_1898)
);

AOI222xp33_ASAP7_75t_L g1899 ( 
.A1(n_1730),
.A2(n_620),
.B1(n_446),
.B2(n_621),
.C1(n_455),
.C2(n_443),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1700),
.A2(n_878),
.B(n_876),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1730),
.A2(n_1306),
.B(n_1283),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1730),
.A2(n_939),
.B(n_933),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1746),
.B(n_0),
.Y(n_1903)
);

OA21x2_ASAP7_75t_L g1904 ( 
.A1(n_1746),
.A2(n_939),
.B(n_933),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1751),
.B(n_1306),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1746),
.B(n_550),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1751),
.B(n_949),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1679),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1679),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1679),
.Y(n_1910)
);

AO21x2_ASAP7_75t_L g1911 ( 
.A1(n_1741),
.A2(n_880),
.B(n_879),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1764),
.Y(n_1912)
);

AO21x2_ASAP7_75t_L g1913 ( 
.A1(n_1848),
.A2(n_880),
.B(n_879),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1767),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1780),
.B(n_0),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1780),
.B(n_2),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1769),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1830),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1773),
.Y(n_1919)
);

AOI21x1_ASAP7_75t_L g1920 ( 
.A1(n_1777),
.A2(n_883),
.B(n_949),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1774),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1775),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1827),
.B(n_1602),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1830),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1908),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1802),
.B(n_3),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1909),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1829),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1910),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1845),
.Y(n_1930)
);

OA21x2_ASAP7_75t_L g1931 ( 
.A1(n_1852),
.A2(n_1853),
.B(n_1838),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1805),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1804),
.B(n_9),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1803),
.B(n_10),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1827),
.B(n_1602),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1813),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1781),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1808),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1845),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1791),
.Y(n_1940)
);

AO21x2_ASAP7_75t_L g1941 ( 
.A1(n_1867),
.A2(n_883),
.B(n_667),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1792),
.Y(n_1942)
);

INVx2_ASAP7_75t_SL g1943 ( 
.A(n_1765),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1803),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1783),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1808),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1818),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1762),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1881),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_SL g1950 ( 
.A1(n_1823),
.A2(n_10),
.B(n_12),
.Y(n_1950)
);

AOI21x1_ASAP7_75t_L g1951 ( 
.A1(n_1777),
.A2(n_620),
.B(n_455),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1818),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1776),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1785),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1881),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1785),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1794),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1794),
.Y(n_1958)
);

AO21x2_ASAP7_75t_L g1959 ( 
.A1(n_1807),
.A2(n_1360),
.B(n_12),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1765),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1803),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1798),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1798),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1793),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1799),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1799),
.Y(n_1966)
);

OA21x2_ASAP7_75t_L g1967 ( 
.A1(n_1835),
.A2(n_442),
.B(n_433),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1790),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1786),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_L g1970 ( 
.A(n_1869),
.B(n_621),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1834),
.B(n_13),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1797),
.B(n_551),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1824),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1826),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1778),
.B(n_558),
.Y(n_1975)
);

OA21x2_ASAP7_75t_L g1976 ( 
.A1(n_1835),
.A2(n_444),
.B(n_442),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1801),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1816),
.B(n_559),
.Y(n_1978)
);

AO21x1_ASAP7_75t_SL g1979 ( 
.A1(n_1831),
.A2(n_1431),
.B(n_14),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1863),
.B(n_562),
.Y(n_1980)
);

OA21x2_ASAP7_75t_L g1981 ( 
.A1(n_1838),
.A2(n_452),
.B(n_444),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1862),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1826),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1868),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1821),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1821),
.Y(n_1986)
);

BUFx3_ASAP7_75t_L g1987 ( 
.A(n_1865),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1846),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1821),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1846),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1847),
.A2(n_843),
.B(n_916),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1836),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1857),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1836),
.Y(n_1994)
);

BUFx2_ASAP7_75t_L g1995 ( 
.A(n_1841),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1841),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1810),
.Y(n_1997)
);

OR2x2_ASAP7_75t_SL g1998 ( 
.A(n_1844),
.B(n_14),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1857),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1886),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1843),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1854),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1833),
.B(n_1840),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1886),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1856),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1888),
.B(n_15),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1787),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1872),
.B(n_15),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1856),
.Y(n_2009)
);

AO21x2_ASAP7_75t_L g2010 ( 
.A1(n_1807),
.A2(n_1360),
.B(n_17),
.Y(n_2010)
);

INVx3_ASAP7_75t_L g2011 ( 
.A(n_1787),
.Y(n_2011)
);

BUFx4f_ASAP7_75t_SL g2012 ( 
.A(n_1762),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1795),
.B(n_19),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1787),
.Y(n_2014)
);

BUFx5_ASAP7_75t_L g2015 ( 
.A(n_1849),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1850),
.B(n_20),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1795),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1841),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1888),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1891),
.B(n_22),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1898),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1766),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1865),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1766),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1847),
.A2(n_843),
.B(n_1360),
.Y(n_2025)
);

OAI21x1_ASAP7_75t_L g2026 ( 
.A1(n_1820),
.A2(n_1861),
.B(n_1809),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1898),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1889),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1871),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1889),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1871),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1768),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1768),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1893),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1877),
.Y(n_2035)
);

OAI21x1_ASAP7_75t_L g2036 ( 
.A1(n_1820),
.A2(n_843),
.B(n_1360),
.Y(n_2036)
);

AO31x2_ASAP7_75t_L g2037 ( 
.A1(n_1823),
.A2(n_25),
.A3(n_23),
.B(n_24),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1761),
.B(n_565),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1789),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1809),
.A2(n_1360),
.B(n_212),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1763),
.B(n_579),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1789),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1893),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1896),
.Y(n_2044)
);

BUFx3_ASAP7_75t_L g2045 ( 
.A(n_1887),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1870),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1870),
.B(n_25),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1870),
.Y(n_2048)
);

OAI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1811),
.A2(n_214),
.B(n_208),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_1875),
.B(n_27),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1888),
.B(n_27),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1888),
.B(n_28),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1888),
.B(n_30),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1885),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1897),
.B(n_32),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1789),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1892),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1903),
.B(n_35),
.Y(n_2058)
);

BUFx2_ASAP7_75t_SL g2059 ( 
.A(n_1760),
.Y(n_2059)
);

AOI222xp33_ASAP7_75t_L g2060 ( 
.A1(n_1970),
.A2(n_1884),
.B1(n_1796),
.B2(n_1825),
.C1(n_1873),
.C2(n_1819),
.Y(n_2060)
);

INVx3_ASAP7_75t_L g2061 ( 
.A(n_1930),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1914),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1914),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1970),
.A2(n_1822),
.B1(n_1842),
.B2(n_1874),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_2056),
.B(n_1903),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_SL g2066 ( 
.A1(n_1998),
.A2(n_1880),
.B1(n_1884),
.B2(n_1828),
.Y(n_2066)
);

BUFx2_ASAP7_75t_L g2067 ( 
.A(n_2045),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1953),
.B(n_1806),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1991),
.A2(n_1896),
.B(n_1779),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1956),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1982),
.B(n_1911),
.Y(n_2071)
);

BUFx3_ASAP7_75t_L g2072 ( 
.A(n_1987),
.Y(n_2072)
);

INVx6_ASAP7_75t_SL g2073 ( 
.A(n_2006),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1956),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_1984),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1917),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1997),
.B(n_1911),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1979),
.A2(n_1842),
.B1(n_1851),
.B2(n_1788),
.Y(n_2078)
);

OAI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2012),
.A2(n_1814),
.B1(n_1770),
.B2(n_1890),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1958),
.Y(n_2080)
);

OAI22xp33_ASAP7_75t_SL g2081 ( 
.A1(n_1971),
.A2(n_2050),
.B1(n_2055),
.B2(n_2016),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_SL g2082 ( 
.A(n_2059),
.B(n_1772),
.Y(n_2082)
);

OAI21xp33_ASAP7_75t_L g2083 ( 
.A1(n_1992),
.A2(n_1899),
.B(n_1869),
.Y(n_2083)
);

AND2x4_ASAP7_75t_SL g2084 ( 
.A(n_2006),
.B(n_1806),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1998),
.A2(n_2059),
.B1(n_1976),
.B2(n_1981),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_1979),
.A2(n_1851),
.B1(n_1906),
.B2(n_1895),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_SL g2087 ( 
.A1(n_1967),
.A2(n_1880),
.B1(n_1772),
.B2(n_1812),
.Y(n_2087)
);

OAI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_1967),
.A2(n_1817),
.B1(n_1904),
.B2(n_1902),
.Y(n_2088)
);

OAI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_1980),
.A2(n_626),
.B1(n_627),
.B2(n_623),
.C(n_622),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_2019),
.B(n_1876),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2045),
.B(n_1784),
.Y(n_2091)
);

NAND4xp25_ASAP7_75t_L g2092 ( 
.A(n_2041),
.B(n_2038),
.C(n_1972),
.D(n_1975),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1987),
.Y(n_2093)
);

OA21x2_ASAP7_75t_L g2094 ( 
.A1(n_2002),
.A2(n_1864),
.B(n_1878),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_1960),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1930),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_SL g2097 ( 
.A1(n_1967),
.A2(n_1772),
.B1(n_1855),
.B2(n_1784),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1942),
.B(n_1911),
.Y(n_2098)
);

AOI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_1950),
.A2(n_1784),
.B1(n_1907),
.B2(n_1837),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1964),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1968),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1968),
.B(n_1817),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1943),
.B(n_1807),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1958),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_1967),
.A2(n_1902),
.B1(n_1904),
.B2(n_1905),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_SL g2106 ( 
.A1(n_1976),
.A2(n_1902),
.B1(n_1904),
.B2(n_1905),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_1950),
.A2(n_1907),
.B1(n_1771),
.B2(n_623),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1917),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1919),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1930),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2048),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2005),
.B(n_1882),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_2006),
.A2(n_626),
.B1(n_627),
.B2(n_622),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2005),
.B(n_1882),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1919),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2017),
.B(n_1882),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1943),
.B(n_1860),
.Y(n_2117)
);

OAI22xp33_ASAP7_75t_L g2118 ( 
.A1(n_1951),
.A2(n_1860),
.B1(n_1901),
.B2(n_1839),
.Y(n_2118)
);

OAI221xp5_ASAP7_75t_L g2119 ( 
.A1(n_1951),
.A2(n_640),
.B1(n_642),
.B2(n_634),
.C(n_631),
.Y(n_2119)
);

OAI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_1930),
.A2(n_634),
.B1(n_640),
.B2(n_631),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1976),
.A2(n_646),
.B1(n_650),
.B2(n_642),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_1939),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_2023),
.Y(n_2123)
);

INVx3_ASAP7_75t_L g2124 ( 
.A(n_1930),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1921),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_1994),
.A2(n_650),
.B1(n_651),
.B2(n_646),
.Y(n_2126)
);

OR2x6_ASAP7_75t_L g2127 ( 
.A(n_2019),
.B(n_1900),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1939),
.B(n_1859),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_SL g2129 ( 
.A1(n_1976),
.A2(n_658),
.B1(n_659),
.B2(n_651),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2056),
.B(n_1900),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1995),
.B(n_1859),
.Y(n_2131)
);

INVxp67_ASAP7_75t_L g2132 ( 
.A(n_1969),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_2023),
.Y(n_2133)
);

OAI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_1978),
.A2(n_662),
.B1(n_664),
.B2(n_659),
.C(n_658),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_1981),
.A2(n_1859),
.B(n_1832),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2035),
.B(n_1832),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1966),
.Y(n_2137)
);

AOI211xp5_ASAP7_75t_L g2138 ( 
.A1(n_2051),
.A2(n_664),
.B(n_666),
.C(n_662),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_1988),
.A2(n_674),
.B1(n_675),
.B2(n_666),
.Y(n_2139)
);

OAI21x1_ASAP7_75t_L g2140 ( 
.A1(n_1991),
.A2(n_1866),
.B(n_1815),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_1990),
.A2(n_675),
.B1(n_679),
.B2(n_674),
.Y(n_2141)
);

OAI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_1971),
.A2(n_686),
.B1(n_688),
.B2(n_683),
.C(n_679),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_1981),
.A2(n_1832),
.B(n_1858),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_2001),
.A2(n_686),
.B1(n_688),
.B2(n_683),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1921),
.Y(n_2145)
);

A2O1A1Ixp33_ASAP7_75t_L g2146 ( 
.A1(n_2051),
.A2(n_693),
.B(n_697),
.C(n_692),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1981),
.A2(n_693),
.B1(n_697),
.B2(n_692),
.Y(n_2147)
);

NAND3xp33_ASAP7_75t_L g2148 ( 
.A(n_2001),
.B(n_698),
.C(n_587),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1948),
.A2(n_698),
.B1(n_592),
.B2(n_597),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_2029),
.A2(n_604),
.B1(n_606),
.B2(n_584),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1948),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2031),
.A2(n_616),
.B1(n_618),
.B2(n_610),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1922),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2056),
.B(n_1866),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2009),
.A2(n_453),
.B1(n_457),
.B2(n_452),
.Y(n_2155)
);

NAND3xp33_ASAP7_75t_L g2156 ( 
.A(n_2009),
.B(n_457),
.C(n_453),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_1954),
.B(n_1858),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_1934),
.A2(n_636),
.B1(n_637),
.B2(n_630),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2002),
.B(n_1815),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1969),
.B(n_1815),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_1934),
.A2(n_636),
.B1(n_637),
.B2(n_630),
.Y(n_2161)
);

AOI22xp33_ASAP7_75t_L g2162 ( 
.A1(n_1934),
.A2(n_649),
.B1(n_665),
.B2(n_643),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_1995),
.B(n_1858),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_SL g2164 ( 
.A1(n_1941),
.A2(n_649),
.B(n_643),
.Y(n_2164)
);

OAI221xp5_ASAP7_75t_SL g2165 ( 
.A1(n_2016),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_2165)
);

A2O1A1Ixp33_ASAP7_75t_L g2166 ( 
.A1(n_2052),
.A2(n_673),
.B(n_678),
.C(n_665),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_1964),
.B(n_36),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1922),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_1945),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2052),
.A2(n_678),
.B1(n_682),
.B2(n_673),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_2039),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_1954),
.B(n_1878),
.Y(n_2172)
);

OAI221xp5_ASAP7_75t_L g2173 ( 
.A1(n_2050),
.A2(n_687),
.B1(n_682),
.B2(n_490),
.C(n_492),
.Y(n_2173)
);

AO21x2_ASAP7_75t_L g2174 ( 
.A1(n_1985),
.A2(n_1883),
.B(n_1879),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_SL g2175 ( 
.A1(n_2039),
.A2(n_687),
.B1(n_486),
.B2(n_497),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_1937),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1949),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_1996),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1996),
.B(n_1894),
.Y(n_2179)
);

OAI211xp5_ASAP7_75t_L g2180 ( 
.A1(n_2055),
.A2(n_499),
.B(n_511),
.C(n_482),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1932),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_2053),
.A2(n_513),
.B1(n_520),
.B2(n_512),
.Y(n_2182)
);

OAI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2058),
.A2(n_531),
.B1(n_535),
.B2(n_522),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2058),
.A2(n_542),
.B1(n_545),
.B2(n_537),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1932),
.Y(n_2185)
);

OAI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2039),
.A2(n_566),
.B1(n_568),
.B2(n_556),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2053),
.A2(n_572),
.B1(n_573),
.B2(n_570),
.Y(n_2187)
);

AOI221xp5_ASAP7_75t_L g2188 ( 
.A1(n_2013),
.A2(n_617),
.B1(n_607),
.B2(n_590),
.C(n_588),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1940),
.B(n_1879),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2013),
.A2(n_575),
.B1(n_577),
.B2(n_574),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2020),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_2039),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_1933),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.C(n_48),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_1957),
.B(n_1883),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2014),
.B(n_1894),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2007),
.A2(n_947),
.B1(n_943),
.B2(n_1782),
.Y(n_2196)
);

AOI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2007),
.A2(n_947),
.B1(n_943),
.B2(n_1782),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2022),
.B(n_1800),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1949),
.Y(n_2199)
);

INVx4_ASAP7_75t_SL g2200 ( 
.A(n_2039),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2020),
.A2(n_50),
.B1(n_45),
.B2(n_49),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1966),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2007),
.A2(n_947),
.B1(n_943),
.B2(n_1800),
.Y(n_2203)
);

AOI33xp33_ASAP7_75t_L g2204 ( 
.A1(n_1933),
.A2(n_49),
.A3(n_50),
.B1(n_51),
.B2(n_52),
.B3(n_53),
.Y(n_2204)
);

OAI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_2008),
.A2(n_54),
.B1(n_51),
.B2(n_52),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1949),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2011),
.A2(n_947),
.B1(n_943),
.B2(n_915),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1957),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_1962),
.B(n_55),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2062),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2200),
.B(n_2046),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2092),
.B(n_2008),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2068),
.B(n_2024),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2063),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_2122),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2208),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2065),
.B(n_2018),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2076),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2081),
.B(n_1912),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2108),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2109),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2075),
.B(n_2032),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2115),
.Y(n_2223)
);

INVx2_ASAP7_75t_SL g2224 ( 
.A(n_2171),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2065),
.B(n_2018),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2125),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_2178),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2169),
.B(n_1925),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_2151),
.Y(n_2229)
);

NAND2x1_ASAP7_75t_L g2230 ( 
.A(n_2067),
.B(n_1944),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2101),
.B(n_2018),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2176),
.B(n_1927),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2098),
.B(n_2033),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2095),
.B(n_1929),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2145),
.Y(n_2235)
);

INVxp67_ASAP7_75t_SL g2236 ( 
.A(n_2159),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2132),
.B(n_1977),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2153),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2168),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2070),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2064),
.A2(n_2042),
.B1(n_2011),
.B2(n_1955),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2177),
.B(n_1944),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2181),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2185),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2200),
.B(n_1944),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2074),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2080),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2129),
.A2(n_2042),
.B1(n_2011),
.B2(n_1955),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2104),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2137),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2111),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2202),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2172),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2198),
.B(n_2054),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2177),
.B(n_1961),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2085),
.B(n_2061),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2085),
.B(n_1915),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2189),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2061),
.B(n_1915),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2189),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2096),
.B(n_1916),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_2073),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2209),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_SL g2264 ( 
.A1(n_2066),
.A2(n_1941),
.B1(n_1926),
.B2(n_1959),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2199),
.B(n_1961),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2194),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_2100),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2157),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2071),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2199),
.B(n_1961),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2077),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2073),
.Y(n_2272)
);

BUFx2_ASAP7_75t_SL g2273 ( 
.A(n_2123),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2096),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_2060),
.A2(n_1941),
.B1(n_2010),
.B2(n_1959),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2110),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2110),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2136),
.B(n_2054),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2124),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2124),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_2171),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2116),
.B(n_2112),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2087),
.B(n_1916),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2195),
.B(n_2091),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2160),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2160),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2114),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2103),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_2163),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2102),
.B(n_1949),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2171),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2206),
.B(n_1949),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2094),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2117),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2084),
.B(n_2072),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2159),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2090),
.B(n_1955),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_2200),
.B(n_2042),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2192),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2192),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2192),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2090),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2090),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2179),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2131),
.B(n_1955),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2128),
.Y(n_2306)
);

BUFx2_ASAP7_75t_L g2307 ( 
.A(n_2093),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2130),
.B(n_1955),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2123),
.B(n_2133),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2094),
.Y(n_2310)
);

NOR2x1p5_ASAP7_75t_L g2311 ( 
.A(n_2133),
.B(n_2042),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2130),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2100),
.B(n_2042),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2100),
.B(n_1962),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2099),
.B(n_1963),
.Y(n_2315)
);

OAI22xp5_ASAP7_75t_SL g2316 ( 
.A1(n_2167),
.A2(n_1923),
.B1(n_1935),
.B2(n_2057),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2127),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2127),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2121),
.B(n_2047),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_SL g2320 ( 
.A1(n_2086),
.A2(n_1923),
.B1(n_1935),
.B2(n_2057),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2127),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2154),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2082),
.Y(n_2323)
);

AND2x2_ASAP7_75t_SL g2324 ( 
.A(n_2204),
.B(n_2047),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2154),
.B(n_1963),
.Y(n_2325)
);

INVx2_ASAP7_75t_SL g2326 ( 
.A(n_2174),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2174),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2105),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2105),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2078),
.B(n_1965),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2069),
.B(n_1936),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2088),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2140),
.Y(n_2333)
);

AOI22xp33_ASAP7_75t_L g2334 ( 
.A1(n_2060),
.A2(n_1959),
.B1(n_2010),
.B2(n_1926),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2088),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2219),
.B(n_1965),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2264),
.B(n_2241),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2308),
.B(n_1923),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2210),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_2251),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2257),
.B(n_1928),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2211),
.B(n_1936),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2214),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2218),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2220),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2330),
.B(n_2212),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_2212),
.B(n_2092),
.Y(n_2347)
);

OR2x2_ASAP7_75t_L g2348 ( 
.A(n_2315),
.B(n_1928),
.Y(n_2348)
);

OAI21xp5_ASAP7_75t_SL g2349 ( 
.A1(n_2264),
.A2(n_2083),
.B(n_2193),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2221),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2223),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2226),
.Y(n_2352)
);

OAI221xp5_ASAP7_75t_L g2353 ( 
.A1(n_2334),
.A2(n_2165),
.B1(n_2089),
.B2(n_2138),
.C(n_2164),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2235),
.Y(n_2354)
);

INVx4_ASAP7_75t_L g2355 ( 
.A(n_2267),
.Y(n_2355)
);

OR2x2_ASAP7_75t_L g2356 ( 
.A(n_2213),
.B(n_1918),
.Y(n_2356)
);

BUFx2_ASAP7_75t_L g2357 ( 
.A(n_2215),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2263),
.B(n_2121),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2238),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2283),
.B(n_2147),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2308),
.B(n_1923),
.Y(n_2361)
);

NOR2x1_ASAP7_75t_SL g2362 ( 
.A(n_2215),
.B(n_2147),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2239),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2326),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2328),
.B(n_2079),
.Y(n_2365)
);

AND2x4_ASAP7_75t_L g2366 ( 
.A(n_2211),
.B(n_1935),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2329),
.B(n_2107),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2297),
.B(n_1935),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2243),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2326),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2319),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2244),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2297),
.B(n_2106),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2237),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2228),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2211),
.B(n_1985),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2293),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2305),
.B(n_2097),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2232),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2305),
.B(n_2015),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2332),
.B(n_2118),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2298),
.B(n_2311),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2245),
.B(n_2015),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2234),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2216),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2230),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2216),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_2251),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2314),
.B(n_2148),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2293),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2227),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2227),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2217),
.B(n_1918),
.Y(n_2393)
);

NOR2xp67_ASAP7_75t_L g2394 ( 
.A(n_2256),
.B(n_2205),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2299),
.B(n_2037),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2310),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2225),
.B(n_1924),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2222),
.Y(n_2398)
);

OR2x6_ASAP7_75t_SL g2399 ( 
.A(n_2229),
.B(n_2205),
.Y(n_2399)
);

BUFx2_ASAP7_75t_L g2400 ( 
.A(n_2298),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2262),
.B(n_1924),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2245),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2246),
.Y(n_2403)
);

INVxp67_ASAP7_75t_SL g2404 ( 
.A(n_2335),
.Y(n_2404)
);

INVxp67_ASAP7_75t_SL g2405 ( 
.A(n_2335),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2272),
.B(n_2313),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2245),
.B(n_2015),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2298),
.B(n_1986),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2306),
.B(n_2015),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2284),
.B(n_1973),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2289),
.B(n_2015),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2300),
.B(n_2037),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2233),
.B(n_1973),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2259),
.B(n_2003),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2289),
.B(n_2015),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2247),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2249),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2250),
.Y(n_2418)
);

INVx4_ASAP7_75t_L g2419 ( 
.A(n_2267),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2302),
.B(n_2015),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2310),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2301),
.B(n_2037),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2303),
.B(n_2015),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2319),
.B(n_2037),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2312),
.B(n_1974),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2252),
.Y(n_2426)
);

BUFx2_ASAP7_75t_L g2427 ( 
.A(n_2309),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2331),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2242),
.B(n_1974),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2322),
.Y(n_2430)
);

INVxp33_ASAP7_75t_L g2431 ( 
.A(n_2320),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2242),
.B(n_1983),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2331),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2331),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2325),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2318),
.B(n_1983),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2261),
.B(n_2037),
.Y(n_2437)
);

BUFx2_ASAP7_75t_L g2438 ( 
.A(n_2307),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2240),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2240),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2318),
.B(n_1993),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2254),
.B(n_2003),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_2224),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2224),
.B(n_2281),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2281),
.B(n_2191),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_2304),
.B(n_1993),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2290),
.B(n_2113),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_2317),
.B(n_2321),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2438),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2349),
.A2(n_2324),
.B(n_2248),
.Y(n_2450)
);

AOI33xp33_ASAP7_75t_L g2451 ( 
.A1(n_2399),
.A2(n_2334),
.A3(n_2275),
.B1(n_2144),
.B2(n_2126),
.B3(n_2120),
.Y(n_2451)
);

OAI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_2431),
.A2(n_2275),
.B1(n_2324),
.B2(n_2273),
.Y(n_2452)
);

OR2x2_ASAP7_75t_L g2453 ( 
.A(n_2371),
.B(n_2282),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2406),
.B(n_2292),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2357),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2340),
.Y(n_2456)
);

BUFx2_ASAP7_75t_L g2457 ( 
.A(n_2382),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_SL g2458 ( 
.A1(n_2362),
.A2(n_2201),
.B(n_2191),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2400),
.B(n_2322),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2382),
.B(n_2322),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2382),
.B(n_2231),
.Y(n_2461)
);

OAI31xp33_ASAP7_75t_SL g2462 ( 
.A1(n_2337),
.A2(n_2201),
.A3(n_2180),
.B(n_2323),
.Y(n_2462)
);

AO21x2_ASAP7_75t_L g2463 ( 
.A1(n_2337),
.A2(n_2236),
.B(n_2327),
.Y(n_2463)
);

OR2x2_ASAP7_75t_L g2464 ( 
.A(n_2398),
.B(n_2278),
.Y(n_2464)
);

OAI221xp5_ASAP7_75t_L g2465 ( 
.A1(n_2347),
.A2(n_2316),
.B1(n_2149),
.B2(n_2134),
.C(n_2146),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2399),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2340),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2368),
.B(n_2295),
.Y(n_2468)
);

OAI33xp33_ASAP7_75t_L g2469 ( 
.A1(n_2360),
.A2(n_2260),
.A3(n_2258),
.B1(n_2285),
.B2(n_2286),
.B3(n_2296),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2388),
.Y(n_2470)
);

INVx1_ASAP7_75t_SL g2471 ( 
.A(n_2427),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2430),
.Y(n_2472)
);

OAI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2431),
.A2(n_2291),
.B1(n_2294),
.B2(n_2170),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2355),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_L g2475 ( 
.A(n_2347),
.B(n_2119),
.C(n_2142),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2368),
.B(n_2291),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_2353),
.A2(n_2173),
.B1(n_2188),
.B2(n_2156),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2388),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_2394),
.A2(n_2367),
.B1(n_2346),
.B2(n_2365),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_SL g2480 ( 
.A(n_2358),
.B(n_2229),
.C(n_2149),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2338),
.B(n_2255),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2391),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2391),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2430),
.Y(n_2484)
);

AOI221xp5_ASAP7_75t_L g2485 ( 
.A1(n_2404),
.A2(n_2236),
.B1(n_2184),
.B2(n_2183),
.C(n_2266),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2392),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2445),
.B(n_2447),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2392),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2375),
.B(n_2379),
.Y(n_2489)
);

OAI321xp33_ASAP7_75t_L g2490 ( 
.A1(n_2424),
.A2(n_2333),
.A3(n_2175),
.B1(n_2183),
.B2(n_2184),
.C(n_2162),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2430),
.Y(n_2491)
);

AOI221x1_ASAP7_75t_L g2492 ( 
.A1(n_2355),
.A2(n_2277),
.B1(n_2279),
.B2(n_2276),
.C(n_2274),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2402),
.B(n_2288),
.Y(n_2493)
);

AOI211xp5_ASAP7_75t_L g2494 ( 
.A1(n_2405),
.A2(n_2381),
.B(n_2378),
.C(n_2373),
.Y(n_2494)
);

OAI211xp5_ASAP7_75t_L g2495 ( 
.A1(n_2378),
.A2(n_2166),
.B(n_2161),
.C(n_2158),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2402),
.B(n_2373),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2389),
.B(n_2374),
.C(n_2395),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2428),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2338),
.B(n_2265),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2339),
.Y(n_2500)
);

NOR3xp33_ASAP7_75t_SL g2501 ( 
.A(n_2444),
.B(n_2186),
.C(n_2280),
.Y(n_2501)
);

AOI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2384),
.A2(n_2269),
.B1(n_2287),
.B2(n_2288),
.Y(n_2502)
);

OR2x2_ASAP7_75t_L g2503 ( 
.A(n_2414),
.B(n_2271),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2343),
.Y(n_2504)
);

AOI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_2437),
.A2(n_2448),
.B1(n_2187),
.B2(n_2182),
.Y(n_2505)
);

AOI211xp5_ASAP7_75t_L g2506 ( 
.A1(n_2412),
.A2(n_2333),
.B(n_2268),
.C(n_2271),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2344),
.Y(n_2507)
);

OAI22xp5_ASAP7_75t_SL g2508 ( 
.A1(n_2355),
.A2(n_2190),
.B1(n_2141),
.B2(n_2139),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2345),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2350),
.Y(n_2510)
);

HB1xp67_ASAP7_75t_L g2511 ( 
.A(n_2377),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2351),
.Y(n_2512)
);

INVx5_ASAP7_75t_SL g2513 ( 
.A(n_2366),
.Y(n_2513)
);

INVx1_ASAP7_75t_SL g2514 ( 
.A(n_2443),
.Y(n_2514)
);

INVx1_ASAP7_75t_SL g2515 ( 
.A(n_2419),
.Y(n_2515)
);

OR2x2_ASAP7_75t_L g2516 ( 
.A(n_2341),
.B(n_2268),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2352),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2354),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2359),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2419),
.A2(n_2253),
.B1(n_2270),
.B2(n_2150),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2386),
.Y(n_2521)
);

NAND3xp33_ASAP7_75t_L g2522 ( 
.A(n_2422),
.B(n_2152),
.C(n_2253),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2361),
.B(n_1999),
.Y(n_2523)
);

OAI221xp5_ASAP7_75t_L g2524 ( 
.A1(n_2336),
.A2(n_2155),
.B1(n_2203),
.B2(n_2197),
.C(n_2196),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2361),
.B(n_1999),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2428),
.Y(n_2526)
);

OAI21x1_ASAP7_75t_L g2527 ( 
.A1(n_2386),
.A2(n_2143),
.B(n_1989),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2419),
.B(n_2000),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2433),
.Y(n_2529)
);

INVx4_ASAP7_75t_L g2530 ( 
.A(n_2386),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2366),
.B(n_1986),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2435),
.B(n_2000),
.Y(n_2532)
);

OAI21x1_ASAP7_75t_L g2533 ( 
.A1(n_2364),
.A2(n_1989),
.B(n_2135),
.Y(n_2533)
);

OAI33xp33_ASAP7_75t_L g2534 ( 
.A1(n_2363),
.A2(n_2027),
.A3(n_2043),
.B1(n_2034),
.B2(n_2030),
.B3(n_2004),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2366),
.B(n_2004),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_2342),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2457),
.B(n_2496),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2496),
.B(n_2448),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2454),
.B(n_2448),
.Y(n_2539)
);

AND2x4_ASAP7_75t_L g2540 ( 
.A(n_2530),
.B(n_2342),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2450),
.B(n_2435),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2521),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2511),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2511),
.Y(n_2544)
);

INVx1_ASAP7_75t_SL g2545 ( 
.A(n_2471),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2456),
.Y(n_2546)
);

OAI21xp5_ASAP7_75t_SL g2547 ( 
.A1(n_2462),
.A2(n_2407),
.B(n_2383),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2468),
.B(n_2342),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2460),
.B(n_2383),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2467),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2521),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2521),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2470),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2449),
.B(n_2369),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2449),
.B(n_2372),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2460),
.B(n_2407),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2487),
.B(n_2348),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2478),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2514),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2513),
.B(n_2380),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2455),
.B(n_2410),
.Y(n_2561)
);

NOR3xp33_ASAP7_75t_L g2562 ( 
.A(n_2451),
.B(n_2390),
.C(n_2377),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2474),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2482),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2483),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2455),
.B(n_2401),
.Y(n_2566)
);

NAND3xp33_ASAP7_75t_L g2567 ( 
.A(n_2480),
.B(n_2396),
.C(n_2390),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2513),
.B(n_2461),
.Y(n_2568)
);

OAI21xp5_ASAP7_75t_SL g2569 ( 
.A1(n_2452),
.A2(n_2380),
.B(n_2411),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2486),
.Y(n_2570)
);

OR2x6_ASAP7_75t_SL g2571 ( 
.A(n_2475),
.B(n_2396),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2513),
.B(n_2393),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2515),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2488),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2500),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2530),
.B(n_2433),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2451),
.B(n_2403),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2453),
.B(n_2416),
.Y(n_2578)
);

INVxp67_ASAP7_75t_SL g2579 ( 
.A(n_2466),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2504),
.Y(n_2580)
);

HB1xp67_ASAP7_75t_L g2581 ( 
.A(n_2463),
.Y(n_2581)
);

NAND2x1p5_ASAP7_75t_L g2582 ( 
.A(n_2530),
.B(n_1920),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2476),
.B(n_2481),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2459),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2459),
.B(n_2434),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2499),
.B(n_2434),
.Y(n_2586)
);

NAND2x1p5_ASAP7_75t_L g2587 ( 
.A(n_2466),
.B(n_1920),
.Y(n_2587)
);

AOI33xp33_ASAP7_75t_L g2588 ( 
.A1(n_2479),
.A2(n_2421),
.A3(n_2426),
.B1(n_2417),
.B2(n_2418),
.B3(n_2439),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2536),
.B(n_2408),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2493),
.B(n_2535),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2479),
.B(n_2425),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2472),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2507),
.Y(n_2593)
);

AO21x2_ASAP7_75t_L g2594 ( 
.A1(n_2463),
.A2(n_2370),
.B(n_2364),
.Y(n_2594)
);

OR2x2_ASAP7_75t_L g2595 ( 
.A(n_2464),
.B(n_2442),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2494),
.B(n_2425),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2472),
.B(n_2408),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2484),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2493),
.B(n_2408),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2505),
.B(n_2429),
.Y(n_2600)
);

O2A1O1Ixp33_ASAP7_75t_L g2601 ( 
.A1(n_2490),
.A2(n_2421),
.B(n_2370),
.C(n_2387),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2535),
.B(n_2420),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2509),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2484),
.B(n_2420),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2520),
.B(n_2397),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2491),
.B(n_2440),
.Y(n_2606)
);

AND2x4_ASAP7_75t_SL g2607 ( 
.A(n_2480),
.B(n_2376),
.Y(n_2607)
);

NOR2x1_ASAP7_75t_L g2608 ( 
.A(n_2458),
.B(n_2440),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2510),
.Y(n_2609)
);

AOI21xp33_ASAP7_75t_L g2610 ( 
.A1(n_2522),
.A2(n_2495),
.B(n_2497),
.Y(n_2610)
);

OAI222xp33_ASAP7_75t_L g2611 ( 
.A1(n_2505),
.A2(n_2411),
.B1(n_2415),
.B2(n_2423),
.C1(n_2385),
.C2(n_2356),
.Y(n_2611)
);

NAND4xp25_ASAP7_75t_SL g2612 ( 
.A(n_2458),
.B(n_2415),
.C(n_2423),
.D(n_2409),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2512),
.Y(n_2613)
);

BUFx2_ASAP7_75t_L g2614 ( 
.A(n_2491),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2523),
.B(n_2429),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2498),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2473),
.B(n_2432),
.Y(n_2617)
);

NAND2x1p5_ASAP7_75t_L g2618 ( 
.A(n_2498),
.B(n_2049),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2543),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2571),
.B(n_2517),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2544),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2571),
.B(n_2518),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2537),
.B(n_2501),
.Y(n_2623)
);

AOI21xp33_ASAP7_75t_L g2624 ( 
.A1(n_2608),
.A2(n_2465),
.B(n_2477),
.Y(n_2624)
);

INVx2_ASAP7_75t_SL g2625 ( 
.A(n_2540),
.Y(n_2625)
);

OR2x2_ASAP7_75t_L g2626 ( 
.A(n_2545),
.B(n_2489),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2616),
.Y(n_2627)
);

NAND2x1p5_ASAP7_75t_L g2628 ( 
.A(n_2559),
.B(n_2526),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2573),
.B(n_2591),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2537),
.B(n_2501),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2540),
.Y(n_2631)
);

NAND2xp67_ASAP7_75t_L g2632 ( 
.A(n_2563),
.B(n_2526),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2616),
.Y(n_2633)
);

OR2x2_ASAP7_75t_L g2634 ( 
.A(n_2579),
.B(n_2516),
.Y(n_2634)
);

HB1xp67_ASAP7_75t_L g2635 ( 
.A(n_2579),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2584),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2541),
.B(n_2503),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2584),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2598),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2540),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2592),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2598),
.Y(n_2642)
);

OR2x2_ASAP7_75t_L g2643 ( 
.A(n_2600),
.B(n_2519),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2610),
.B(n_2469),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2578),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2576),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2561),
.B(n_2529),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2546),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2550),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2553),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2617),
.B(n_2529),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2596),
.B(n_2502),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2566),
.B(n_2532),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2538),
.B(n_2525),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2539),
.B(n_2485),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2563),
.B(n_2477),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2568),
.B(n_2492),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2583),
.B(n_2531),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2562),
.B(n_2506),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2562),
.B(n_2528),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2588),
.B(n_2531),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2588),
.B(n_2436),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2558),
.B(n_2564),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2576),
.B(n_2376),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2548),
.B(n_2432),
.Y(n_2665)
);

INVxp67_ASAP7_75t_L g2666 ( 
.A(n_2585),
.Y(n_2666)
);

NAND2x2_ASAP7_75t_L g2667 ( 
.A(n_2577),
.B(n_2508),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2576),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2542),
.Y(n_2669)
);

NAND2xp33_ASAP7_75t_SL g2670 ( 
.A(n_2581),
.B(n_2413),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2548),
.B(n_2590),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2595),
.B(n_2436),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2557),
.B(n_2446),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2554),
.B(n_2441),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2565),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2555),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2590),
.B(n_2572),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2570),
.Y(n_2678)
);

OR2x2_ASAP7_75t_L g2679 ( 
.A(n_2567),
.B(n_2441),
.Y(n_2679)
);

OAI21xp5_ASAP7_75t_SL g2680 ( 
.A1(n_2607),
.A2(n_2611),
.B(n_2547),
.Y(n_2680)
);

INVx1_ASAP7_75t_SL g2681 ( 
.A(n_2641),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2635),
.B(n_2574),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2641),
.B(n_2668),
.Y(n_2683)
);

NOR2x2_ASAP7_75t_L g2684 ( 
.A(n_2631),
.B(n_2542),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2634),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2646),
.Y(n_2686)
);

OAI21xp5_ASAP7_75t_SL g2687 ( 
.A1(n_2624),
.A2(n_2607),
.B(n_2569),
.Y(n_2687)
);

OR2x2_ASAP7_75t_L g2688 ( 
.A(n_2629),
.B(n_2605),
.Y(n_2688)
);

OAI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2659),
.A2(n_2581),
.B1(n_2587),
.B2(n_2601),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2632),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2636),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2628),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2638),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2671),
.B(n_2560),
.Y(n_2694)
);

A2O1A1Ixp33_ASAP7_75t_L g2695 ( 
.A1(n_2624),
.A2(n_2560),
.B(n_2580),
.C(n_2575),
.Y(n_2695)
);

OR2x2_ASAP7_75t_L g2696 ( 
.A(n_2656),
.B(n_2593),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2646),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2627),
.Y(n_2698)
);

OR2x2_ASAP7_75t_L g2699 ( 
.A(n_2626),
.B(n_2603),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2633),
.Y(n_2700)
);

OR2x2_ASAP7_75t_L g2701 ( 
.A(n_2637),
.B(n_2609),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2644),
.A2(n_2612),
.B1(n_2586),
.B2(n_2585),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2639),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2623),
.B(n_2613),
.Y(n_2704)
);

AOI211xp5_ASAP7_75t_L g2705 ( 
.A1(n_2680),
.A2(n_2589),
.B(n_2614),
.C(n_2524),
.Y(n_2705)
);

AOI21xp33_ASAP7_75t_L g2706 ( 
.A1(n_2659),
.A2(n_2594),
.B(n_2552),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2630),
.B(n_2655),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2666),
.B(n_2586),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2625),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2620),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2677),
.B(n_2549),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2642),
.Y(n_2712)
);

O2A1O1Ixp33_ASAP7_75t_SL g2713 ( 
.A1(n_2680),
.A2(n_2552),
.B(n_2551),
.C(n_2594),
.Y(n_2713)
);

INVxp67_ASAP7_75t_SL g2714 ( 
.A(n_2620),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2669),
.Y(n_2715)
);

OAI31xp33_ASAP7_75t_L g2716 ( 
.A1(n_2657),
.A2(n_2587),
.A3(n_2589),
.B(n_2618),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2651),
.B(n_2551),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2652),
.A2(n_2618),
.B1(n_2582),
.B2(n_2599),
.Y(n_2718)
);

AOI21xp33_ASAP7_75t_L g2719 ( 
.A1(n_2622),
.A2(n_2606),
.B(n_2597),
.Y(n_2719)
);

NAND2x1p5_ASAP7_75t_L g2720 ( 
.A(n_2640),
.B(n_2599),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2647),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2657),
.B(n_2597),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2654),
.B(n_2658),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2645),
.B(n_2549),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2663),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2663),
.Y(n_2726)
);

INVxp67_ASAP7_75t_L g2727 ( 
.A(n_2622),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2681),
.B(n_2676),
.Y(n_2728)
);

INVx2_ASAP7_75t_SL g2729 ( 
.A(n_2720),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2720),
.Y(n_2730)
);

OAI21xp33_ASAP7_75t_L g2731 ( 
.A1(n_2687),
.A2(n_2702),
.B(n_2707),
.Y(n_2731)
);

INVxp67_ASAP7_75t_L g2732 ( 
.A(n_2722),
.Y(n_2732)
);

OR2x2_ASAP7_75t_L g2733 ( 
.A(n_2681),
.B(n_2662),
.Y(n_2733)
);

AOI32xp33_ASAP7_75t_SL g2734 ( 
.A1(n_2714),
.A2(n_2685),
.A3(n_2660),
.B1(n_2700),
.B2(n_2698),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2683),
.B(n_2662),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2708),
.Y(n_2736)
);

INVx2_ASAP7_75t_SL g2737 ( 
.A(n_2686),
.Y(n_2737)
);

O2A1O1Ixp33_ASAP7_75t_L g2738 ( 
.A1(n_2713),
.A2(n_2660),
.B(n_2661),
.C(n_2643),
.Y(n_2738)
);

AOI33xp33_ASAP7_75t_L g2739 ( 
.A1(n_2710),
.A2(n_2621),
.A3(n_2619),
.B1(n_2675),
.B2(n_2648),
.B3(n_2649),
.Y(n_2739)
);

OAI221xp5_ASAP7_75t_L g2740 ( 
.A1(n_2727),
.A2(n_2667),
.B1(n_2705),
.B2(n_2689),
.C(n_2710),
.Y(n_2740)
);

INVx1_ASAP7_75t_SL g2741 ( 
.A(n_2684),
.Y(n_2741)
);

INVxp67_ASAP7_75t_SL g2742 ( 
.A(n_2692),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_SL g2743 ( 
.A1(n_2689),
.A2(n_2679),
.B1(n_2658),
.B2(n_2664),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2697),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2724),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2682),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2694),
.A2(n_2670),
.B1(n_2664),
.B2(n_2665),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2721),
.Y(n_2748)
);

OAI221xp5_ASAP7_75t_L g2749 ( 
.A1(n_2716),
.A2(n_2653),
.B1(n_2674),
.B2(n_2650),
.C(n_2678),
.Y(n_2749)
);

AOI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2711),
.A2(n_2556),
.B1(n_2672),
.B2(n_2597),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2699),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2717),
.Y(n_2752)
);

OAI321xp33_ASAP7_75t_L g2753 ( 
.A1(n_2696),
.A2(n_2673),
.A3(n_2582),
.B1(n_2556),
.B2(n_2604),
.C(n_2602),
.Y(n_2753)
);

NOR3xp33_ASAP7_75t_SL g2754 ( 
.A(n_2695),
.B(n_2534),
.C(n_2606),
.Y(n_2754)
);

O2A1O1Ixp33_ASAP7_75t_L g2755 ( 
.A1(n_2706),
.A2(n_2606),
.B(n_2604),
.C(n_2602),
.Y(n_2755)
);

OAI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2688),
.A2(n_2615),
.B1(n_2376),
.B2(n_2409),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2709),
.Y(n_2757)
);

OAI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2690),
.A2(n_2027),
.B1(n_2028),
.B2(n_2021),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2723),
.A2(n_2527),
.B1(n_2533),
.B2(n_2010),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2719),
.B(n_2533),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2701),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2704),
.B(n_2527),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2719),
.B(n_56),
.Y(n_2763)
);

OAI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2706),
.A2(n_2049),
.B(n_2040),
.Y(n_2764)
);

NOR4xp25_ASAP7_75t_SL g2765 ( 
.A(n_2715),
.B(n_58),
.C(n_56),
.D(n_57),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2741),
.B(n_2691),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2741),
.B(n_2693),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2728),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2742),
.B(n_2725),
.Y(n_2769)
);

AOI221xp5_ASAP7_75t_L g2770 ( 
.A1(n_2740),
.A2(n_2726),
.B1(n_2712),
.B2(n_2703),
.C(n_2718),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2732),
.B(n_2731),
.Y(n_2771)
);

NOR2xp67_ASAP7_75t_L g2772 ( 
.A(n_2729),
.B(n_2718),
.Y(n_2772)
);

AOI221xp5_ASAP7_75t_L g2773 ( 
.A1(n_2738),
.A2(n_2207),
.B1(n_60),
.B2(n_61),
.C(n_62),
.Y(n_2773)
);

O2A1O1Ixp33_ASAP7_75t_SL g2774 ( 
.A1(n_2763),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2752),
.Y(n_2775)
);

INVx1_ASAP7_75t_SL g2776 ( 
.A(n_2730),
.Y(n_2776)
);

OAI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2743),
.A2(n_2040),
.B(n_2025),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2757),
.Y(n_2778)
);

OAI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2747),
.A2(n_2028),
.B1(n_2030),
.B2(n_2021),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_2733),
.Y(n_2780)
);

OAI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2735),
.A2(n_2043),
.B1(n_2044),
.B2(n_2034),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2737),
.Y(n_2782)
);

OAI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2750),
.A2(n_2044),
.B1(n_1938),
.B2(n_1947),
.Y(n_2783)
);

OAI321xp33_ASAP7_75t_L g2784 ( 
.A1(n_2749),
.A2(n_62),
.A3(n_63),
.B1(n_64),
.B2(n_65),
.C(n_66),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2739),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2761),
.Y(n_2786)
);

AOI22xp33_ASAP7_75t_SL g2787 ( 
.A1(n_2751),
.A2(n_1913),
.B1(n_1931),
.B2(n_1938),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2744),
.B(n_63),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2748),
.B(n_2745),
.Y(n_2789)
);

INVx1_ASAP7_75t_SL g2790 ( 
.A(n_2760),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2765),
.B(n_65),
.Y(n_2791)
);

AOI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2756),
.A2(n_2736),
.B1(n_2754),
.B2(n_2746),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2762),
.B(n_2765),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2755),
.B(n_66),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2758),
.Y(n_2795)
);

NOR3xp33_ASAP7_75t_L g2796 ( 
.A(n_2753),
.B(n_67),
.C(n_68),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2764),
.B(n_2734),
.Y(n_2797)
);

AOI21xp33_ASAP7_75t_L g2798 ( 
.A1(n_2780),
.A2(n_2753),
.B(n_2759),
.Y(n_2798)
);

AOI221xp5_ASAP7_75t_L g2799 ( 
.A1(n_2796),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.C(n_74),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2772),
.B(n_2776),
.Y(n_2800)
);

OAI21xp5_ASAP7_75t_SL g2801 ( 
.A1(n_2792),
.A2(n_69),
.B(n_74),
.Y(n_2801)
);

NAND4xp25_ASAP7_75t_L g2802 ( 
.A(n_2771),
.B(n_77),
.C(n_75),
.D(n_76),
.Y(n_2802)
);

AOI221xp5_ASAP7_75t_L g2803 ( 
.A1(n_2773),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.C(n_82),
.Y(n_2803)
);

OAI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2780),
.A2(n_1946),
.B1(n_1952),
.B2(n_1947),
.Y(n_2804)
);

NOR3xp33_ASAP7_75t_L g2805 ( 
.A(n_2784),
.B(n_78),
.C(n_79),
.Y(n_2805)
);

AOI33xp33_ASAP7_75t_L g2806 ( 
.A1(n_2785),
.A2(n_82),
.A3(n_83),
.B1(n_85),
.B2(n_86),
.B3(n_88),
.Y(n_2806)
);

AOI322xp5_ASAP7_75t_L g2807 ( 
.A1(n_2770),
.A2(n_1946),
.A3(n_1952),
.B1(n_88),
.B2(n_89),
.C1(n_90),
.C2(n_91),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2776),
.B(n_83),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2797),
.A2(n_1913),
.B(n_85),
.Y(n_2809)
);

NAND3xp33_ASAP7_75t_L g2810 ( 
.A(n_2793),
.B(n_90),
.C(n_92),
.Y(n_2810)
);

AOI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2794),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.C(n_98),
.Y(n_2811)
);

AOI21xp5_ASAP7_75t_SL g2812 ( 
.A1(n_2791),
.A2(n_2766),
.B(n_2788),
.Y(n_2812)
);

OAI21xp33_ASAP7_75t_L g2813 ( 
.A1(n_2768),
.A2(n_2025),
.B(n_2026),
.Y(n_2813)
);

NAND3xp33_ASAP7_75t_SL g2814 ( 
.A(n_2767),
.B(n_94),
.C(n_95),
.Y(n_2814)
);

OAI31xp33_ASAP7_75t_L g2815 ( 
.A1(n_2790),
.A2(n_97),
.A3(n_98),
.B(n_99),
.Y(n_2815)
);

AOI221xp5_ASAP7_75t_L g2816 ( 
.A1(n_2790),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.C(n_103),
.Y(n_2816)
);

NOR3xp33_ASAP7_75t_L g2817 ( 
.A(n_2786),
.B(n_101),
.C(n_104),
.Y(n_2817)
);

OAI211xp5_ASAP7_75t_L g2818 ( 
.A1(n_2775),
.A2(n_104),
.B(n_106),
.C(n_107),
.Y(n_2818)
);

AOI211xp5_ASAP7_75t_L g2819 ( 
.A1(n_2769),
.A2(n_107),
.B(n_108),
.C(n_109),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2782),
.Y(n_2820)
);

OAI21xp5_ASAP7_75t_SL g2821 ( 
.A1(n_2778),
.A2(n_111),
.B(n_112),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2774),
.B(n_2795),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2800),
.Y(n_2823)
);

AOI211xp5_ASAP7_75t_L g2824 ( 
.A1(n_2798),
.A2(n_2789),
.B(n_2777),
.C(n_2779),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2808),
.B(n_2781),
.Y(n_2825)
);

AOI211x1_ASAP7_75t_L g2826 ( 
.A1(n_2810),
.A2(n_2783),
.B(n_2787),
.C(n_115),
.Y(n_2826)
);

OAI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2801),
.A2(n_111),
.B(n_114),
.Y(n_2827)
);

AOI21xp33_ASAP7_75t_L g2828 ( 
.A1(n_2822),
.A2(n_116),
.B(n_117),
.Y(n_2828)
);

OAI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2820),
.A2(n_1931),
.B1(n_117),
.B2(n_118),
.Y(n_2829)
);

A2O1A1Ixp33_ASAP7_75t_L g2830 ( 
.A1(n_2799),
.A2(n_116),
.B(n_118),
.C(n_119),
.Y(n_2830)
);

HB1xp67_ASAP7_75t_L g2831 ( 
.A(n_2814),
.Y(n_2831)
);

AOI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2805),
.A2(n_1913),
.B1(n_1931),
.B2(n_2036),
.Y(n_2832)
);

AOI221xp5_ASAP7_75t_L g2833 ( 
.A1(n_2812),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.C(n_124),
.Y(n_2833)
);

OAI32xp33_ASAP7_75t_L g2834 ( 
.A1(n_2817),
.A2(n_2802),
.A3(n_2807),
.B1(n_2806),
.B2(n_2815),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2809),
.A2(n_120),
.B(n_123),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2819),
.B(n_124),
.Y(n_2836)
);

OAI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2821),
.A2(n_125),
.B(n_126),
.Y(n_2837)
);

AOI21xp33_ASAP7_75t_SL g2838 ( 
.A1(n_2818),
.A2(n_126),
.B(n_130),
.Y(n_2838)
);

NOR3xp33_ASAP7_75t_L g2839 ( 
.A(n_2803),
.B(n_131),
.C(n_132),
.Y(n_2839)
);

INVxp33_ASAP7_75t_SL g2840 ( 
.A(n_2811),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2816),
.B(n_131),
.Y(n_2841)
);

AOI221xp5_ASAP7_75t_L g2842 ( 
.A1(n_2834),
.A2(n_2804),
.B1(n_2813),
.B2(n_134),
.C(n_135),
.Y(n_2842)
);

O2A1O1Ixp33_ASAP7_75t_L g2843 ( 
.A1(n_2838),
.A2(n_132),
.B(n_133),
.C(n_136),
.Y(n_2843)
);

OAI221xp5_ASAP7_75t_L g2844 ( 
.A1(n_2824),
.A2(n_133),
.B1(n_136),
.B2(n_138),
.C(n_139),
.Y(n_2844)
);

AOI32xp33_ASAP7_75t_L g2845 ( 
.A1(n_2823),
.A2(n_138),
.A3(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_2845)
);

OAI21xp33_ASAP7_75t_L g2846 ( 
.A1(n_2840),
.A2(n_2036),
.B(n_2026),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2831),
.Y(n_2847)
);

AOI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2839),
.A2(n_1931),
.B1(n_142),
.B2(n_143),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2836),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2825),
.Y(n_2850)
);

AOI211xp5_ASAP7_75t_L g2851 ( 
.A1(n_2828),
.A2(n_140),
.B(n_143),
.C(n_144),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2841),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_2852)
);

OAI221xp5_ASAP7_75t_L g2853 ( 
.A1(n_2833),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.C(n_149),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2837),
.Y(n_2854)
);

NOR3xp33_ASAP7_75t_L g2855 ( 
.A(n_2847),
.B(n_2833),
.C(n_2827),
.Y(n_2855)
);

OAI211xp5_ASAP7_75t_SL g2856 ( 
.A1(n_2842),
.A2(n_2835),
.B(n_2830),
.C(n_2832),
.Y(n_2856)
);

AOI31xp33_ASAP7_75t_L g2857 ( 
.A1(n_2851),
.A2(n_2829),
.A3(n_2826),
.B(n_152),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2845),
.B(n_2852),
.Y(n_2858)
);

NOR2xp67_ASAP7_75t_L g2859 ( 
.A(n_2854),
.B(n_150),
.Y(n_2859)
);

XNOR2x1_ASAP7_75t_L g2860 ( 
.A(n_2850),
.B(n_151),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2844),
.A2(n_154),
.B1(n_156),
.B2(n_158),
.Y(n_2861)
);

AOI211xp5_ASAP7_75t_L g2862 ( 
.A1(n_2843),
.A2(n_154),
.B(n_159),
.C(n_160),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2853),
.B(n_159),
.Y(n_2863)
);

O2A1O1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2849),
.A2(n_160),
.B(n_161),
.C(n_162),
.Y(n_2864)
);

AO22x2_ASAP7_75t_L g2865 ( 
.A1(n_2848),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_2865)
);

OAI21xp5_ASAP7_75t_SL g2866 ( 
.A1(n_2846),
.A2(n_165),
.B(n_166),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2847),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2867),
.B(n_167),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2859),
.Y(n_2869)
);

NOR2x1_ASAP7_75t_L g2870 ( 
.A(n_2860),
.B(n_168),
.Y(n_2870)
);

INVxp33_ASAP7_75t_SL g2871 ( 
.A(n_2855),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2865),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2863),
.B(n_168),
.Y(n_2873)
);

INVxp67_ASAP7_75t_L g2874 ( 
.A(n_2865),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2858),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2864),
.Y(n_2876)
);

OAI221xp5_ASAP7_75t_L g2877 ( 
.A1(n_2866),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.C(n_173),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2856),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_2878)
);

OR2x2_ASAP7_75t_L g2879 ( 
.A(n_2861),
.B(n_174),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2862),
.B(n_175),
.Y(n_2880)
);

AOI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2857),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2859),
.B(n_178),
.Y(n_2882)
);

OAI211xp5_ASAP7_75t_SL g2883 ( 
.A1(n_2858),
.A2(n_179),
.B(n_180),
.C(n_181),
.Y(n_2883)
);

AND2x4_ASAP7_75t_L g2884 ( 
.A(n_2859),
.B(n_179),
.Y(n_2884)
);

INVxp33_ASAP7_75t_SL g2885 ( 
.A(n_2870),
.Y(n_2885)
);

NOR2x1_ASAP7_75t_L g2886 ( 
.A(n_2884),
.B(n_182),
.Y(n_2886)
);

NOR2xp67_ASAP7_75t_L g2887 ( 
.A(n_2874),
.B(n_183),
.Y(n_2887)
);

NOR3xp33_ASAP7_75t_L g2888 ( 
.A(n_2875),
.B(n_183),
.C(n_186),
.Y(n_2888)
);

NAND4xp75_ASAP7_75t_L g2889 ( 
.A(n_2869),
.B(n_188),
.C(n_189),
.D(n_191),
.Y(n_2889)
);

NAND4xp75_ASAP7_75t_L g2890 ( 
.A(n_2881),
.B(n_188),
.C(n_189),
.D(n_194),
.Y(n_2890)
);

NAND2x1p5_ASAP7_75t_L g2891 ( 
.A(n_2884),
.B(n_194),
.Y(n_2891)
);

OR3x2_ASAP7_75t_L g2892 ( 
.A(n_2876),
.B(n_195),
.C(n_197),
.Y(n_2892)
);

NOR2x1_ASAP7_75t_L g2893 ( 
.A(n_2882),
.B(n_195),
.Y(n_2893)
);

OAI22xp5_ASAP7_75t_SL g2894 ( 
.A1(n_2871),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2868),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2872),
.Y(n_2896)
);

INVx1_ASAP7_75t_SL g2897 ( 
.A(n_2879),
.Y(n_2897)
);

NOR2xp67_ASAP7_75t_L g2898 ( 
.A(n_2877),
.B(n_198),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2878),
.Y(n_2899)
);

NOR3xp33_ASAP7_75t_SL g2900 ( 
.A(n_2896),
.B(n_2883),
.C(n_2873),
.Y(n_2900)
);

OR3x2_ASAP7_75t_L g2901 ( 
.A(n_2899),
.B(n_2895),
.C(n_2892),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2891),
.Y(n_2902)
);

NOR3xp33_ASAP7_75t_L g2903 ( 
.A(n_2897),
.B(n_2880),
.C(n_217),
.Y(n_2903)
);

NAND3x1_ASAP7_75t_L g2904 ( 
.A(n_2886),
.B(n_215),
.C(n_221),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2887),
.B(n_223),
.Y(n_2905)
);

OAI221xp5_ASAP7_75t_R g2906 ( 
.A1(n_2885),
.A2(n_225),
.B1(n_226),
.B2(n_230),
.C(n_231),
.Y(n_2906)
);

NAND5xp2_ASAP7_75t_L g2907 ( 
.A(n_2888),
.B(n_237),
.C(n_238),
.D(n_239),
.E(n_248),
.Y(n_2907)
);

OAI221xp5_ASAP7_75t_SL g2908 ( 
.A1(n_2898),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.C(n_264),
.Y(n_2908)
);

NAND5xp2_ASAP7_75t_L g2909 ( 
.A(n_2893),
.B(n_265),
.C(n_267),
.D(n_272),
.E(n_276),
.Y(n_2909)
);

HB1xp67_ASAP7_75t_L g2910 ( 
.A(n_2889),
.Y(n_2910)
);

INVx1_ASAP7_75t_SL g2911 ( 
.A(n_2894),
.Y(n_2911)
);

INVx4_ASAP7_75t_L g2912 ( 
.A(n_2902),
.Y(n_2912)
);

AND3x1_ASAP7_75t_L g2913 ( 
.A(n_2900),
.B(n_2890),
.C(n_279),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2910),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2904),
.Y(n_2915)
);

OR2x2_ASAP7_75t_L g2916 ( 
.A(n_2909),
.B(n_278),
.Y(n_2916)
);

XNOR2xp5_ASAP7_75t_L g2917 ( 
.A(n_2911),
.B(n_283),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2905),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2903),
.B(n_285),
.Y(n_2919)
);

BUFx12f_ASAP7_75t_L g2920 ( 
.A(n_2901),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2907),
.Y(n_2921)
);

INVx1_ASAP7_75t_SL g2922 ( 
.A(n_2906),
.Y(n_2922)
);

OR3x1_ASAP7_75t_L g2923 ( 
.A(n_2914),
.B(n_2908),
.C(n_293),
.Y(n_2923)
);

NAND3xp33_ASAP7_75t_L g2924 ( 
.A(n_2912),
.B(n_947),
.C(n_910),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2917),
.B(n_287),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2916),
.Y(n_2926)
);

HB1xp67_ASAP7_75t_L g2927 ( 
.A(n_2913),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2919),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2915),
.B(n_2921),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2922),
.B(n_296),
.Y(n_2930)
);

BUFx2_ASAP7_75t_L g2931 ( 
.A(n_2920),
.Y(n_2931)
);

OAI21xp5_ASAP7_75t_SL g2932 ( 
.A1(n_2918),
.A2(n_298),
.B(n_299),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2917),
.Y(n_2933)
);

HB1xp67_ASAP7_75t_L g2934 ( 
.A(n_2917),
.Y(n_2934)
);

AOI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2930),
.A2(n_921),
.B(n_915),
.Y(n_2935)
);

AOI22xp33_ASAP7_75t_L g2936 ( 
.A1(n_2931),
.A2(n_915),
.B1(n_910),
.B2(n_921),
.Y(n_2936)
);

XNOR2xp5_ASAP7_75t_L g2937 ( 
.A(n_2923),
.B(n_301),
.Y(n_2937)
);

HB1xp67_ASAP7_75t_L g2938 ( 
.A(n_2925),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2928),
.B(n_304),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2934),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2927),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_SL g2942 ( 
.A1(n_2933),
.A2(n_1226),
.B1(n_311),
.B2(n_316),
.Y(n_2942)
);

XNOR2xp5_ASAP7_75t_L g2943 ( 
.A(n_2937),
.B(n_2929),
.Y(n_2943)
);

AOI22x1_ASAP7_75t_L g2944 ( 
.A1(n_2940),
.A2(n_2929),
.B1(n_2926),
.B2(n_2932),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2939),
.Y(n_2945)
);

AND2x4_ASAP7_75t_L g2946 ( 
.A(n_2941),
.B(n_2924),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2938),
.B(n_306),
.Y(n_2947)
);

INVx3_ASAP7_75t_SL g2948 ( 
.A(n_2935),
.Y(n_2948)
);

OAI22x1_ASAP7_75t_L g2949 ( 
.A1(n_2942),
.A2(n_317),
.B1(n_320),
.B2(n_324),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2936),
.Y(n_2950)
);

NOR2x1p5_ASAP7_75t_L g2951 ( 
.A(n_2939),
.B(n_921),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2937),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2941),
.A2(n_1289),
.B1(n_1241),
.B2(n_1239),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2941),
.A2(n_1226),
.B1(n_910),
.B2(n_921),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2937),
.Y(n_2955)
);

XNOR2x2_ASAP7_75t_L g2956 ( 
.A(n_2937),
.B(n_325),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2937),
.Y(n_2957)
);

OAI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2941),
.A2(n_915),
.B1(n_910),
.B2(n_882),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2937),
.B(n_327),
.Y(n_2959)
);

AND2x4_ASAP7_75t_L g2960 ( 
.A(n_2957),
.B(n_2952),
.Y(n_2960)
);

OAI22xp5_ASAP7_75t_SL g2961 ( 
.A1(n_2959),
.A2(n_328),
.B1(n_329),
.B2(n_331),
.Y(n_2961)
);

NOR2x1_ASAP7_75t_L g2962 ( 
.A(n_2947),
.B(n_332),
.Y(n_2962)
);

BUFx6f_ASAP7_75t_L g2963 ( 
.A(n_2955),
.Y(n_2963)
);

XNOR2xp5_ASAP7_75t_L g2964 ( 
.A(n_2943),
.B(n_334),
.Y(n_2964)
);

AO22x2_ASAP7_75t_L g2965 ( 
.A1(n_2945),
.A2(n_340),
.B1(n_342),
.B2(n_344),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2951),
.B(n_347),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2956),
.Y(n_2967)
);

OAI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2944),
.A2(n_2950),
.B1(n_2946),
.B2(n_2948),
.Y(n_2968)
);

NOR2x1_ASAP7_75t_L g2969 ( 
.A(n_2954),
.B(n_349),
.Y(n_2969)
);

BUFx2_ASAP7_75t_L g2970 ( 
.A(n_2949),
.Y(n_2970)
);

INVxp67_ASAP7_75t_SL g2971 ( 
.A(n_2958),
.Y(n_2971)
);

OAI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2953),
.A2(n_915),
.B1(n_889),
.B2(n_882),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2959),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2963),
.A2(n_889),
.B1(n_868),
.B2(n_882),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2962),
.B(n_354),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2966),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2964),
.B(n_355),
.Y(n_2977)
);

AOI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2968),
.A2(n_889),
.B(n_882),
.Y(n_2978)
);

AOI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2967),
.A2(n_889),
.B(n_882),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2965),
.Y(n_2980)
);

OAI22xp5_ASAP7_75t_L g2981 ( 
.A1(n_2970),
.A2(n_889),
.B1(n_868),
.B2(n_861),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2969),
.B(n_356),
.Y(n_2982)
);

OAI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2960),
.A2(n_868),
.B1(n_861),
.B2(n_859),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2973),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_2975),
.B(n_2971),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_SL g2986 ( 
.A1(n_2982),
.A2(n_2972),
.B(n_2961),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2980),
.B(n_2977),
.Y(n_2987)
);

AOI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2984),
.A2(n_868),
.B(n_923),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2976),
.A2(n_2978),
.B(n_2979),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2981),
.B(n_358),
.Y(n_2990)
);

AOI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2983),
.A2(n_2974),
.B1(n_1289),
.B2(n_1241),
.Y(n_2991)
);

XNOR2xp5_ASAP7_75t_L g2992 ( 
.A(n_2987),
.B(n_359),
.Y(n_2992)
);

OAI21xp5_ASAP7_75t_SL g2993 ( 
.A1(n_2985),
.A2(n_362),
.B(n_365),
.Y(n_2993)
);

AOI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2990),
.A2(n_1289),
.B1(n_1241),
.B2(n_1239),
.Y(n_2994)
);

AOI222xp33_ASAP7_75t_L g2995 ( 
.A1(n_2993),
.A2(n_2986),
.B1(n_2991),
.B2(n_2989),
.C1(n_2988),
.C2(n_1289),
.Y(n_2995)
);

AOI22xp33_ASAP7_75t_L g2996 ( 
.A1(n_2992),
.A2(n_962),
.B1(n_1239),
.B2(n_1241),
.Y(n_2996)
);

AO21x2_ASAP7_75t_L g2997 ( 
.A1(n_2995),
.A2(n_2994),
.B(n_962),
.Y(n_2997)
);

AOI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_2997),
.A2(n_2996),
.B(n_923),
.Y(n_2998)
);

AOI211xp5_ASAP7_75t_L g2999 ( 
.A1(n_2998),
.A2(n_861),
.B(n_859),
.C(n_854),
.Y(n_2999)
);


endmodule