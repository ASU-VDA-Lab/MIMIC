module fake_jpeg_11812_n_64 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_16),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_28),
.B1(n_11),
.B2(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_21),
.B1(n_17),
.B2(n_8),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_20),
.B1(n_17),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_8),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_20),
.B1(n_22),
.B2(n_12),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_20),
.B1(n_1),
.B2(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_3),
.Y(n_43)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_38),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_44),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_41),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_48),
.Y(n_57)
);

AOI31xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.A3(n_51),
.B(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_52),
.Y(n_58)
);

MAJx2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_60),
.C(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_43),
.B1(n_35),
.B2(n_39),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_39),
.B(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_7),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_1),
.Y(n_64)
);


endmodule