module fake_jpeg_16941_n_69 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_44),
.B1(n_9),
.B2(n_10),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_12),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_45),
.B1(n_17),
.B2(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.C(n_56),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_59),
.Y(n_69)
);


endmodule