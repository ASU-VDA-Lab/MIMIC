module real_aes_6603_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_140;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g470 ( .A(n_1), .Y(n_470) );
INVx1_ASAP7_75t_L g254 ( .A(n_2), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_3), .A2(n_38), .B1(n_204), .B2(n_509), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_4), .B(n_447), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g215 ( .A1(n_5), .A2(n_137), .B(n_216), .Y(n_215) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_6), .B(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_6), .B(n_159), .Y(n_495) );
AND2x6_ASAP7_75t_L g142 ( .A(n_7), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_8), .A2(n_136), .B(n_144), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_9), .B(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_9), .B(n_39), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_10), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g221 ( .A(n_11), .Y(n_221) );
INVx1_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
INVx1_ASAP7_75t_L g464 ( .A(n_13), .Y(n_464) );
INVx1_ASAP7_75t_L g154 ( .A(n_14), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_15), .B(n_228), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_16), .B(n_160), .Y(n_497) );
AO32x2_ASAP7_75t_L g543 ( .A1(n_17), .A2(n_159), .A3(n_175), .B1(n_483), .B2(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_18), .B(n_204), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_19), .B(n_171), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_20), .B(n_160), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_21), .A2(n_50), .B1(n_204), .B2(n_509), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_22), .B(n_137), .Y(n_164) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_23), .A2(n_78), .B1(n_204), .B2(n_228), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_24), .B(n_204), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_25), .B(n_214), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_26), .A2(n_151), .B(n_153), .C(n_155), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_27), .A2(n_105), .B1(n_117), .B2(n_750), .Y(n_104) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_28), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_29), .B(n_130), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_30), .B(n_186), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_31), .A2(n_102), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_31), .Y(n_738) );
INVx1_ASAP7_75t_L g233 ( .A(n_32), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_33), .B(n_130), .Y(n_521) );
INVx2_ASAP7_75t_L g140 ( .A(n_34), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_35), .B(n_204), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_36), .B(n_130), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_37), .A2(n_142), .B(n_147), .C(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g116 ( .A(n_39), .Y(n_116) );
INVx1_ASAP7_75t_L g231 ( .A(n_40), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_41), .B(n_186), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_42), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_42), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_43), .B(n_204), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_44), .A2(n_88), .B1(n_156), .B2(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_45), .B(n_204), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_46), .B(n_204), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_47), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_48), .B(n_469), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_49), .B(n_137), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_51), .A2(n_61), .B1(n_204), .B2(n_228), .Y(n_501) );
OAI22xp5_ASAP7_75t_SL g432 ( .A1(n_52), .A2(n_433), .B1(n_436), .B2(n_437), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_52), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_53), .A2(n_147), .B1(n_228), .B2(n_230), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_54), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_55), .B(n_204), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_56), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_57), .B(n_204), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_58), .A2(n_219), .B(n_220), .C(n_222), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_59), .Y(n_190) );
INVx1_ASAP7_75t_L g217 ( .A(n_60), .Y(n_217) );
INVx1_ASAP7_75t_L g143 ( .A(n_62), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_63), .A2(n_736), .B1(n_739), .B2(n_740), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_63), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_64), .B(n_204), .Y(n_471) );
INVx1_ASAP7_75t_L g133 ( .A(n_65), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g433 ( .A1(n_66), .A2(n_77), .B1(n_434), .B2(n_435), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_66), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
AO32x2_ASAP7_75t_L g506 ( .A1(n_68), .A2(n_159), .A3(n_196), .B1(n_483), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g481 ( .A(n_69), .Y(n_481) );
INVx1_ASAP7_75t_L g516 ( .A(n_70), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_SL g241 ( .A1(n_71), .A2(n_171), .B(n_222), .C(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g243 ( .A(n_72), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_73), .B(n_228), .Y(n_517) );
INVx1_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_75), .Y(n_236) );
INVx1_ASAP7_75t_L g181 ( .A(n_76), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_77), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_79), .A2(n_142), .B(n_147), .C(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_80), .B(n_509), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_81), .B(n_228), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_82), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_84), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_85), .B(n_228), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_86), .A2(n_142), .B(n_147), .C(n_253), .Y(n_252) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_87), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g442 ( .A(n_87), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g452 ( .A(n_87), .B(n_444), .Y(n_452) );
INVx2_ASAP7_75t_L g730 ( .A(n_87), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_89), .A2(n_103), .B1(n_228), .B2(n_229), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_90), .B(n_130), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_91), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_92), .A2(n_142), .B(n_147), .C(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_93), .Y(n_207) );
INVx1_ASAP7_75t_L g240 ( .A(n_94), .Y(n_240) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_95), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_96), .B(n_168), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_97), .B(n_228), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_98), .B(n_159), .Y(n_158) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_99), .A2(n_451), .B1(n_731), .B2(n_732), .C1(n_741), .C2(n_744), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_101), .A2(n_137), .B(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_102), .Y(n_737) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g752 ( .A(n_107), .Y(n_752) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_114), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g444 ( .A(n_110), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_120), .B(n_449), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g749 ( .A(n_119), .Y(n_749) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_439), .B(n_446), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_431), .B1(n_432), .B2(n_438), .Y(n_122) );
INVx2_ASAP7_75t_SL g438 ( .A(n_123), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_123), .A2(n_452), .B1(n_454), .B2(n_742), .Y(n_741) );
OR4x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_327), .C(n_386), .D(n_413), .Y(n_123) );
NAND3xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_269), .C(n_294), .Y(n_124) );
O2A1O1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_192), .B(n_212), .C(n_245), .Y(n_125) );
AOI211xp5_ASAP7_75t_SL g417 ( .A1(n_126), .A2(n_418), .B(n_420), .C(n_423), .Y(n_417) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_161), .Y(n_126) );
INVx1_ASAP7_75t_L g292 ( .A(n_127), .Y(n_292) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g267 ( .A(n_128), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g299 ( .A(n_128), .Y(n_299) );
AND2x2_ASAP7_75t_L g354 ( .A(n_128), .B(n_323), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_128), .B(n_210), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_128), .B(n_211), .Y(n_412) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g273 ( .A(n_129), .Y(n_273) );
AND2x2_ASAP7_75t_L g316 ( .A(n_129), .B(n_179), .Y(n_316) );
AND2x2_ASAP7_75t_L g334 ( .A(n_129), .B(n_211), .Y(n_334) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_135), .B(n_158), .Y(n_129) );
INVx1_ASAP7_75t_L g191 ( .A(n_130), .Y(n_191) );
INVx2_ASAP7_75t_L g196 ( .A(n_130), .Y(n_196) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_130), .A2(n_514), .B(n_521), .Y(n_513) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_130), .A2(n_523), .B(n_531), .Y(n_522) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_L g160 ( .A(n_131), .B(n_132), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_138), .B(n_142), .Y(n_182) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g469 ( .A(n_139), .Y(n_469) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx1_ASAP7_75t_L g229 ( .A(n_140), .Y(n_229) );
INVx1_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
INVx3_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
INVx4_ASAP7_75t_SL g157 ( .A(n_142), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_142), .A2(n_463), .B(n_467), .Y(n_462) );
BUFx3_ASAP7_75t_L g483 ( .A(n_142), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_142), .A2(n_489), .B(n_492), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_142), .A2(n_515), .B(n_518), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_142), .A2(n_524), .B(n_528), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_150), .C(n_157), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_146), .A2(n_157), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_146), .A2(n_157), .B(n_240), .C(n_241), .Y(n_239) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_148), .Y(n_204) );
INVx1_ASAP7_75t_L g509 ( .A(n_148), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_151), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g466 ( .A(n_151), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_151), .A2(n_519), .B(n_520), .Y(n_518) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g230 ( .A1(n_152), .A2(n_231), .B1(n_232), .B2(n_233), .Y(n_230) );
INVx2_ASAP7_75t_L g232 ( .A(n_152), .Y(n_232) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_157), .A2(n_182), .B1(n_227), .B2(n_234), .Y(n_226) );
INVx4_ASAP7_75t_L g178 ( .A(n_159), .Y(n_178) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_159), .A2(n_238), .B(n_244), .Y(n_237) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_159), .A2(n_488), .B(n_495), .Y(n_487) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g175 ( .A(n_160), .Y(n_175) );
INVx4_ASAP7_75t_L g266 ( .A(n_161), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_161), .A2(n_322), .B(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_L g402 ( .A(n_161), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_179), .Y(n_161) );
INVx1_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
AND2x2_ASAP7_75t_L g271 ( .A(n_162), .B(n_211), .Y(n_271) );
OR2x2_ASAP7_75t_L g300 ( .A(n_162), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g314 ( .A(n_162), .Y(n_314) );
INVx3_ASAP7_75t_L g323 ( .A(n_162), .Y(n_323) );
AND2x2_ASAP7_75t_L g333 ( .A(n_162), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g366 ( .A(n_162), .B(n_272), .Y(n_366) );
AND2x2_ASAP7_75t_L g390 ( .A(n_162), .B(n_346), .Y(n_390) );
OR2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_176), .Y(n_162) );
AOI21xp5_ASAP7_75t_SL g163 ( .A1(n_164), .A2(n_165), .B(n_174), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_172), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_168), .A2(n_254), .B(n_255), .C(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g472 ( .A(n_168), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_168), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_168), .A2(n_490), .B(n_491), .Y(n_489) );
O2A1O1Ixp5_ASAP7_75t_SL g515 ( .A1(n_168), .A2(n_222), .B(n_516), .C(n_517), .Y(n_515) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_169), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_169), .B(n_243), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g507 ( .A1(n_169), .A2(n_186), .B1(n_508), .B2(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g527 ( .A(n_171), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_172), .A2(n_185), .B(n_187), .Y(n_184) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g188 ( .A(n_174), .Y(n_188) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_174), .A2(n_462), .B(n_473), .Y(n_461) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_174), .A2(n_476), .B(n_484), .Y(n_475) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_175), .A2(n_226), .B(n_235), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_175), .B(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_175), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx3_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_178), .B(n_483), .C(n_499), .Y(n_498) );
AO21x1_ASAP7_75t_L g577 ( .A1(n_178), .A2(n_499), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
AND2x2_ASAP7_75t_L g426 ( .A(n_179), .B(n_268), .Y(n_426) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_188), .B(n_189), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_182), .A2(n_251), .B(n_252), .Y(n_250) );
INVx4_ASAP7_75t_L g202 ( .A(n_186), .Y(n_202) );
INVx2_ASAP7_75t_L g219 ( .A(n_186), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_186), .A2(n_472), .B1(n_500), .B2(n_501), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_186), .A2(n_472), .B1(n_545), .B2(n_546), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_191), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_191), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_208), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_194), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g346 ( .A(n_194), .B(n_334), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_194), .B(n_323), .Y(n_408) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g268 ( .A(n_195), .Y(n_268) );
AND2x2_ASAP7_75t_L g272 ( .A(n_195), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g313 ( .A(n_195), .B(n_314), .Y(n_313) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_206), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_205), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_203), .Y(n_199) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g222 ( .A(n_204), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_208), .B(n_309), .Y(n_331) );
INVx1_ASAP7_75t_L g370 ( .A(n_208), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_208), .B(n_297), .Y(n_414) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AND2x2_ASAP7_75t_L g277 ( .A(n_209), .B(n_272), .Y(n_277) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_211), .B(n_268), .Y(n_301) );
INVx1_ASAP7_75t_L g380 ( .A(n_211), .Y(n_380) );
AOI322xp5_ASAP7_75t_L g404 ( .A1(n_212), .A2(n_319), .A3(n_379), .B1(n_405), .B2(n_407), .C1(n_409), .C2(n_411), .Y(n_404) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_213), .B(n_224), .Y(n_212) );
AND2x2_ASAP7_75t_L g259 ( .A(n_213), .B(n_237), .Y(n_259) );
INVx1_ASAP7_75t_SL g262 ( .A(n_213), .Y(n_262) );
AND2x2_ASAP7_75t_L g264 ( .A(n_213), .B(n_225), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_213), .B(n_281), .Y(n_287) );
INVx2_ASAP7_75t_L g306 ( .A(n_213), .Y(n_306) );
AND2x2_ASAP7_75t_L g319 ( .A(n_213), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g357 ( .A(n_213), .B(n_281), .Y(n_357) );
BUFx2_ASAP7_75t_L g374 ( .A(n_213), .Y(n_374) );
AND2x2_ASAP7_75t_L g388 ( .A(n_213), .B(n_248), .Y(n_388) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_223), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_L g480 ( .A1(n_219), .A2(n_468), .B(n_481), .C(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_219), .A2(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_224), .B(n_276), .Y(n_303) );
AND2x2_ASAP7_75t_L g430 ( .A(n_224), .B(n_306), .Y(n_430) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_237), .Y(n_224) );
OR2x2_ASAP7_75t_L g275 ( .A(n_225), .B(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
AND2x2_ASAP7_75t_L g326 ( .A(n_225), .B(n_249), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_225), .B(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_225), .Y(n_410) );
INVx2_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g261 ( .A(n_237), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
BUFx2_ASAP7_75t_L g289 ( .A(n_237), .Y(n_289) );
AND2x2_ASAP7_75t_L g308 ( .A(n_237), .B(n_281), .Y(n_308) );
INVx3_ASAP7_75t_L g320 ( .A(n_237), .Y(n_320) );
OR2x2_ASAP7_75t_L g330 ( .A(n_237), .B(n_281), .Y(n_330) );
AOI31xp33_ASAP7_75t_SL g245 ( .A1(n_246), .A2(n_260), .A3(n_263), .B(n_265), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_259), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_247), .B(n_282), .Y(n_293) );
OR2x2_ASAP7_75t_L g317 ( .A(n_247), .B(n_287), .Y(n_317) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_248), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g338 ( .A(n_248), .B(n_330), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_248), .B(n_320), .Y(n_348) );
AND2x2_ASAP7_75t_L g355 ( .A(n_248), .B(n_356), .Y(n_355) );
NAND2x1_ASAP7_75t_L g383 ( .A(n_248), .B(n_319), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_248), .B(n_374), .Y(n_384) );
AND2x2_ASAP7_75t_L g396 ( .A(n_248), .B(n_281), .Y(n_396) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g276 ( .A(n_249), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_256), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g342 ( .A(n_259), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_259), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_261), .B(n_337), .Y(n_371) );
AND2x4_ASAP7_75t_L g282 ( .A(n_262), .B(n_283), .Y(n_282) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g361 ( .A(n_267), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_267), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_299), .Y(n_309) );
AND2x2_ASAP7_75t_L g403 ( .A(n_268), .B(n_273), .Y(n_403) );
INVx1_ASAP7_75t_L g428 ( .A(n_268), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .B1(n_277), .B2(n_278), .C(n_284), .Y(n_269) );
CKINVDCx14_ASAP7_75t_R g290 ( .A(n_270), .Y(n_290) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_271), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_274), .B(n_325), .Y(n_344) );
INVx3_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g393 ( .A(n_275), .B(n_289), .Y(n_393) );
AND2x2_ASAP7_75t_L g307 ( .A(n_276), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g337 ( .A(n_276), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_276), .B(n_320), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_276), .B(n_377), .C(n_408), .Y(n_407) );
AOI211xp5_ASAP7_75t_SL g340 ( .A1(n_277), .A2(n_341), .B(n_343), .C(n_351), .Y(n_340) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp33_ASAP7_75t_L g329 ( .A1(n_279), .A2(n_330), .B1(n_331), .B2(n_332), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_280), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_280), .B(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g422 ( .A(n_282), .B(n_396), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_290), .B1(n_291), .B2(n_293), .Y(n_284) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_288), .B(n_337), .Y(n_368) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_291), .A2(n_383), .B1(n_414), .B2(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_302), .B1(n_304), .B2(n_309), .C(n_310), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI221xp5_ASAP7_75t_L g310 ( .A1(n_300), .A2(n_311), .B1(n_317), .B2(n_318), .C(n_321), .Y(n_310) );
INVx1_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_SL g325 ( .A(n_306), .Y(n_325) );
OR2x2_ASAP7_75t_L g398 ( .A(n_306), .B(n_330), .Y(n_398) );
AND2x2_ASAP7_75t_L g400 ( .A(n_306), .B(n_308), .Y(n_400) );
INVx1_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_312), .A2(n_370), .B(n_371), .Y(n_369) );
OR2x2_ASAP7_75t_L g376 ( .A(n_312), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_334), .Y(n_350) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_318), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_319), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_320), .B(n_356), .Y(n_419) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_323), .A2(n_336), .B(n_338), .C(n_339), .Y(n_335) );
NAND2x1_ASAP7_75t_SL g360 ( .A(n_323), .B(n_361), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_324), .A2(n_373), .B1(n_375), .B2(n_378), .Y(n_372) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_326), .B(n_416), .Y(n_415) );
NAND5xp2_ASAP7_75t_L g327 ( .A(n_328), .B(n_340), .C(n_358), .D(n_372), .E(n_381), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_329), .B(n_335), .Y(n_328) );
INVx1_ASAP7_75t_L g385 ( .A(n_331), .Y(n_385) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_333), .A2(n_352), .B1(n_392), .B2(n_394), .C(n_397), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_334), .B(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_337), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_337), .B(n_403), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B1(n_347), .B2(n_349), .Y(n_343) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g425 ( .A(n_354), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_366), .B2(n_367), .C(n_369), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g409 ( .A(n_364), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g416 ( .A(n_374), .Y(n_416) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_384), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_389), .B(n_391), .C(n_404), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_414), .B(n_415), .C(n_417), .Y(n_413) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_393), .B(n_395), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_427), .B(n_429), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_433), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_438), .A2(n_452), .B1(n_453), .B2(n_729), .Y(n_451) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_442), .Y(n_448) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_443), .B(n_730), .Y(n_746) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g729 ( .A(n_444), .B(n_730), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_446), .B(n_450), .C(n_747), .Y(n_449) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR5x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_620), .C(n_678), .D(n_714), .E(n_721), .Y(n_456) );
NAND3xp33_ASAP7_75t_SL g457 ( .A(n_458), .B(n_566), .C(n_590), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_502), .B1(n_532), .B2(n_537), .C(n_547), .Y(n_458) );
OAI21xp5_ASAP7_75t_SL g700 ( .A1(n_459), .A2(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_485), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_460), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_474), .Y(n_460) );
INVx2_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
AND2x2_ASAP7_75t_L g549 ( .A(n_461), .B(n_487), .Y(n_549) );
AND2x2_ASAP7_75t_L g603 ( .A(n_461), .B(n_486), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_461), .B(n_475), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B(n_471), .C(n_472), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_472), .A2(n_493), .B(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g636 ( .A(n_474), .B(n_577), .Y(n_636) );
AND2x2_ASAP7_75t_L g669 ( .A(n_474), .B(n_487), .Y(n_669) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g576 ( .A(n_475), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g589 ( .A(n_475), .B(n_487), .Y(n_589) );
AND2x2_ASAP7_75t_L g596 ( .A(n_475), .B(n_577), .Y(n_596) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_475), .Y(n_605) );
AND2x2_ASAP7_75t_L g612 ( .A(n_475), .B(n_486), .Y(n_612) );
INVx1_ASAP7_75t_L g643 ( .A(n_475), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_480), .B(n_483), .Y(n_476) );
INVx1_ASAP7_75t_L g619 ( .A(n_485), .Y(n_619) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
INVx2_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
AND2x2_ASAP7_75t_L g597 ( .A(n_486), .B(n_536), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_486), .B(n_643), .Y(n_648) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_487), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g720 ( .A(n_487), .B(n_684), .Y(n_720) );
INVx2_ASAP7_75t_L g534 ( .A(n_496), .Y(n_534) );
INVx3_ASAP7_75t_L g635 ( .A(n_496), .Y(n_635) );
OR2x2_ASAP7_75t_L g665 ( .A(n_496), .B(n_666), .Y(n_665) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_496), .B(n_575), .Y(n_691) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g578 ( .A(n_497), .Y(n_578) );
AOI33xp33_ASAP7_75t_L g711 ( .A1(n_502), .A2(n_549), .A3(n_563), .B1(n_635), .B2(n_712), .B3(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_511), .Y(n_503) );
OR2x2_ASAP7_75t_L g564 ( .A(n_504), .B(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_504), .B(n_561), .Y(n_623) );
OR2x2_ASAP7_75t_L g676 ( .A(n_504), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g602 ( .A(n_505), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g627 ( .A(n_505), .B(n_511), .Y(n_627) );
AND2x2_ASAP7_75t_L g694 ( .A(n_505), .B(n_539), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_505), .A2(n_594), .B(n_720), .Y(n_719) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
INVx1_ASAP7_75t_L g554 ( .A(n_506), .Y(n_554) );
AND2x2_ASAP7_75t_L g573 ( .A(n_506), .B(n_543), .Y(n_573) );
AND2x2_ASAP7_75t_L g622 ( .A(n_506), .B(n_542), .Y(n_622) );
INVx2_ASAP7_75t_SL g664 ( .A(n_511), .Y(n_664) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
INVx2_ASAP7_75t_L g584 ( .A(n_512), .Y(n_584) );
INVx1_ASAP7_75t_L g715 ( .A(n_512), .Y(n_715) );
AND2x2_ASAP7_75t_L g728 ( .A(n_512), .B(n_609), .Y(n_728) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g555 ( .A(n_513), .Y(n_555) );
OR2x2_ASAP7_75t_L g561 ( .A(n_513), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_513), .Y(n_572) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_522), .Y(n_539) );
AND2x2_ASAP7_75t_L g556 ( .A(n_522), .B(n_542), .Y(n_556) );
INVx1_ASAP7_75t_L g562 ( .A(n_522), .Y(n_562) );
INVx1_ASAP7_75t_L g569 ( .A(n_522), .Y(n_569) );
AND2x2_ASAP7_75t_L g594 ( .A(n_522), .B(n_543), .Y(n_594) );
INVx2_ASAP7_75t_L g610 ( .A(n_522), .Y(n_610) );
AND2x2_ASAP7_75t_L g703 ( .A(n_522), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_522), .B(n_584), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_527), .Y(n_524) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g558 ( .A(n_534), .Y(n_558) );
INVx1_ASAP7_75t_L g587 ( .A(n_534), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_534), .B(n_618), .Y(n_684) );
INVx1_ASAP7_75t_SL g644 ( .A(n_535), .Y(n_644) );
INVx2_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
AND2x2_ASAP7_75t_L g634 ( .A(n_536), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g650 ( .A(n_536), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g712 ( .A(n_538), .Y(n_712) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g567 ( .A(n_540), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g670 ( .A(n_540), .B(n_660), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_540), .A2(n_681), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g583 ( .A(n_541), .B(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
INVx1_ASAP7_75t_L g632 ( .A(n_541), .Y(n_632) );
OR2x2_ASAP7_75t_L g696 ( .A(n_542), .B(n_555), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_542), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g609 ( .A(n_543), .B(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g616 ( .A(n_543), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_550), .B1(n_557), .B2(n_559), .Y(n_547) );
OR2x2_ASAP7_75t_L g626 ( .A(n_548), .B(n_576), .Y(n_626) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_549), .A2(n_668), .B1(n_670), .B2(n_671), .C1(n_672), .C2(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g614 ( .A(n_553), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_555), .B(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_555), .Y(n_639) );
AND2x2_ASAP7_75t_L g687 ( .A(n_555), .B(n_556), .Y(n_687) );
INVx1_ASAP7_75t_L g705 ( .A(n_555), .Y(n_705) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g671 ( .A(n_558), .B(n_597), .Y(n_671) );
AND2x2_ASAP7_75t_L g713 ( .A(n_558), .B(n_589), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_560), .B(n_608), .Y(n_695) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_561), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g588 ( .A(n_565), .B(n_589), .Y(n_588) );
INVx3_ASAP7_75t_L g656 ( .A(n_565), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_570), .B(n_574), .C(n_579), .Y(n_566) );
INVxp67_ASAP7_75t_L g580 ( .A(n_567), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_568), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_568), .B(n_615), .Y(n_710) );
BUFx3_ASAP7_75t_L g674 ( .A(n_569), .Y(n_674) );
INVx1_ASAP7_75t_L g581 ( .A(n_570), .Y(n_581) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g600 ( .A(n_572), .B(n_594), .Y(n_600) );
INVx1_ASAP7_75t_SL g640 ( .A(n_573), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g630 ( .A(n_575), .Y(n_630) );
AND2x2_ASAP7_75t_L g653 ( .A(n_575), .B(n_636), .Y(n_653) );
INVx1_ASAP7_75t_SL g624 ( .A(n_576), .Y(n_624) );
INVx1_ASAP7_75t_L g651 ( .A(n_577), .Y(n_651) );
AOI31xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .A3(n_582), .B(n_585), .Y(n_579) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g672 ( .A(n_583), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g646 ( .A(n_584), .Y(n_646) );
BUFx2_ASAP7_75t_L g660 ( .A(n_584), .Y(n_660) );
AND2x2_ASAP7_75t_L g688 ( .A(n_584), .B(n_609), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_SL g661 ( .A(n_588), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_589), .B(n_656), .Y(n_702) );
AND2x2_ASAP7_75t_L g709 ( .A(n_589), .B(n_635), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_595), .B(n_598), .C(n_613), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_595), .A2(n_622), .B1(n_623), .B2(n_624), .C(n_625), .Y(n_621) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g629 ( .A(n_596), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g666 ( .A(n_597), .Y(n_666) );
OAI32xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .A3(n_604), .B1(n_606), .B2(n_611), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_600), .A2(n_653), .B(n_654), .C(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_608), .A2(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g677 ( .A(n_609), .Y(n_677) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_615), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g663 ( .A(n_615), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g680 ( .A(n_617), .Y(n_680) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NAND4xp25_ASAP7_75t_SL g620 ( .A(n_621), .B(n_633), .C(n_652), .D(n_667), .Y(n_620) );
AND2x2_ASAP7_75t_L g659 ( .A(n_622), .B(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g681 ( .A(n_622), .B(n_674), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_624), .B(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_628), .B2(n_631), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_626), .A2(n_677), .B1(n_708), .B2(n_710), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g714 ( .A1(n_626), .A2(n_715), .B(n_716), .C(n_719), .Y(n_714) );
INVx2_ASAP7_75t_L g685 ( .A(n_627), .Y(n_685) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_629), .A2(n_663), .B1(n_680), .B2(n_681), .C1(n_682), .C2(n_685), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_637), .C(n_641), .Y(n_633) );
INVx1_ASAP7_75t_L g699 ( .A(n_634), .Y(n_699) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_638), .A2(n_642), .B1(n_645), .B2(n_647), .Y(n_641) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g668 ( .A(n_650), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g726 ( .A(n_653), .Y(n_726) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_662), .B2(n_665), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_660), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g717 ( .A(n_665), .Y(n_717) );
INVx1_ASAP7_75t_L g698 ( .A(n_669), .Y(n_698) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_671), .Y(n_725) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND5xp2_ASAP7_75t_L g678 ( .A(n_679), .B(n_686), .C(n_700), .D(n_706), .E(n_711), .Y(n_678) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B(n_689), .C(n_692), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI31xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .A3(n_696), .B(n_697), .Y(n_692) );
INVx1_ASAP7_75t_L g718 ( .A(n_694), .Y(n_718) );
OR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI222xp33_ASAP7_75t_L g721 ( .A1(n_708), .A2(n_710), .B1(n_722), .B2(n_725), .C1(n_726), .C2(n_727), .Y(n_721) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g743 ( .A(n_729), .Y(n_743) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g739 ( .A(n_736), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
endmodule