module fake_jpeg_17494_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_28),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_12),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_18),
.B(n_17),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_24),
.B(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_23),
.B1(n_15),
.B2(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_17),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_53),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_25),
.B(n_2),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_31),
.B1(n_27),
.B2(n_16),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_55),
.B1(n_42),
.B2(n_13),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_14),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_37),
.B(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_19),
.C(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_19),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_15),
.B1(n_16),
.B2(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_42),
.B1(n_53),
.B2(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_66),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_10),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_45),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_72),
.B1(n_71),
.B2(n_75),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_65),
.B1(n_57),
.B2(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_52),
.B1(n_34),
.B2(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_59),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_49),
.C(n_46),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_78),
.C(n_54),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_1),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_82),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_78),
.B1(n_76),
.B2(n_4),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_5),
.C(n_8),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_87),
.B(n_79),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_93),
.B(n_3),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_86),
.B1(n_80),
.B2(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_1),
.B(n_3),
.Y(n_98)
);

AOI21x1_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_88),
.B(n_89),
.Y(n_99)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_9),
.B(n_11),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_98),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_101),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.B(n_1),
.Y(n_108)
);


endmodule