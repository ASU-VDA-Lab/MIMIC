module fake_netlist_1_202_n_22 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_22;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_9), .B(n_5), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_17), .B(n_11), .C(n_12), .Y(n_18) );
NAND4xp25_ASAP7_75t_L g19 ( .A(n_18), .B(n_14), .C(n_1), .D(n_2), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_19), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_22) );
endmodule