module fake_jpeg_29696_n_330 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_49),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_68),
.Y(n_106)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_32),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_8),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_76),
.B(n_37),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_42),
.B1(n_65),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_77),
.A2(n_85),
.B1(n_90),
.B2(n_111),
.Y(n_157)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_83),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_42),
.B1(n_31),
.B2(n_36),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_29),
.B(n_25),
.C(n_43),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_31),
.B(n_32),
.C(n_39),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_31),
.B1(n_36),
.B2(n_32),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_95),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_109),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_43),
.B1(n_28),
.B2(n_38),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_51),
.B1(n_46),
.B2(n_39),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_61),
.B(n_29),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_47),
.A2(n_38),
.B1(n_28),
.B2(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_64),
.A3(n_18),
.B1(n_37),
.B2(n_30),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_97),
.B(n_107),
.C(n_20),
.D(n_12),
.Y(n_173)
);

NOR2x1_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_52),
.Y(n_120)
);

OAI21x1_ASAP7_75t_SL g178 ( 
.A1(n_120),
.A2(n_128),
.B(n_147),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_126),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_47),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_135),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_81),
.A2(n_53),
.B(n_32),
.C(n_8),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_77),
.B(n_90),
.C(n_10),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_73),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_141),
.C(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_53),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_67),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_58),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_67),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_53),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_110),
.A3(n_20),
.B1(n_111),
.B2(n_82),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_51),
.C(n_46),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_100),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_158),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_92),
.A2(n_46),
.B1(n_20),
.B2(n_39),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_154),
.B1(n_101),
.B2(n_110),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_74),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_115),
.B1(n_96),
.B2(n_104),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_74),
.A2(n_20),
.B1(n_39),
.B2(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_84),
.B(n_7),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_159),
.B(n_166),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_162),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_110),
.B(n_82),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_161),
.A2(n_165),
.B(n_176),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_168),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_164),
.B(n_138),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_101),
.B(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_84),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_189),
.B1(n_195),
.B2(n_144),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_174),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_173),
.B(n_118),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_122),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_102),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_146),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_142),
.B(n_157),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_102),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_193),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_96),
.B1(n_103),
.B2(n_104),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_156),
.B1(n_133),
.B2(n_121),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_103),
.B1(n_87),
.B2(n_7),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_87),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_132),
.B(n_6),
.C(n_11),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_128),
.A2(n_14),
.B1(n_10),
.B2(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_147),
.A3(n_157),
.B1(n_152),
.B2(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_212),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_198),
.A2(n_205),
.B1(n_206),
.B2(n_210),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

AOI22x1_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_152),
.B1(n_118),
.B2(n_148),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_213),
.B(n_214),
.Y(n_240)
);

NAND2x1_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_150),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_184),
.B(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_171),
.A2(n_143),
.B1(n_140),
.B2(n_155),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_188),
.B1(n_161),
.B2(n_167),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_226),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_133),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_182),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_149),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_167),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_192),
.B1(n_169),
.B2(n_131),
.Y(n_254)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_138),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_188),
.B1(n_165),
.B2(n_159),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_239),
.B1(n_241),
.B2(n_250),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_203),
.B(n_213),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_159),
.B1(n_190),
.B2(n_160),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_197),
.A2(n_189),
.B1(n_179),
.B2(n_175),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_164),
.B(n_170),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_253),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_179),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.C(n_251),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_252),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_173),
.B1(n_181),
.B2(n_174),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_181),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_244),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_172),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_202),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_206),
.B1(n_219),
.B2(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_220),
.Y(n_259)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_264),
.C(n_267),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_210),
.C(n_205),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_262),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_208),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_225),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_273),
.B(n_276),
.Y(n_287)
);

OA21x2_ASAP7_75t_SL g273 ( 
.A1(n_253),
.A2(n_220),
.B(n_217),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_208),
.C(n_214),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_239),
.C(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

BUFx12_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_241),
.B1(n_243),
.B2(n_235),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_285),
.B1(n_263),
.B2(n_269),
.Y(n_293)
);

AOI211xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_250),
.B(n_209),
.C(n_233),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_260),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_219),
.B1(n_233),
.B2(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_232),
.C(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_267),
.C(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_249),
.C(n_246),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_230),
.B(n_218),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_278),
.C(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_301),
.C(n_302),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_268),
.B1(n_258),
.B2(n_272),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_298),
.Y(n_309)
);

BUFx4f_ASAP7_75t_SL g298 ( 
.A(n_279),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_183),
.B(n_216),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_303),
.B1(n_277),
.B2(n_196),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_266),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_255),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_255),
.C(n_236),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_290),
.C(n_281),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_307),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_287),
.B(n_283),
.C(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_310),
.A2(n_296),
.B(n_1),
.C(n_3),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_194),
.B(n_238),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_298),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_192),
.C(n_215),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_222),
.A3(n_199),
.B1(n_169),
.B2(n_183),
.C1(n_186),
.C2(n_131),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_319),
.B1(n_306),
.B2(n_305),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_310),
.B1(n_308),
.B2(n_4),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_301),
.A3(n_302),
.B1(n_296),
.B2(n_186),
.C1(n_6),
.C2(n_5),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_0),
.C(n_1),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_323),
.B(n_325),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_317),
.Y(n_321)
);

OAI221xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_4),
.B1(n_324),
.B2(n_320),
.C(n_322),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_308),
.C(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_326),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);


endmodule