module fake_jpeg_29008_n_365 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_365);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_365;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_49),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_24),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_79),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_32),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_70),
.A2(n_28),
.B1(n_38),
.B2(n_35),
.Y(n_137)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_12),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_83),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_12),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_86),
.B(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx6f_ASAP7_75t_SL g150 ( 
.A(n_88),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_90),
.Y(n_129)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_92),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_25),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_31),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_39),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_45),
.B1(n_39),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_101),
.A2(n_112),
.B1(n_118),
.B2(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_135),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_103),
.B(n_121),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_45),
.B1(n_47),
.B2(n_46),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_53),
.A2(n_48),
.B1(n_47),
.B2(n_43),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_31),
.C(n_42),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_57),
.A2(n_30),
.B1(n_42),
.B2(n_38),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_97),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_74),
.A2(n_77),
.B1(n_68),
.B2(n_56),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_92),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_143),
.B1(n_8),
.B2(n_111),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_48),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_144),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_49),
.A2(n_19),
.B1(n_33),
.B2(n_28),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_140),
.A2(n_61),
.B1(n_54),
.B2(n_5),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_51),
.A2(n_35),
.B1(n_33),
.B2(n_25),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_23),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_82),
.A2(n_23),
.B(n_22),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_9),
.B(n_4),
.C(n_5),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_64),
.B1(n_65),
.B2(n_88),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_158),
.B1(n_159),
.B2(n_162),
.Y(n_213)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_104),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_160),
.Y(n_203)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_156),
.Y(n_200)
);

OR2x6_ASAP7_75t_SL g157 ( 
.A(n_113),
.B(n_97),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_175),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_89),
.B1(n_19),
.B2(n_22),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_61),
.B1(n_54),
.B2(n_21),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_165),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_147),
.B1(n_127),
.B2(n_145),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_105),
.B(n_100),
.Y(n_196)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_1),
.B(n_3),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_150),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_82),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_181),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_180),
.B(n_150),
.Y(n_210)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_179),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_124),
.B1(n_142),
.B2(n_128),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_113),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_129),
.B(n_109),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_149),
.B1(n_116),
.B2(n_108),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_130),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_108),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_148),
.C(n_117),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_205),
.C(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_105),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_161),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_196),
.B(n_158),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_148),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_212),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_126),
.C(n_119),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_126),
.C(n_149),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_171),
.Y(n_237)
);

BUFx24_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_110),
.B(n_115),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_166),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_128),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_165),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_219),
.Y(n_252)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_184),
.A3(n_180),
.B1(n_151),
.B2(n_183),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_238),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_240),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_156),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_164),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_153),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_211),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_173),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_183),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_241),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_190),
.B(n_116),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_205),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_220),
.C(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

CKINVDCx12_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_213),
.B1(n_208),
.B2(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_255),
.B(n_219),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_210),
.B(n_199),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_221),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_236),
.B(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_266),
.C(n_271),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_226),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_221),
.B(n_199),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_279),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_220),
.C(n_239),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_231),
.C(n_240),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_221),
.B(n_199),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_229),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_281),
.C(n_282),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_224),
.B(n_233),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_251),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_207),
.C(n_202),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_201),
.C(n_213),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_201),
.C(n_216),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_283),
.B(n_244),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_252),
.B1(n_254),
.B2(n_253),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_290),
.B1(n_295),
.B2(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_285),
.B(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_261),
.B1(n_257),
.B2(n_259),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_291),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_260),
.B1(n_212),
.B2(n_228),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_282),
.A2(n_225),
.B1(n_256),
.B2(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_283),
.B1(n_225),
.B2(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_299),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_260),
.B1(n_249),
.B2(n_243),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_306),
.B1(n_308),
.B2(n_313),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_266),
.C(n_277),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_309),
.C(n_312),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_267),
.B1(n_280),
.B2(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_269),
.B1(n_276),
.B2(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_223),
.C(n_222),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_250),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_262),
.C(n_200),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_194),
.B1(n_242),
.B2(n_262),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_250),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_297),
.A2(n_188),
.B(n_187),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_299),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_295),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_319),
.Y(n_336)
);

NAND2x1p5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_294),
.Y(n_317)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_294),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_286),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_322),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_289),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_297),
.C(n_291),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_314),
.C(n_301),
.Y(n_332)
);

AOI221xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_315),
.B1(n_302),
.B2(n_300),
.C(n_301),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_288),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_289),
.C(n_194),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_309),
.B(n_305),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_317),
.B(n_242),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_332),
.B(n_335),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_334),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_294),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_320),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_320),
.C(n_324),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_345),
.B(n_215),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_342),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_329),
.B1(n_328),
.B2(n_327),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_344),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_328),
.A2(n_334),
.B1(n_336),
.B2(n_188),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_214),
.C(n_217),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_217),
.C(n_214),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_349),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_351),
.Y(n_353)
);

AOI322xp5_ASAP7_75t_L g349 ( 
.A1(n_344),
.A2(n_191),
.A3(n_174),
.B1(n_181),
.B2(n_154),
.C1(n_215),
.C2(n_242),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_339),
.B(n_176),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_340),
.B(n_189),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_189),
.B(n_123),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_345),
.C(n_191),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_350),
.A2(n_186),
.B(n_179),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_349),
.C(n_100),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_136),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_360),
.C(n_356),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_361),
.A2(n_362),
.B(n_120),
.Y(n_363)
);

O2A1O1Ixp33_ASAP7_75t_SL g362 ( 
.A1(n_359),
.A2(n_353),
.B(n_136),
.C(n_120),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_142),
.C(n_130),
.Y(n_364)
);

BUFx24_ASAP7_75t_SL g365 ( 
.A(n_364),
.Y(n_365)
);


endmodule