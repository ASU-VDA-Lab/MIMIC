module fake_jpeg_6500_n_52 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_0),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_11),
.B(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_18),
.B(n_6),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_19),
.A2(n_7),
.B1(n_30),
.B2(n_29),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_16),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_28),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_33),
.B1(n_31),
.B2(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_42),
.B2(n_40),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_37),
.B1(n_41),
.B2(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

NAND2x1_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_42),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_48),
.C(n_47),
.Y(n_50)
);

A2O1A1O1Ixp25_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_43),
.B(n_40),
.C(n_23),
.D(n_27),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_16),
.B(n_27),
.Y(n_52)
);


endmodule