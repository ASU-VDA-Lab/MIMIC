module real_jpeg_29647_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_53),
.Y(n_74)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_1),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_5),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_22),
.B1(n_48),
.B2(n_52),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_SL g97 ( 
.A1(n_5),
.A2(n_28),
.B(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_5),
.B(n_123),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_6),
.B(n_48),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_8),
.B(n_31),
.C(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_48),
.B1(n_52),
.B2(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_9),
.A2(n_48),
.B1(n_52),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_10),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_102),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_100),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_85),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_85),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_76),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_45),
.B2(n_66),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_17),
.A2(n_18),
.B1(n_93),
.B2(n_94),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_33),
.B2(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_44),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_19),
.A2(n_20),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

AOI211xp5_ASAP7_75t_L g107 ( 
.A1(n_20),
.A2(n_58),
.B(n_84),
.C(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_22),
.A2(n_23),
.B(n_29),
.C(n_97),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_22),
.A2(n_39),
.B(n_61),
.C(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_22),
.B(n_60),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_146),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_22),
.A2(n_38),
.B(n_40),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_40),
.Y(n_42)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_33),
.A2(n_44),
.B1(n_58),
.B2(n_91),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_33),
.B(n_98),
.C(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_33),
.A2(n_44),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_43),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_35),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_39),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_91),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_44),
.A2(n_91),
.B(n_158),
.C(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_58),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_58),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_52),
.B(n_145),
.Y(n_144)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_80),
.B1(n_91),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_58),
.A2(n_91),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_91),
.B1(n_131),
.B2(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_58),
.B(n_98),
.C(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_58),
.A2(n_91),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_58),
.B(n_164),
.C(n_170),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_62),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_75),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B(n_83),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_84),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.C(n_92),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_92),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_99),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_98),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_98),
.A2(n_99),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_98),
.A2(n_99),
.B1(n_121),
.B2(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_124),
.B(n_181),
.C(n_186),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_104),
.B(n_113),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_112),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_182)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_120),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_114),
.A2(n_115),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_117),
.B1(n_154),
.B2(n_158),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_180),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_173),
.B(n_179),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_160),
.B(n_172),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_151),
.B(n_159),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_139),
.B(n_150),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);


endmodule