module fake_jpeg_32131_n_118 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_45),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_17),
.B(n_25),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_35),
.C(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_17),
.B1(n_13),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_13),
.B1(n_20),
.B2(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_39),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_31),
.B1(n_20),
.B2(n_15),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_17),
.B(n_22),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_3),
.B(n_25),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_61),
.C(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_27),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_28),
.C(n_32),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_64),
.B1(n_24),
.B2(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_26),
.B1(n_24),
.B2(n_19),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_71),
.B1(n_78),
.B2(n_80),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_75),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_27),
.B(n_18),
.C(n_38),
.Y(n_68)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_50),
.B(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_53),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_18),
.B1(n_3),
.B2(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_83),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_67),
.B1(n_63),
.B2(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_96),
.B1(n_90),
.B2(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_71),
.B1(n_77),
.B2(n_75),
.Y(n_96)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_78),
.B(n_70),
.C(n_55),
.D(n_79),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_82),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_86),
.B(n_87),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_99),
.B(n_100),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_82),
.B(n_86),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_93),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_60),
.C(n_65),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_106),
.C(n_96),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_5),
.C(n_9),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_109),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_102),
.B(n_97),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_94),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_113),
.A2(n_114),
.B(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_112),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);


endmodule