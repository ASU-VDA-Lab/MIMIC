module fake_jpeg_11893_n_245 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_13),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_32),
.B1(n_37),
.B2(n_34),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_66),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_85),
.B1(n_95),
.B2(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_80),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_28),
.B1(n_34),
.B2(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_27),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_24),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_39),
.B1(n_30),
.B2(n_29),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_111),
.B1(n_125),
.B2(n_82),
.Y(n_149)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_61),
.B1(n_57),
.B2(n_62),
.Y(n_108)
);

OAI22x1_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_85),
.B1(n_48),
.B2(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_66),
.A2(n_63),
.B1(n_49),
.B2(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_118),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_20),
.B(n_30),
.C(n_29),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_106),
.A3(n_104),
.B1(n_114),
.B2(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_27),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_117),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_122),
.Y(n_131)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_23),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_23),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_20),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_107),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_118),
.B1(n_103),
.B2(n_70),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_73),
.B1(n_89),
.B2(n_65),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_146),
.B1(n_143),
.B2(n_136),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_77),
.C(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_143),
.C(n_133),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_82),
.B(n_92),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_89),
.C(n_73),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_121),
.B1(n_113),
.B2(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_96),
.B1(n_70),
.B2(n_65),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_101),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_138),
.C(n_140),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_154),
.C(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_117),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_135),
.B1(n_148),
.B2(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_99),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_166),
.B1(n_171),
.B2(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_168),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_130),
.A2(n_24),
.B1(n_6),
.B2(n_7),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_4),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_4),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_129),
.B1(n_144),
.B2(n_147),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_180),
.B(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_128),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_185),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_139),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_164),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_137),
.B1(n_148),
.B2(n_149),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_139),
.B(n_7),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_6),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_159),
.B1(n_170),
.B2(n_144),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_147),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_160),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_203),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_180),
.B(n_167),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_206),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_178),
.B(n_188),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_6),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_178),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_210),
.B(n_211),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_174),
.B(n_186),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_177),
.B(n_181),
.C(n_192),
.D(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_195),
.C(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_226),
.C(n_216),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_207),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_214),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_218),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_222),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_205),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_224),
.B(n_213),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_201),
.C(n_190),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_196),
.B(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_8),
.B(n_9),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_228),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_190),
.B1(n_191),
.B2(n_175),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_233),
.B1(n_223),
.B2(n_220),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_221),
.B1(n_9),
.B2(n_11),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_238),
.B(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_234),
.B(n_232),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_243),
.Y(n_245)
);


endmodule