module fake_jpeg_13764_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_75),
.Y(n_87)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_0),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_85),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_47),
.B1(n_49),
.B2(n_54),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_90),
.B(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_48),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_91),
.C(n_86),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_106),
.B(n_111),
.C(n_0),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_103),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_65),
.A3(n_62),
.B1(n_61),
.B2(n_51),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_35),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_53),
.B1(n_42),
.B2(n_3),
.Y(n_121)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_112),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_51),
.B(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_129),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_55),
.B1(n_60),
.B2(n_57),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_9),
.B(n_13),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_128),
.B1(n_117),
.B2(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_30),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_27),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_124),
.C(n_125),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_7),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_15),
.Y(n_145)
);

OR2x6_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_8),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_40),
.B(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_140),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_141),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_147),
.B(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_145),
.B(n_146),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_26),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_145),
.B(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_144),
.B1(n_131),
.B2(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_139),
.C(n_142),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_149),
.B(n_148),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_148),
.B(n_156),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_151),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_31),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_34),
.Y(n_163)
);


endmodule