module real_jpeg_4524_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_1),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_1),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_1),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_1),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_1),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_1),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_1),
.B(n_328),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_2),
.Y(n_98)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_2),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_2),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_2),
.Y(n_309)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_2),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_2),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_3),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_3),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_3),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_3),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_3),
.B(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_5),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_5),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_5),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_5),
.B(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_7),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_11),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_11),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_11),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_11),
.B(n_72),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_11),
.Y(n_432)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_12),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_13),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_13),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_13),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_13),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_14),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_14),
.B(n_143),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_14),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_14),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_14),
.B(n_488),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_15),
.Y(n_126)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_15),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_16),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_16),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_16),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_17),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_17),
.B(n_113),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_17),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_17),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_17),
.B(n_72),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_17),
.B(n_97),
.Y(n_470)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_499),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_478),
.B(n_498),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_423),
.B(n_475),
.Y(n_26)
);

AO21x2_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_277),
.B(n_311),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_234),
.B(n_276),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_206),
.B(n_233),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_30),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_166),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_31),
.B(n_166),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_109),
.C(n_150),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_32),
.B(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_32),
.Y(n_516)
);

FAx1_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_74),
.CI(n_91),
.CON(n_32),
.SN(n_32)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_33),
.B(n_74),
.C(n_91),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_50),
.C(n_64),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_34),
.B(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_45),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_36),
.B(n_41),
.C(n_45),
.Y(n_165)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_39),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_40),
.Y(n_358)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_49),
.Y(n_164)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_49),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_49),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_50),
.A2(n_64),
.B1(n_65),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_50),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_61),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_51),
.A2(n_61),
.B1(n_185),
.B2(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_51),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_51),
.A2(n_215),
.B1(n_224),
.B2(n_257),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_51),
.A2(n_111),
.B1(n_112),
.B2(n_215),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_51),
.B(n_224),
.C(n_283),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_77),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_52),
.B(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_52),
.B(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_55),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_61),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_61),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_61),
.B(n_186),
.C(n_190),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_62),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_63),
.Y(n_226)
);

BUFx8_ASAP7_75t_L g383 ( 
.A(n_63),
.Y(n_383)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_227)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_69),
.Y(n_375)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_73),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_75),
.A2(n_76),
.B1(n_111),
.B2(n_112),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_75),
.B(n_112),
.C(n_470),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_75),
.A2(n_76),
.B1(n_173),
.B2(n_174),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_75),
.B(n_174),
.C(n_296),
.Y(n_505)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_76),
.B(n_83),
.C(n_88),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_79),
.Y(n_244)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_79),
.Y(n_337)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_83),
.A2(n_90),
.B1(n_134),
.B2(n_135),
.Y(n_343)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_100),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_93),
.B(n_95),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_92),
.B(n_101),
.C(n_104),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_99),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_105),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_105),
.B(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_105),
.B(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_108),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_109),
.B(n_150),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_129),
.C(n_131),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_110),
.A2(n_129),
.B1(n_130),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_128),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_117),
.C(n_122),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_112),
.B(n_215),
.C(n_447),
.Y(n_467)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_121),
.A2(n_122),
.B1(n_242),
.B2(n_249),
.Y(n_241)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_122),
.B(n_243),
.C(n_245),
.Y(n_289)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_126),
.Y(n_366)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_131),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.C(n_145),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_132),
.A2(n_133),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_139),
.A2(n_140),
.B1(n_145),
.B2(n_146),
.Y(n_411)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_165),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_153),
.C(n_165),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_156),
.C(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_155),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_155),
.Y(n_295)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_164),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_167),
.B(n_169),
.C(n_205),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_192),
.B1(n_204),
.B2(n_205),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_182),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_171),
.B(n_172),
.C(n_182),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_181),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_173),
.A2(n_174),
.B1(n_253),
.B2(n_254),
.Y(n_507)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_174),
.B(n_273),
.C(n_274),
.Y(n_272)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_179),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_189),
.B2(n_190),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_186),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_186),
.A2(n_188),
.B1(n_224),
.B2(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_186),
.B(n_224),
.C(n_254),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_186),
.A2(n_188),
.B1(n_334),
.B2(n_335),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_188),
.B(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_189),
.A2(n_190),
.B1(n_435),
.B2(n_439),
.Y(n_434)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_190),
.B(n_430),
.C(n_435),
.Y(n_465)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_202),
.C(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_231),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_207),
.B(n_231),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_228),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_208),
.A2(n_209),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_212),
.B(n_228),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.C(n_227),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_213),
.B(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_216),
.B(n_227),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_224),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_331)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_220),
.Y(n_328)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_224),
.A2(n_257),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_235),
.B(n_277),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_278),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_237),
.B(n_278),
.Y(n_422)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_259),
.CI(n_275),
.CON(n_237),
.SN(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_252),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_250),
.B2(n_251),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_240),
.B(n_251),
.C(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_248),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_258),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_262),
.C(n_264),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_265)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_270),
.C(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_271),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_268),
.A2(n_271),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_268),
.B(n_461),
.C(n_465),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_271),
.B(n_305),
.C(n_308),
.Y(n_428)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_279),
.B(n_281),
.C(n_298),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_298),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_282),
.B(n_289),
.C(n_290),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_296),
.B2(n_297),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_452)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_296),
.A2(n_297),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_310),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_299),
.B(n_302),
.C(n_304),
.Y(n_453)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

OAI31xp33_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_419),
.A3(n_420),
.B(n_422),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_413),
.B(n_418),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_398),
.B(n_412),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_353),
.B(n_397),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_344),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_344),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_332),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_329),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_318),
.B(n_329),
.C(n_332),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.C(n_326),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_346)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_326),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_333),
.B(n_407),
.C(n_408),
.Y(n_406)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.C(n_352),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_352),
.B1(n_389),
.B2(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_349),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_391),
.B(n_396),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_377),
.B(n_390),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_362),
.B(n_376),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_372),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_372),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_367),
.B(n_371),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_367),
.Y(n_371)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_379),
.B1(n_384),
.B2(n_385),
.Y(n_378)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_386),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_386),
.Y(n_390)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_379),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_380),
.A2(n_381),
.B(n_384),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_388),
.B(n_389),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_393),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_400),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_404),
.B2(n_405),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_406),
.C(n_409),
.Y(n_414)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_415),
.Y(n_418)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_416),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_472),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_424),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_454),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_454),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_444),
.C(n_453),
.Y(n_425)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_426),
.B(n_444),
.CI(n_453),
.CON(n_474),
.SN(n_474)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_426)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_429),
.C(n_443),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_433),
.B1(n_434),
.B2(n_440),
.Y(n_429)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_430),
.A2(n_440),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_449),
.B2(n_450),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_451),
.C(n_452),
.Y(n_456)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_454),
.Y(n_513)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_456),
.CI(n_457),
.CON(n_454),
.SN(n_454)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_455),
.B(n_456),
.C(n_457),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_466),
.B2(n_471),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_458),
.B(n_467),
.C(n_468),
.Y(n_496)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_465),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_462),
.Y(n_461)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_466),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_473),
.B(n_474),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_474),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_497),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_497),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_496),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_483),
.C(n_496),
.Y(n_511)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_492),
.B2(n_493),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_487),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_489),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_490),
.C(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_495),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_512),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_511),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_511),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_509),
.B2(n_510),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_505),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_506),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_507),
.Y(n_508)
);


endmodule