module real_aes_9945_n_5 (n_4, n_0, n_3, n_2, n_1, n_5);
input n_4;
input n_0;
input n_3;
input n_2;
input n_1;
output n_5;
wire n_17;
wire n_13;
wire n_6;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_18;
wire n_7;
wire n_8;
wire n_10;
OAI21xp33_ASAP7_75t_SL g6 ( .A1(n_0), .A2(n_1), .B(n_7), .Y(n_6) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_1), .A2(n_13), .B(n_14), .Y(n_12) );
AOI22xp33_ASAP7_75t_L g5 ( .A1(n_2), .A2(n_6), .B1(n_15), .B2(n_19), .Y(n_5) );
INVx1_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_11), .Y(n_14) );
BUFx2_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_11), .B(n_12), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_9), .Y(n_8) );
BUFx8_ASAP7_75t_SL g9 ( .A(n_10), .Y(n_9) );
INVx4_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
NOR3xp33_ASAP7_75t_L g15 ( .A(n_16), .B(n_17), .C(n_18), .Y(n_15) );
endmodule