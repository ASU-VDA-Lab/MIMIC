module fake_jpeg_20629_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_149;
wire n_35;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_36),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_43),
.B1(n_39),
.B2(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_25),
.B1(n_33),
.B2(n_31),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_72),
.B1(n_81),
.B2(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_77),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_67),
.B(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_25),
.B1(n_43),
.B2(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_86),
.B1(n_92),
.B2(n_98),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_28),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_78),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_37),
.B(n_23),
.Y(n_130)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_18),
.B1(n_27),
.B2(n_36),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_43),
.B1(n_44),
.B2(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_43),
.B1(n_30),
.B2(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_96),
.B1(n_40),
.B2(n_39),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_45),
.B1(n_37),
.B2(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_45),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_99),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_39),
.B1(n_40),
.B2(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_29),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_40),
.B1(n_45),
.B2(n_37),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_20),
.B(n_29),
.C(n_45),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_131),
.B1(n_133),
.B2(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_122),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_130),
.B(n_102),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_20),
.B(n_23),
.C(n_22),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_85),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_37),
.B1(n_21),
.B2(n_19),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_69),
.A2(n_21),
.B1(n_19),
.B2(n_37),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_92),
.B1(n_76),
.B2(n_84),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_136),
.A2(n_151),
.B1(n_162),
.B2(n_109),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_95),
.C(n_79),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_132),
.C(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_148),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_164),
.B(n_119),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_79),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_150),
.B(n_155),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_79),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_103),
.B1(n_96),
.B2(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_91),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_91),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_88),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_125),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_80),
.B(n_87),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_68),
.B1(n_71),
.B2(n_89),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_89),
.B1(n_88),
.B2(n_21),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_131),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_35),
.Y(n_164)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_107),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_167),
.B(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_175),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_185),
.C(n_137),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_109),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_177),
.B(n_181),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_142),
.B(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_186),
.B1(n_142),
.B2(n_164),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_111),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_115),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_115),
.C(n_125),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_110),
.B1(n_112),
.B2(n_126),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_120),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_190),
.B(n_191),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_146),
.B(n_150),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_120),
.B(n_123),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_211),
.C(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_205),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_171),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_151),
.B1(n_163),
.B2(n_159),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_139),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_143),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_145),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_159),
.C(n_144),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_117),
.B1(n_120),
.B2(n_87),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_165),
.A2(n_117),
.B1(n_35),
.B2(n_26),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_192),
.B1(n_179),
.B2(n_170),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_35),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_180),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_26),
.C(n_16),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_26),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_188),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_191),
.B(n_174),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_227),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_218),
.Y(n_243)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_233),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_174),
.B(n_189),
.Y(n_233)
);

AOI211xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_165),
.B(n_189),
.C(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_193),
.C(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_193),
.C(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_237),
.A2(n_205),
.B1(n_198),
.B2(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_192),
.C(n_16),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_194),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_244),
.B1(n_232),
.B2(n_223),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_213),
.B1(n_212),
.B2(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_222),
.B1(n_219),
.B2(n_221),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_248),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_226),
.A2(n_209),
.B1(n_202),
.B2(n_211),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_217),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_253),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_195),
.B1(n_216),
.B2(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_215),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_207),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_194),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.C(n_228),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_214),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_261),
.B1(n_267),
.B2(n_242),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_265),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_241),
.A2(n_219),
.B(n_231),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_266),
.B(n_6),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_234),
.B1(n_1),
.B2(n_2),
.Y(n_261)
);

AO22x1_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_0),
.C(n_3),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_4),
.B(n_5),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_254),
.B(n_243),
.C(n_247),
.D(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_276),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_278),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_6),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_10),
.B(n_11),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_267),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_7),
.B(n_9),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_270),
.Y(n_286)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_274),
.A3(n_267),
.B1(n_262),
.B2(n_257),
.C1(n_15),
.C2(n_13),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_268),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_280),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_288),
.B(n_280),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_284),
.B(n_262),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_292),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_281),
.B(n_12),
.Y(n_299)
);


endmodule