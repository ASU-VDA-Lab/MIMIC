module fake_jpeg_31446_n_553 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_553);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_18),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_17),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_54),
.B(n_91),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_55),
.B(n_90),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_56),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_17),
.B1(n_16),
.B2(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_63),
.A2(n_23),
.B1(n_24),
.B2(n_49),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_72),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_22),
.B(n_16),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_74),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_82),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_77),
.Y(n_135)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx11_ASAP7_75t_SL g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_89),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_0),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_0),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_103),
.Y(n_120)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_40),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_23),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_108),
.B(n_124),
.Y(n_189)
);

NAND2x1_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_40),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_122),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_24),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_126),
.B(n_138),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_67),
.A2(n_53),
.B1(n_39),
.B2(n_42),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_53),
.B1(n_39),
.B2(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_21),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_25),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_59),
.B(n_25),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_30),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_63),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_104),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_68),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_56),
.B(n_30),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_32),
.Y(n_162)
);

BUFx16f_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_109),
.B(n_48),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_171),
.B(n_197),
.C(n_211),
.Y(n_269)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_105),
.B1(n_80),
.B2(n_95),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_174),
.A2(n_223),
.B1(n_159),
.B2(n_19),
.Y(n_272)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_107),
.B1(n_93),
.B2(n_61),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_178),
.A2(n_204),
.B1(n_0),
.B2(n_2),
.Y(n_274)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_181),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_195),
.Y(n_252)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_115),
.B(n_32),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_114),
.A2(n_35),
.B(n_36),
.C(n_51),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_196),
.B(n_215),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_48),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_198),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_130),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_199),
.B(n_231),
.Y(n_275)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_203),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_120),
.B(n_49),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_154),
.A2(n_65),
.B1(n_66),
.B2(n_75),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_70),
.B1(n_69),
.B2(n_40),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_205),
.A2(n_127),
.B1(n_156),
.B2(n_128),
.Y(n_247)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

CKINVDCx12_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_208),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_144),
.B(n_35),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_210),
.B(n_216),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_110),
.B(n_51),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_36),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_218),
.Y(n_270)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_220),
.B1(n_229),
.B2(n_230),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_222),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_117),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_123),
.A2(n_101),
.B1(n_79),
.B2(n_62),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_125),
.B(n_99),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_227),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_157),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_125),
.B(n_19),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_153),
.Y(n_235)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_129),
.Y(n_229)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_81),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_259),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_196),
.A2(n_168),
.B1(n_116),
.B2(n_142),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_236),
.A2(n_247),
.B1(n_254),
.B2(n_255),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_116),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_163),
.C(n_143),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_248),
.Y(n_285)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_153),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_180),
.A2(n_168),
.B1(n_142),
.B2(n_113),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_250),
.A2(n_266),
.B1(n_205),
.B2(n_192),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_134),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_186),
.A2(n_134),
.B1(n_118),
.B2(n_131),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_186),
.A2(n_131),
.B1(n_118),
.B2(n_148),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_148),
.B1(n_121),
.B2(n_71),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_181),
.A2(n_135),
.B1(n_121),
.B2(n_143),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_199),
.B(n_213),
.C(n_188),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_261),
.B(n_248),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_174),
.A2(n_129),
.B1(n_19),
.B2(n_152),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_272),
.A2(n_274),
.B1(n_176),
.B2(n_219),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_218),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_189),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_296),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_222),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_287),
.B(n_292),
.Y(n_363)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_178),
.B(n_204),
.C(n_221),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_289),
.A2(n_251),
.B(n_233),
.Y(n_349)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_184),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_192),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_295),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_294),
.A2(n_274),
.B1(n_246),
.B2(n_271),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_183),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_216),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_256),
.B(n_198),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_298),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_230),
.B(n_173),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_301),
.B(n_243),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_208),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_198),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_202),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_308),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_273),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_306),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_202),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_309),
.A2(n_240),
.B1(n_257),
.B2(n_271),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_261),
.B(n_237),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_276),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_311),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_208),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_244),
.C(n_248),
.Y(n_329)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_229),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_318),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_232),
.B(n_217),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_316),
.Y(n_364)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_232),
.B(n_209),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_320),
.Y(n_354)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_238),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_259),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_269),
.B(n_191),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_323),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_237),
.B(n_194),
.Y(n_323)
);

INVx4_ASAP7_75t_SL g324 ( 
.A(n_278),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_324),
.A2(n_271),
.B1(n_279),
.B2(n_243),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_330),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_247),
.C(n_255),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_254),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_332),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_258),
.C(n_264),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_333),
.B(n_357),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_284),
.A2(n_272),
.B(n_270),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_336),
.A2(n_337),
.B(n_342),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_284),
.A2(n_262),
.B(n_259),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_308),
.B1(n_315),
.B2(n_303),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_284),
.A2(n_182),
.B1(n_264),
.B2(n_258),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_343),
.A2(n_359),
.B1(n_297),
.B2(n_317),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_349),
.B1(n_355),
.B2(n_289),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_296),
.B1(n_286),
.B2(n_299),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_251),
.C(n_239),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_220),
.B1(n_240),
.B2(n_265),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_361),
.B1(n_294),
.B2(n_324),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_281),
.A2(n_240),
.B1(n_265),
.B2(n_239),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_354),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_382),
.Y(n_400)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_311),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_369),
.Y(n_419)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_306),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_372),
.B(n_379),
.Y(n_402)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_385),
.B1(n_389),
.B2(n_360),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_305),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_281),
.Y(n_380)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_326),
.B(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_335),
.Y(n_382)
);

INVx13_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_387),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_290),
.Y(n_384)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_283),
.B1(n_303),
.B2(n_291),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_334),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_393),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_328),
.B(n_301),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_392),
.B(n_395),
.Y(n_418)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_345),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_396),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_352),
.B(n_282),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

AOI21xp33_ASAP7_75t_L g427 ( 
.A1(n_397),
.A2(n_398),
.B(n_341),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_391),
.B(n_352),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_398),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_378),
.B(n_329),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_406),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_333),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_331),
.C(n_357),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_412),
.C(n_431),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_411),
.A2(n_339),
.B1(n_384),
.B2(n_381),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_330),
.C(n_332),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_342),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_397),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_336),
.B1(n_337),
.B2(n_353),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_422),
.A2(n_428),
.B1(n_368),
.B2(n_371),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_427),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_353),
.B1(n_349),
.B2(n_283),
.Y(n_428)
);

AOI221xp5_ASAP7_75t_L g429 ( 
.A1(n_382),
.A2(n_358),
.B1(n_365),
.B2(n_388),
.C(n_387),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_388),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_364),
.C(n_343),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_436),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_434),
.B(n_451),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_380),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_439),
.C(n_446),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_408),
.A2(n_389),
.B1(n_367),
.B2(n_374),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_408),
.A2(n_359),
.B1(n_364),
.B2(n_377),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_441),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_448),
.B1(n_454),
.B2(n_456),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_358),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_363),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_418),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_445),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_366),
.Y(n_443)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_282),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_396),
.C(n_393),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_282),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_449),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_327),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_450),
.A2(n_458),
.B(n_417),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_403),
.B(n_362),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_455),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_373),
.B1(n_370),
.B2(n_325),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_362),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_423),
.A2(n_356),
.B1(n_325),
.B2(n_344),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_411),
.A2(n_422),
.B1(n_428),
.B2(n_415),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_421),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_426),
.A2(n_356),
.B1(n_344),
.B2(n_288),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_415),
.A2(n_409),
.B(n_430),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_459),
.A2(n_443),
.B(n_448),
.Y(n_471)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_464),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_452),
.Y(n_467)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_467),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_431),
.C(n_409),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_470),
.C(n_476),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_430),
.C(n_426),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_454),
.B(n_456),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_474),
.A2(n_457),
.B1(n_434),
.B2(n_451),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_432),
.B(n_421),
.C(n_424),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_459),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_424),
.C(n_417),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_481),
.C(n_482),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_413),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_444),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_413),
.C(n_407),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_439),
.B(n_407),
.C(n_268),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_483),
.B(n_488),
.Y(n_515)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_475),
.Y(n_485)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_485),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_471),
.A2(n_436),
.B(n_437),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_487),
.A2(n_498),
.B(n_460),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_473),
.B(n_455),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_493),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_472),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_480),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_468),
.A2(n_405),
.B1(n_314),
.B2(n_307),
.Y(n_494)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_468),
.Y(n_495)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_499),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_461),
.C(n_470),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_478),
.C(n_469),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_462),
.A2(n_383),
.B(n_405),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_486),
.B(n_465),
.Y(n_501)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_501),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_502),
.B(n_504),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_514),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_487),
.A2(n_460),
.B(n_481),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_510),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_461),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_508),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_500),
.A2(n_482),
.B(n_466),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_479),
.C(n_466),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_513),
.C(n_492),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_472),
.C(n_320),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_313),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_516),
.A2(n_484),
.B1(n_495),
.B2(n_485),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_521),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_518),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_524),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_494),
.B1(n_499),
.B2(n_498),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_SL g522 ( 
.A1(n_512),
.A2(n_483),
.B(n_491),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_522),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_515),
.A2(n_279),
.B1(n_234),
.B2(n_6),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_506),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_529),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_504),
.A2(n_234),
.B1(n_7),
.B2(n_8),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_505),
.Y(n_530)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_502),
.B1(n_511),
.B2(n_513),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_520),
.C(n_519),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_514),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_536),
.B(n_537),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_SL g537 ( 
.A(n_525),
.B(n_515),
.C(n_503),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_538),
.A2(n_524),
.B(n_522),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_541),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_533),
.A2(n_528),
.B(n_11),
.Y(n_542)
);

AOI21xp33_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_535),
.B(n_534),
.Y(n_544)
);

OAI21xp33_ASAP7_75t_L g548 ( 
.A1(n_544),
.A2(n_546),
.B(n_543),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_SL g546 ( 
.A(n_540),
.B(n_537),
.C(n_532),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_545),
.B(n_532),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_547),
.A2(n_548),
.B(n_9),
.Y(n_549)
);

AOI322xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_548),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_9),
.B(n_12),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_9),
.C(n_12),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_552),
.B(n_13),
.Y(n_553)
);


endmodule