module fake_jpeg_12659_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_62),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_29),
.B(n_10),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_68),
.Y(n_136)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_73),
.Y(n_199)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_76),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_77),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_29),
.B(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_82),
.B(n_86),
.Y(n_149)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_9),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_128),
.Y(n_154)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_37),
.B(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_92),
.B(n_105),
.Y(n_166)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_93),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_95),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_98),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_103),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_104),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_42),
.B(n_9),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_9),
.B(n_2),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_28),
.C(n_53),
.Y(n_184)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_42),
.B(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_120),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_20),
.B(n_25),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_123),
.Y(n_147)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

CKINVDCx6p67_ASAP7_75t_R g215 ( 
.A(n_117),
.Y(n_215)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_118),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_49),
.B(n_11),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_25),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_126),
.B(n_58),
.Y(n_217)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_11),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_18),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_130),
.B(n_15),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_44),
.B1(n_34),
.B2(n_40),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_137),
.A2(n_139),
.B1(n_179),
.B2(n_191),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_34),
.B1(n_40),
.B2(n_46),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_138),
.A2(n_172),
.B1(n_35),
.B2(n_38),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_73),
.A2(n_34),
.B1(n_40),
.B2(n_46),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_46),
.B1(n_54),
.B2(n_26),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_145),
.A2(n_41),
.B1(n_35),
.B2(n_125),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_54),
.B1(n_46),
.B2(n_57),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_161),
.A2(n_189),
.B1(n_213),
.B2(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_26),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_168),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_94),
.B(n_50),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_80),
.B(n_50),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_181),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_54),
.B1(n_59),
.B2(n_28),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_66),
.A2(n_54),
.B1(n_59),
.B2(n_33),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_39),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_184),
.B(n_217),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_77),
.A2(n_28),
.B1(n_53),
.B2(n_52),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_118),
.B(n_39),
.C(n_33),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_212),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_91),
.A2(n_59),
.B1(n_33),
.B2(n_53),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_127),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_122),
.Y(n_249)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_60),
.B(n_52),
.C(n_51),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_63),
.A2(n_58),
.B1(n_35),
.B2(n_51),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_81),
.A2(n_52),
.B1(n_51),
.B2(n_48),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_107),
.B(n_48),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_223),
.Y(n_344)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_226),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_228),
.Y(n_346)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_234),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_238),
.B(n_246),
.Y(n_333)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_147),
.A2(n_90),
.B(n_71),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_244),
.A2(n_163),
.B(n_152),
.Y(n_348)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_247),
.B(n_248),
.Y(n_350)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_215),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_250),
.Y(n_309)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_70),
.B1(n_76),
.B2(n_119),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_253),
.A2(n_298),
.B1(n_141),
.B2(n_144),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_136),
.B(n_126),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_254),
.B(n_258),
.Y(n_341)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_138),
.A2(n_104),
.B1(n_84),
.B2(n_113),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_257),
.A2(n_269),
.B1(n_276),
.B2(n_203),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_154),
.B(n_122),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_149),
.B(n_48),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_264),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_140),
.A2(n_41),
.B(n_38),
.C(n_58),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_260),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_354)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_261),
.B(n_275),
.Y(n_356)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_262),
.Y(n_353)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_166),
.B(n_38),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_186),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_274),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_164),
.Y(n_267)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_270),
.Y(n_323)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_156),
.Y(n_271)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_151),
.Y(n_272)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_287),
.B1(n_292),
.B2(n_293),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_188),
.B(n_41),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_139),
.A2(n_111),
.B1(n_110),
.B2(n_103),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_148),
.B(n_12),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_277),
.B(n_281),
.Y(n_355)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_155),
.B(n_193),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_132),
.Y(n_282)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_282),
.Y(n_332)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_165),
.Y(n_283)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_177),
.B(n_0),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_290),
.Y(n_300)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_180),
.Y(n_285)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_197),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_286),
.B(n_288),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_198),
.B(n_12),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_205),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_160),
.B(n_12),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_146),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_291),
.Y(n_334)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_208),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_199),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_172),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_187),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g295 ( 
.A(n_199),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_202),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_194),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_221),
.A2(n_99),
.B1(n_62),
.B2(n_3),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_171),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g308 ( 
.A1(n_232),
.A2(n_135),
.B1(n_179),
.B2(n_137),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_308),
.A2(n_326),
.B(n_348),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_233),
.A2(n_191),
.B1(n_160),
.B2(n_187),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_311),
.A2(n_359),
.B1(n_292),
.B2(n_295),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_284),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_276),
.A2(n_135),
.B1(n_131),
.B2(n_150),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_221),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_335),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_322),
.A2(n_345),
.B1(n_352),
.B2(n_357),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_SL g326 ( 
.A(n_255),
.B(n_215),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_230),
.B(n_205),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_233),
.A2(n_194),
.B1(n_144),
.B2(n_141),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_336),
.A2(n_342),
.B1(n_347),
.B2(n_287),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_244),
.A2(n_203),
.B(n_208),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_337),
.A2(n_278),
.B(n_251),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_229),
.B(n_163),
.CI(n_196),
.CON(n_339),
.SN(n_339)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_227),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_257),
.A2(n_185),
.B1(n_206),
.B2(n_157),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_265),
.A2(n_185),
.B1(n_206),
.B2(n_157),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_278),
.A2(n_152),
.B1(n_142),
.B2(n_216),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_0),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_273),
.A2(n_142),
.B1(n_4),
.B2(n_5),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_253),
.A2(n_265),
.B1(n_260),
.B2(n_273),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_360),
.A2(n_363),
.B(n_374),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_361),
.B(n_390),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_300),
.B(n_284),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_350),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_376),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_235),
.C(n_222),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_368),
.B(n_371),
.C(n_394),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_224),
.B1(n_289),
.B2(n_268),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_369),
.Y(n_424)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_370),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_243),
.C(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_349),
.Y(n_372)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_322),
.A2(n_298),
.B1(n_297),
.B2(n_286),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_330),
.B1(n_329),
.B2(n_332),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_310),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_350),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_383),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_300),
.B(n_285),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_323),
.B(n_237),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_341),
.C(n_356),
.Y(n_413)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_239),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_382),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_333),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_252),
.B1(n_262),
.B2(n_283),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_384),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_385),
.A2(n_386),
.B1(n_400),
.B2(n_402),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_342),
.A2(n_245),
.B1(n_280),
.B2(n_236),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_238),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_396),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_309),
.A2(n_308),
.B1(n_317),
.B2(n_314),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_388),
.A2(n_395),
.B(n_313),
.Y(n_426)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_267),
.C(n_226),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_309),
.A2(n_228),
.B1(n_293),
.B2(n_234),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_271),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_324),
.B(n_291),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_399),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_231),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_270),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_334),
.C(n_332),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_308),
.A2(n_250),
.B1(n_295),
.B2(n_6),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_301),
.Y(n_403)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_323),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_348),
.A2(n_13),
.B1(n_4),
.B2(n_6),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_405),
.A2(n_316),
.B1(n_305),
.B2(n_314),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_341),
.A2(n_223),
.B1(n_8),
.B2(n_12),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_406),
.A2(n_374),
.B(n_399),
.Y(n_414)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_363),
.C(n_398),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_414),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_339),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_419),
.B(n_420),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_379),
.Y(n_420)
);

MAJx2_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_337),
.C(n_339),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_362),
.C(n_380),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_365),
.B(n_356),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_429),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_383),
.B(n_352),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_396),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_422),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_394),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_392),
.A2(n_314),
.B1(n_329),
.B2(n_334),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_436),
.A2(n_385),
.B1(n_402),
.B2(n_386),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_368),
.B(n_304),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_325),
.C(n_351),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_438),
.A2(n_445),
.B1(n_373),
.B2(n_393),
.Y(n_469)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_439),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_371),
.B(n_325),
.C(n_328),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_360),
.C(n_401),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_400),
.A2(n_305),
.B1(n_304),
.B2(n_328),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_407),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_446),
.B(n_447),
.C(n_448),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_380),
.Y(n_448)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_423),
.C(n_422),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_439),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_450),
.B(n_455),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_378),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_452),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_453),
.A2(n_458),
.B1(n_416),
.B2(n_430),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_361),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_463),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_409),
.A2(n_366),
.B(n_361),
.Y(n_457)
);

AO21x1_ASAP7_75t_L g492 ( 
.A1(n_457),
.A2(n_461),
.B(n_467),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_409),
.A2(n_405),
.B1(n_392),
.B2(n_390),
.Y(n_458)
);

AO21x1_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_391),
.B(n_389),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_439),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_460),
.B(n_462),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_410),
.A2(n_406),
.B(n_367),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_412),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_428),
.B(n_377),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_410),
.B(n_375),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_469),
.B1(n_475),
.B2(n_436),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_414),
.A2(n_364),
.B(n_370),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_417),
.B(n_420),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_472),
.B(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_408),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_416),
.A2(n_372),
.B1(n_397),
.B2(n_381),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_408),
.Y(n_478)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_411),
.Y(n_479)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_479),
.Y(n_504)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_435),
.Y(n_486)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_476),
.Y(n_482)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_484),
.A2(n_453),
.B1(n_454),
.B2(n_457),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_511),
.Y(n_524)
);

XNOR2x1_ASAP7_75t_L g528 ( 
.A(n_489),
.B(n_441),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_490),
.A2(n_469),
.B1(n_477),
.B2(n_463),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_466),
.A2(n_445),
.B1(n_438),
.B2(n_424),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_493),
.A2(n_494),
.B1(n_499),
.B2(n_404),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_424),
.B1(n_434),
.B2(n_426),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_429),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_496),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_458),
.A2(n_434),
.B1(n_423),
.B2(n_440),
.Y(n_499)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_454),
.A2(n_440),
.B(n_421),
.C(n_442),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_500),
.A2(n_320),
.B(n_353),
.Y(n_533)
);

AOI21xp33_ASAP7_75t_L g502 ( 
.A1(n_461),
.A2(n_444),
.B(n_431),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_468),
.A2(n_459),
.B1(n_470),
.B2(n_475),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_451),
.B(n_415),
.Y(n_507)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_507),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_471),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_510),
.Y(n_534)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_480),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_448),
.B(n_421),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_468),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_513),
.B(n_515),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_456),
.B(n_442),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_447),
.C(n_452),
.Y(n_517)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_517),
.B(n_535),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_481),
.C(n_446),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_530),
.C(n_537),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_520),
.A2(n_523),
.B1(n_525),
.B2(n_545),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_492),
.A2(n_477),
.B(n_464),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_521),
.A2(n_529),
.B(n_543),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_522),
.A2(n_509),
.B1(n_490),
.B2(n_507),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_504),
.A2(n_418),
.B1(n_415),
.B2(n_432),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_488),
.A2(n_418),
.B1(n_432),
.B2(n_441),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_492),
.B(n_449),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_527),
.B(n_536),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_487),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_488),
.A2(n_443),
.B(n_425),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_425),
.C(n_320),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g569 ( 
.A(n_533),
.B(n_344),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_331),
.Y(n_535)
);

XOR2x1_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_404),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_353),
.C(n_301),
.Y(n_537)
);

CKINVDCx14_ASAP7_75t_R g538 ( 
.A(n_512),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_538),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_495),
.B(n_403),
.Y(n_540)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_540),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_541),
.A2(n_312),
.B1(n_344),
.B2(n_302),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_485),
.B(n_351),
.C(n_303),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_514),
.C(n_483),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_496),
.A2(n_346),
.B(n_302),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_496),
.A2(n_319),
.B1(n_346),
.B2(n_340),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_532),
.B(n_508),
.Y(n_546)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_546),
.Y(n_574)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_548),
.B(n_549),
.Y(n_582)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_544),
.Y(n_549)
);

A2O1A1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_527),
.A2(n_497),
.B(n_500),
.C(n_501),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_555),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_551),
.C(n_560),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_530),
.B(n_485),
.C(n_487),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g572 ( 
.A(n_556),
.B(n_524),
.Y(n_572)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_557),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_558),
.A2(n_562),
.B1(n_567),
.B2(n_545),
.Y(n_588)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_516),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_559),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_539),
.A2(n_493),
.B1(n_494),
.B2(n_500),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_561),
.A2(n_563),
.B1(n_565),
.B2(n_570),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_539),
.A2(n_500),
.B1(n_482),
.B2(n_498),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_520),
.A2(n_489),
.B1(n_491),
.B2(n_319),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_521),
.A2(n_340),
.B1(n_303),
.B2(n_312),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_531),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_568),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_533),
.Y(n_576)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_566),
.A2(n_526),
.B(n_517),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_571),
.B(n_575),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_572),
.B(n_581),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_518),
.Y(n_575)
);

XOR2x2_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_554),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_564),
.A2(n_529),
.B(n_519),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_577),
.B(n_579),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_524),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_535),
.C(n_542),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_585),
.B(n_586),
.C(n_587),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_536),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_541),
.Y(n_587)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_588),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_553),
.B(n_528),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_552),
.C(n_558),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_552),
.B(n_537),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_590),
.B(n_569),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_580),
.A2(n_564),
.B(n_550),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_592),
.A2(n_593),
.B(n_600),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_547),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_595),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_582),
.B(n_584),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_599),
.Y(n_614)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_573),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_576),
.A2(n_519),
.B(n_562),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_587),
.A2(n_554),
.B1(n_574),
.B2(n_561),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_601),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_573),
.B(n_546),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_605),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_604),
.B(n_589),
.Y(n_612)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_583),
.Y(n_605)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_583),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_607),
.B(n_559),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_603),
.A2(n_585),
.B(n_578),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_610),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_598),
.A2(n_569),
.B1(n_565),
.B2(n_586),
.Y(n_609)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_609),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_592),
.A2(n_567),
.B(n_543),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_611),
.B(n_612),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_606),
.B(n_581),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_SL g624 ( 
.A(n_613),
.B(n_606),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_598),
.A2(n_572),
.B1(n_306),
.B2(n_223),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_617),
.B(n_619),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_306),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_601),
.B(n_8),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_620),
.B(n_17),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_602),
.Y(n_622)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_622),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_624),
.B(n_625),
.Y(n_632)
);

OAI211xp5_ASAP7_75t_L g625 ( 
.A1(n_616),
.A2(n_618),
.B(n_600),
.C(n_617),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_615),
.B(n_591),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_629),
.B(n_630),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_621),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_631),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_623),
.B(n_616),
.C(n_621),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_633),
.B(n_16),
.C(n_634),
.Y(n_642)
);

AOI321xp33_ASAP7_75t_SL g636 ( 
.A1(n_628),
.A2(n_595),
.A3(n_609),
.B1(n_594),
.B2(n_591),
.C(n_610),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_636),
.A2(n_638),
.B1(n_16),
.B2(n_0),
.Y(n_641)
);

AO21x1_ASAP7_75t_SL g638 ( 
.A1(n_622),
.A2(n_13),
.B(n_15),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_637),
.Y(n_639)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_639),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_632),
.A2(n_626),
.B(n_627),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_640),
.A2(n_641),
.B(n_642),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_635),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_643),
.Y(n_646)
);

NAND2x1p5_ASAP7_75t_SL g647 ( 
.A(n_646),
.B(n_636),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_16),
.Y(n_648)
);


endmodule