module real_jpeg_20427_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_73;
wire n_65;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_31;
wire n_58;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_71;
wire n_47;
wire n_45;
wire n_25;
wire n_51;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_70;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_74;
wire n_16;
wire n_15;
wire n_13;

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_0),
.A2(n_16),
.B1(n_20),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_1),
.A2(n_16),
.B1(n_20),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_2),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_69)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_16),
.B1(n_20),
.B2(n_41),
.Y(n_45)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_8),
.B(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_15),
.B1(n_45),
.B2(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_33),
.B(n_37),
.C(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_16),
.B1(n_20),
.B2(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_55),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_42),
.B(n_54),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_26),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_13),
.B(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_15),
.A2(n_19),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_15),
.A2(n_24),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_28),
.B(n_34),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_32),
.A2(n_33),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_53),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_74),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_70),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);


endmodule