module fake_netlist_5_1573_n_1759 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1759);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1759;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g157 ( 
.A(n_5),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_0),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_80),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_124),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_8),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_91),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_43),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_82),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_84),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_33),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_42),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_109),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_34),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_83),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_29),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_78),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_72),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_68),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_66),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_100),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_32),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_20),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_131),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_127),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_102),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_22),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_95),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_21),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_81),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_23),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_19),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_29),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_34),
.Y(n_204)
);

BUFx8_ASAP7_75t_SL g205 ( 
.A(n_93),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_50),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_28),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_13),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_43),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_120),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_44),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_18),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_94),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_103),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_11),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_41),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_48),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_36),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_137),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_1),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_128),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_3),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_111),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_105),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_19),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_46),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_133),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_17),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_79),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_48),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_108),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_10),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_23),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_85),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_119),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_21),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_76),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_154),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_122),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_15),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_55),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_126),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_38),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_141),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_5),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_8),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_56),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_152),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_27),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_30),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_28),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_77),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_6),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_145),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_74),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_130),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_45),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_24),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_129),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_35),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_30),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_65),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_116),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_138),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_86),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_51),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_42),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_149),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_142),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_98),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_144),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_55),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_104),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_62),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_41),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_18),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_32),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_71),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_92),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_90),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_2),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_135),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_25),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_26),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_6),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_4),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_17),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_196),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_163),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_196),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_166),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_171),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_167),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_167),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_190),
.Y(n_323)
);

BUFx6f_ASAP7_75t_SL g324 ( 
.A(n_212),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_205),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_190),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_243),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_243),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_213),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_233),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_160),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_189),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_213),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_157),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_157),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_165),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_169),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_174),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_159),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_R g345 ( 
.A(n_179),
.B(n_57),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_182),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_159),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_162),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_183),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_162),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_165),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_184),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_175),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_173),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_173),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_201),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_161),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_188),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_210),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_192),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_271),
.B(n_2),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_193),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_202),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_220),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_202),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_218),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_216),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_223),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_223),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_240),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_177),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_236),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_170),
.B(n_4),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_254),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_236),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_177),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_194),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_239),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_275),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_291),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_216),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_195),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_259),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_200),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_208),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_261),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_316),
.B(n_214),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_313),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_319),
.B(n_259),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_314),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_321),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_315),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_221),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_318),
.B(n_225),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_227),
.Y(n_416)
);

BUFx8_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_353),
.B(n_212),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_329),
.A2(n_253),
.B1(n_257),
.B2(n_278),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_350),
.B(n_228),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_336),
.A2(n_197),
.B(n_186),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_323),
.B(n_161),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_326),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_330),
.A2(n_247),
.B(n_239),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_333),
.B(n_297),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_336),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_384),
.A2(n_181),
.B1(n_298),
.B2(n_222),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_338),
.A2(n_248),
.B(n_247),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_338),
.B(n_230),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_351),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_215),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_354),
.B(n_297),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

CKINVDCx11_ASAP7_75t_R g446 ( 
.A(n_334),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_356),
.B(n_235),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_321),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_356),
.B(n_186),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_376),
.B(n_306),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_392),
.B(n_332),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_339),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_397),
.B(n_341),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_398),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_342),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_403),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_418),
.A2(n_370),
.B1(n_203),
.B2(n_267),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_418),
.B(n_344),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_408),
.B(n_452),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_408),
.B(n_346),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_408),
.B(n_349),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_449),
.A2(n_203),
.B1(n_241),
.B2(n_276),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_446),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_403),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_446),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_SL g492 ( 
.A1(n_404),
.A2(n_425),
.B(n_444),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_439),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_452),
.B(n_352),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_439),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_355),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_404),
.B(n_359),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_452),
.B(n_361),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_412),
.B(n_363),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_441),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_390),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_452),
.B(n_197),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_441),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_448),
.B(n_380),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_441),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_448),
.B(n_387),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_448),
.B(n_321),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_436),
.A2(n_284),
.B1(n_211),
.B2(n_279),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_398),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_409),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_412),
.B(n_385),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_449),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_415),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_448),
.B(n_321),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_444),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_452),
.B(n_331),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_390),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_442),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_426),
.B(n_367),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_416),
.B(n_424),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_413),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_444),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_415),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_417),
.B(n_325),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_391),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_416),
.B(n_324),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_424),
.B(n_324),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_445),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_440),
.B(n_383),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_396),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_423),
.B(n_340),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_426),
.B(n_367),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_402),
.Y(n_548)
);

BUFx6f_ASAP7_75t_SL g549 ( 
.A(n_449),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_417),
.B(n_345),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_396),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_396),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_448),
.B(n_238),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_399),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_417),
.B(n_212),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_449),
.A2(n_276),
.B1(n_241),
.B2(n_267),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_402),
.B(n_158),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_449),
.A2(n_248),
.B1(n_263),
.B2(n_264),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_426),
.B(n_368),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_445),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_417),
.B(n_212),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_451),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_391),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_448),
.B(n_242),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_448),
.B(n_245),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_440),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_417),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_447),
.B(n_360),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_391),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_391),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_447),
.B(n_382),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_436),
.B(n_249),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_434),
.B(n_368),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_405),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_393),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_405),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_180),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_417),
.B(n_249),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_388),
.Y(n_586)
);

AND3x2_ASAP7_75t_L g587 ( 
.A(n_393),
.B(n_293),
.C(n_217),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_391),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_423),
.B(n_249),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_407),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_437),
.B(n_246),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_437),
.B(n_407),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_407),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_455),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_449),
.A2(n_229),
.B1(n_244),
.B2(n_237),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_391),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_391),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_437),
.B(n_250),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_388),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_437),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_434),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_437),
.B(n_366),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_456),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_456),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_492),
.A2(n_219),
.B(n_217),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_582),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_SL g609 ( 
.A(n_557),
.B(n_373),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_572),
.A2(n_377),
.B1(n_281),
.B2(n_274),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_533),
.B(n_435),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_435),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_526),
.B(n_435),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_466),
.B(n_164),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_480),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_527),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_582),
.B(n_434),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_526),
.B(n_435),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_474),
.B(n_172),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_535),
.B(n_435),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_535),
.B(n_435),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_457),
.B(n_461),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_484),
.B(n_435),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_573),
.B(n_249),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_499),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_605),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_573),
.B(n_429),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_605),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_506),
.B(n_435),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_548),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_520),
.B(n_191),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_506),
.B(n_435),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_606),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_492),
.A2(n_219),
.B(n_232),
.C(n_234),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_511),
.B(n_438),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_544),
.B(n_199),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_574),
.B(n_578),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_503),
.B(n_180),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_482),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_511),
.B(n_438),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_537),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_606),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_482),
.A2(n_299),
.B1(n_289),
.B2(n_282),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_513),
.B(n_438),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_490),
.A2(n_299),
.B(n_263),
.C(n_264),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_513),
.B(n_438),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_522),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g652 ( 
.A(n_529),
.B(n_224),
.C(n_209),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_528),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_503),
.B(n_180),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_522),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_531),
.B(n_539),
.Y(n_656)
);

BUFx8_ASAP7_75t_L g657 ( 
.A(n_532),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_603),
.B(n_204),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_528),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_532),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_531),
.B(n_438),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_490),
.A2(n_232),
.B(n_234),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_539),
.B(n_438),
.Y(n_663)
);

O2A1O1Ixp5_ASAP7_75t_L g664 ( 
.A1(n_493),
.A2(n_497),
.B(n_465),
.C(n_469),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_486),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_SL g666 ( 
.A1(n_590),
.A2(n_185),
.B1(n_304),
.B2(n_178),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_481),
.B(n_206),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_543),
.B(n_438),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_483),
.B(n_207),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_503),
.B(n_521),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_543),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_558),
.B(n_438),
.Y(n_672)
);

BUFx6f_ASAP7_75t_SL g673 ( 
.A(n_459),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_503),
.B(n_180),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_558),
.B(n_564),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_521),
.A2(n_285),
.B1(n_293),
.B2(n_258),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_495),
.B(n_226),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_468),
.B(n_415),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_564),
.B(n_438),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_567),
.B(n_429),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_547),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_482),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_567),
.B(n_429),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_489),
.A2(n_308),
.B1(n_282),
.B2(n_289),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_502),
.B(n_231),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_534),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_571),
.B(n_429),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_493),
.B(n_251),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_534),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_571),
.B(n_429),
.Y(n_690)
);

NAND2x1_ASAP7_75t_L g691 ( 
.A(n_497),
.B(n_464),
.Y(n_691)
);

NAND2x1_ASAP7_75t_L g692 ( 
.A(n_464),
.B(n_465),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_560),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_459),
.B(n_252),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_536),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_547),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_459),
.B(n_255),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_590),
.B(n_178),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_563),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_521),
.B(n_180),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_577),
.B(n_588),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_536),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_459),
.B(n_256),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_577),
.B(n_588),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_468),
.B(n_369),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_563),
.B(n_277),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_595),
.B(n_432),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_476),
.B(n_260),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_579),
.B(n_178),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_580),
.B(n_277),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_SL g711 ( 
.A(n_566),
.B(n_585),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_595),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_586),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_596),
.B(n_432),
.Y(n_714)
);

NOR2x1_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_509),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_489),
.B(n_391),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_586),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_601),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_489),
.B(n_391),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_469),
.A2(n_477),
.B1(n_473),
.B2(n_458),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_473),
.B(n_432),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_476),
.B(n_178),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_601),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_602),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_458),
.B(n_395),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_602),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_462),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_SL g730 ( 
.A1(n_509),
.A2(n_258),
.B1(n_292),
.B2(n_270),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_458),
.B(n_477),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_580),
.B(n_541),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_510),
.B(n_395),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_542),
.B(n_432),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_476),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_592),
.B(n_432),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_518),
.B(n_369),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_545),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_476),
.B(n_262),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_600),
.B(n_433),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_604),
.B(n_433),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_597),
.B(n_268),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_462),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_509),
.B(n_433),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_510),
.B(n_395),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_509),
.A2(n_265),
.B1(n_294),
.B2(n_287),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_597),
.B(n_272),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_509),
.B(n_433),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_510),
.A2(n_292),
.B(n_288),
.C(n_286),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_479),
.B(n_283),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_486),
.B(n_185),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_549),
.A2(n_296),
.B1(n_273),
.B2(n_285),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_562),
.A2(n_308),
.B1(n_266),
.B2(n_270),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_550),
.A2(n_288),
.B(n_286),
.C(n_280),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_518),
.B(n_371),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_549),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_517),
.B(n_290),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_433),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_559),
.B(n_371),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_467),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_587),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_545),
.B(n_450),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_467),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_552),
.B(n_553),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_523),
.B(n_372),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_550),
.A2(n_266),
.B1(n_280),
.B2(n_454),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_550),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_463),
.B(n_372),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_517),
.B(n_295),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_552),
.B(n_450),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_553),
.Y(n_771)
);

NAND2x1_ASAP7_75t_L g772 ( 
.A(n_599),
.B(n_388),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_488),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_485),
.B(n_277),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_523),
.Y(n_775)
);

OAI221xp5_ASAP7_75t_L g776 ( 
.A1(n_554),
.A2(n_427),
.B1(n_422),
.B2(n_414),
.C(n_430),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_554),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_556),
.B(n_450),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_726),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_623),
.B(n_556),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_664),
.A2(n_514),
.B(n_498),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_662),
.A2(n_512),
.B(n_460),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_633),
.A2(n_460),
.B(n_496),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_632),
.Y(n_784)
);

AND2x2_ASAP7_75t_SL g785 ( 
.A(n_640),
.B(n_584),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_633),
.A2(n_496),
.B(n_460),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_640),
.B(n_561),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_614),
.B(n_561),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_731),
.A2(n_594),
.B(n_591),
.C(n_583),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_614),
.B(n_565),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_728),
.Y(n_791)
);

AND2x4_ASAP7_75t_SL g792 ( 
.A(n_756),
.B(n_185),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_641),
.A2(n_581),
.B(n_594),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_641),
.A2(n_581),
.B(n_591),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_633),
.A2(n_589),
.B(n_460),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_633),
.A2(n_575),
.B(n_496),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_620),
.B(n_565),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_651),
.Y(n_798)
);

BUFx2_ASAP7_75t_R g799 ( 
.A(n_665),
.Y(n_799)
);

CKINVDCx10_ASAP7_75t_R g800 ( 
.A(n_673),
.Y(n_800)
);

INVx11_ASAP7_75t_L g801 ( 
.A(n_657),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_611),
.A2(n_589),
.B(n_496),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_612),
.A2(n_589),
.B(n_575),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_620),
.B(n_732),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_731),
.A2(n_583),
.B(n_538),
.C(n_471),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_717),
.B(n_634),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_696),
.B(n_546),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_634),
.A2(n_546),
.B(n_470),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_639),
.A2(n_569),
.B1(n_555),
.B2(n_570),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_639),
.B(n_463),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_654),
.A2(n_575),
.B(n_589),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_637),
.A2(n_501),
.B(n_471),
.C(n_472),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_628),
.B(n_463),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_630),
.B(n_463),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_742),
.A2(n_494),
.B(n_508),
.C(n_524),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_654),
.A2(n_575),
.B(n_598),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_636),
.B(n_494),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_618),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_674),
.A2(n_507),
.B(n_598),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_674),
.A2(n_507),
.B(n_598),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_742),
.A2(n_494),
.B(n_508),
.C(n_524),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_688),
.A2(n_507),
.B(n_598),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_655),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_716),
.A2(n_507),
.B(n_598),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_671),
.Y(n_825)
);

OAI21xp33_ASAP7_75t_L g826 ( 
.A1(n_757),
.A2(n_305),
.B(n_300),
.Y(n_826)
);

NAND2x1_ASAP7_75t_L g827 ( 
.A(n_682),
.B(n_599),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_757),
.B(n_307),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_712),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_716),
.A2(n_727),
.B(n_721),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_709),
.B(n_516),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_721),
.A2(n_525),
.B(n_487),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_727),
.A2(n_530),
.B(n_576),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_646),
.B(n_494),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_618),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_625),
.A2(n_530),
.B(n_576),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_733),
.A2(n_745),
.B(n_670),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_733),
.A2(n_530),
.B(n_576),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_745),
.A2(n_530),
.B(n_576),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_670),
.A2(n_530),
.B(n_576),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_618),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_657),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_736),
.A2(n_507),
.B(n_568),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_738),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_608),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_682),
.B(n_540),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_769),
.A2(n_310),
.B(n_311),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_747),
.A2(n_508),
.B(n_524),
.C(n_475),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_649),
.A2(n_504),
.B(n_519),
.C(n_515),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_682),
.B(n_540),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_669),
.A2(n_524),
.B1(n_508),
.B2(n_599),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_669),
.B(n_766),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_766),
.B(n_642),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_769),
.B(n_309),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_642),
.B(n_472),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_660),
.B(n_475),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_627),
.B(n_478),
.Y(n_857)
);

AOI21xp33_ASAP7_75t_L g858 ( 
.A1(n_747),
.A2(n_488),
.B(n_422),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_667),
.A2(n_677),
.B(n_685),
.C(n_750),
.Y(n_859)
);

AO21x1_ASAP7_75t_L g860 ( 
.A1(n_607),
.A2(n_711),
.B(n_676),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_627),
.B(n_478),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_681),
.B(n_487),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_775),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_691),
.A2(n_504),
.B(n_500),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_692),
.A2(n_500),
.B(n_501),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_667),
.B(n_515),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_740),
.A2(n_568),
.B(n_540),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_624),
.B(n_519),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_682),
.B(n_540),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_741),
.B(n_540),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_699),
.B(n_568),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_773),
.B(n_185),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_756),
.B(n_759),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_723),
.A2(n_568),
.B(n_491),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_647),
.B(n_568),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_647),
.B(n_450),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_698),
.B(n_599),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_771),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_777),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_656),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_684),
.B(n_453),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_758),
.A2(n_491),
.B(n_406),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_613),
.A2(n_491),
.B(n_406),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_705),
.B(n_9),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_684),
.B(n_453),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_737),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_749),
.A2(n_454),
.B(n_453),
.C(n_414),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_713),
.Y(n_888)
);

AND2x6_ASAP7_75t_L g889 ( 
.A(n_715),
.B(n_375),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_675),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_759),
.B(n_375),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_724),
.B(n_378),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_701),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_619),
.A2(n_491),
.B(n_406),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_645),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_706),
.B(n_453),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_704),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_621),
.A2(n_491),
.B(n_395),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_754),
.A2(n_454),
.B(n_430),
.C(n_427),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_710),
.B(n_454),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_767),
.B(n_419),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_730),
.A2(n_414),
.B(n_427),
.C(n_422),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_622),
.A2(n_491),
.B(n_406),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_767),
.A2(n_722),
.B1(n_693),
.B2(n_744),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_629),
.B(n_406),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_658),
.B(n_428),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_645),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_755),
.Y(n_908)
);

NOR2x1_ASAP7_75t_R g909 ( 
.A(n_735),
.B(n_378),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_658),
.B(n_428),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_677),
.A2(n_430),
.B1(n_428),
.B2(n_421),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_729),
.Y(n_912)
);

NOR2x2_ASAP7_75t_L g913 ( 
.A(n_666),
.B(n_626),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_765),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_694),
.B(n_428),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_694),
.B(n_421),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_743),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_760),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_761),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_644),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_697),
.B(n_421),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_748),
.A2(n_388),
.B(n_389),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_SL g923 ( 
.A1(n_700),
.A2(n_381),
.B(n_389),
.C(n_419),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_697),
.B(n_10),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_774),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_768),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_652),
.B(n_381),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_703),
.B(n_406),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_673),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_703),
.B(n_421),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_708),
.B(n_419),
.Y(n_931)
);

NOR2xp67_ASAP7_75t_L g932 ( 
.A(n_610),
.B(n_87),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_763),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_708),
.B(n_11),
.Y(n_934)
);

AOI21x1_ASAP7_75t_L g935 ( 
.A1(n_734),
.A2(n_389),
.B(n_419),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_700),
.A2(n_401),
.B(n_395),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_764),
.A2(n_401),
.B(n_395),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_739),
.B(n_15),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_739),
.B(n_401),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_645),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_750),
.A2(n_411),
.B(n_389),
.C(n_304),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_685),
.A2(n_411),
.B(n_420),
.C(n_401),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_761),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_722),
.A2(n_406),
.B1(n_401),
.B2(n_400),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_678),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_680),
.B(n_406),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_751),
.B(n_304),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_746),
.A2(n_411),
.B(n_420),
.C(n_401),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_616),
.B(n_304),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_609),
.B(n_406),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_683),
.A2(n_401),
.B(n_400),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_722),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_687),
.A2(n_401),
.B(n_400),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_SL g954 ( 
.A1(n_753),
.A2(n_411),
.B(n_20),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_768),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_690),
.A2(n_401),
.B(n_400),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_707),
.B(n_400),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_772),
.A2(n_778),
.B(n_762),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_753),
.B(n_411),
.Y(n_959)
);

BUFx4f_ASAP7_75t_L g960 ( 
.A(n_768),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_714),
.A2(n_776),
.B(n_672),
.C(n_668),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_631),
.A2(n_400),
.B(n_395),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_615),
.B(n_400),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_617),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_752),
.B(n_400),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_635),
.A2(n_400),
.B(n_395),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_638),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_653),
.B(n_395),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_798),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_859),
.B(n_650),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_870),
.A2(n_782),
.B(n_780),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_852),
.A2(n_661),
.B1(n_643),
.B2(n_663),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_873),
.B(n_768),
.Y(n_973)
);

HAxp5_ASAP7_75t_L g974 ( 
.A(n_808),
.B(n_16),
.CON(n_974),
.SN(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_920),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_804),
.B(n_806),
.Y(n_976)
);

AO22x1_ASAP7_75t_L g977 ( 
.A1(n_828),
.A2(n_768),
.B1(n_648),
.B2(n_679),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_806),
.B(n_702),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_895),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_828),
.A2(n_695),
.B1(n_725),
.B2(n_720),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_895),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_SL g982 ( 
.A1(n_854),
.A2(n_16),
.B1(n_24),
.B2(n_25),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_783),
.A2(n_770),
.B(n_719),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_786),
.A2(n_718),
.B(n_689),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_825),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_863),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_955),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_779),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_795),
.A2(n_686),
.B(n_659),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_914),
.B(n_886),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_854),
.A2(n_420),
.B(n_31),
.C(n_37),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_914),
.B(n_420),
.Y(n_992)
);

NAND2x1p5_ASAP7_75t_L g993 ( 
.A(n_895),
.B(n_420),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_880),
.B(n_420),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_895),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_890),
.B(n_420),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_893),
.B(n_420),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_945),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_823),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_796),
.A2(n_410),
.B(n_420),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_853),
.A2(n_410),
.B(n_73),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_897),
.B(n_410),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_791),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_908),
.B(n_26),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_810),
.A2(n_410),
.B(n_75),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_924),
.A2(n_70),
.B(n_150),
.C(n_147),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_924),
.A2(n_31),
.B(n_37),
.C(n_38),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_829),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_934),
.A2(n_410),
.B1(n_88),
.B2(n_89),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_928),
.A2(n_410),
.B(n_64),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_788),
.B(n_410),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_945),
.B(n_39),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_803),
.A2(n_410),
.B(n_106),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_842),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_SL g1015 ( 
.A1(n_934),
.A2(n_60),
.B(n_146),
.C(n_143),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_784),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_836),
.A2(n_867),
.B(n_843),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_L g1018 ( 
.A(n_940),
.B(n_410),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_888),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_787),
.B(n_39),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_955),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_856),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_818),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_844),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_785),
.A2(n_59),
.B1(n_134),
.B2(n_125),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_925),
.B(n_40),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_952),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_891),
.B(n_868),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_879),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_938),
.A2(n_40),
.B1(n_47),
.B2(n_49),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_790),
.B(n_58),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_785),
.A2(n_107),
.B1(n_121),
.B2(n_117),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_807),
.B(n_49),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_797),
.B(n_139),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_830),
.A2(n_837),
.B(n_821),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_925),
.B(n_50),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_SL g1037 ( 
.A1(n_950),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_891),
.B(n_52),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_938),
.A2(n_53),
.B(n_54),
.C(n_56),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_860),
.A2(n_54),
.B1(n_112),
.B2(n_113),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_868),
.B(n_114),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_967),
.B(n_857),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_907),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_892),
.B(n_904),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_822),
.A2(n_802),
.B(n_811),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_815),
.A2(n_875),
.B(n_848),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_967),
.B(n_857),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_862),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_892),
.B(n_896),
.Y(n_1049)
);

AO22x1_ASAP7_75t_L g1050 ( 
.A1(n_949),
.A2(n_947),
.B1(n_884),
.B2(n_873),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_907),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_939),
.A2(n_900),
.B(n_866),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_878),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_912),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_861),
.B(n_906),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_SL g1056 ( 
.A1(n_858),
.A2(n_831),
.B(n_965),
.C(n_916),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_917),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_855),
.A2(n_816),
.B(n_869),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_918),
.Y(n_1059)
);

OAI22x1_ASAP7_75t_L g1060 ( 
.A1(n_884),
.A2(n_841),
.B1(n_818),
.B2(n_835),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_915),
.A2(n_921),
.B(n_931),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_943),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_861),
.B(n_910),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_846),
.A2(n_850),
.B(n_930),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_877),
.A2(n_871),
.B1(n_960),
.B2(n_881),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_933),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_927),
.B(n_959),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_840),
.A2(n_819),
.B(n_820),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_927),
.B(n_877),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_960),
.B(n_932),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_SL g1071 ( 
.A(n_872),
.B(n_847),
.C(n_826),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_901),
.B(n_889),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_889),
.B(n_964),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_805),
.A2(n_941),
.B(n_954),
.C(n_961),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_835),
.A2(n_841),
.B(n_943),
.C(n_902),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_907),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_SL g1077 ( 
.A1(n_948),
.A2(n_942),
.B(n_834),
.C(n_813),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_919),
.A2(n_923),
.B(n_817),
.C(n_814),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_889),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_955),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_799),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_845),
.B(n_909),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_889),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_958),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_824),
.A2(n_833),
.B(n_839),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_876),
.A2(n_885),
.B(n_789),
.C(n_812),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_SL g1087 ( 
.A(n_940),
.B(n_955),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_889),
.B(n_911),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_792),
.B(n_929),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_926),
.B(n_851),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_827),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_838),
.A2(n_781),
.B(n_874),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_809),
.A2(n_832),
.B(n_793),
.C(n_794),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_963),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_946),
.A2(n_957),
.B(n_922),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_801),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_849),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_800),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_926),
.B(n_944),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_899),
.A2(n_887),
.B(n_968),
.C(n_864),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_SL g1101 ( 
.A1(n_865),
.A2(n_882),
.B(n_936),
.C(n_951),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_913),
.A2(n_905),
.B(n_937),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_883),
.B(n_894),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_935),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_905),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_953),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_962),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_966),
.B(n_956),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_898),
.B(n_903),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_955),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_870),
.A2(n_633),
.B(n_670),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_914),
.B(n_886),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_870),
.A2(n_633),
.B(n_670),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_914),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_859),
.A2(n_640),
.B(n_854),
.C(n_828),
.Y(n_1115)
);

CKINVDCx8_ASAP7_75t_R g1116 ( 
.A(n_800),
.Y(n_1116)
);

OR2x6_ASAP7_75t_SL g1117 ( 
.A(n_929),
.B(n_486),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_976),
.B(n_1115),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1016),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_971),
.A2(n_1052),
.B(n_1045),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_SL g1121 ( 
.A1(n_1067),
.A2(n_1075),
.B(n_1069),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_976),
.A2(n_1044),
.B(n_974),
.C(n_991),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1028),
.B(n_1022),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_1030),
.A2(n_1036),
.B(n_1026),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1048),
.B(n_1042),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_979),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1095),
.A2(n_1092),
.B(n_1035),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_L g1129 ( 
.A(n_1050),
.B(n_1071),
.C(n_1039),
.Y(n_1129)
);

O2A1O1Ixp5_ASAP7_75t_L g1130 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_1034),
.C(n_970),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1047),
.B(n_1055),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1063),
.B(n_978),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1033),
.A2(n_1102),
.B1(n_975),
.B2(n_1082),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1030),
.A2(n_982),
.B(n_1040),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1109),
.A2(n_1093),
.B(n_970),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1074),
.A2(n_1084),
.A3(n_1104),
.B(n_1086),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1068),
.A2(n_1085),
.B(n_1058),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1093),
.A2(n_1101),
.B(n_1103),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1046),
.A2(n_1056),
.B(n_1086),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1089),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_1077),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1099),
.A2(n_972),
.B(n_1011),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1000),
.A2(n_983),
.B(n_984),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_974),
.B(n_990),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_989),
.A2(n_1010),
.B(n_1107),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_973),
.B(n_981),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_991),
.A2(n_1007),
.B(n_1036),
.C(n_1026),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_985),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1082),
.A2(n_986),
.B1(n_998),
.B2(n_1089),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1077),
.A2(n_1108),
.B(n_1064),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1041),
.A2(n_978),
.B(n_1099),
.C(n_1040),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_SL g1152 ( 
.A(n_1096),
.B(n_1081),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1013),
.A2(n_1100),
.B(n_1090),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1065),
.A2(n_1090),
.B(n_1011),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_982),
.A2(n_1020),
.B1(n_1009),
.B2(n_1049),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1106),
.A2(n_977),
.B(n_1070),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1112),
.B(n_1114),
.Y(n_1157)
);

INVx5_ASAP7_75t_L g1158 ( 
.A(n_979),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1054),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1038),
.A2(n_1012),
.B1(n_1114),
.B2(n_1062),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1001),
.A2(n_1060),
.A3(n_1005),
.B(n_1088),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1097),
.A2(n_1072),
.A3(n_980),
.B(n_1073),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1106),
.A2(n_1070),
.B(n_1049),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1059),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_999),
.A2(n_1008),
.B1(n_988),
.B2(n_1003),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1031),
.A2(n_1034),
.B(n_1061),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1106),
.A2(n_997),
.B(n_994),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1066),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_992),
.B(n_1029),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1024),
.B(n_1057),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1106),
.A2(n_994),
.B(n_997),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1094),
.A2(n_996),
.A3(n_1002),
.B(n_1025),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1019),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1078),
.A2(n_993),
.B(n_1018),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_1096),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1027),
.B(n_1023),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1079),
.A2(n_1083),
.B(n_1006),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1079),
.A2(n_1083),
.B(n_1006),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_993),
.A2(n_1021),
.B(n_987),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1032),
.A2(n_1015),
.B(n_973),
.C(n_1023),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_SL g1181 ( 
.A(n_1105),
.B(n_979),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1027),
.B(n_1004),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1043),
.B(n_1076),
.Y(n_1183)
);

AOI221x1_ASAP7_75t_L g1184 ( 
.A1(n_1037),
.A2(n_1015),
.B1(n_987),
.B2(n_1110),
.C(n_1021),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_979),
.Y(n_1185)
);

AO32x2_ASAP7_75t_L g1186 ( 
.A1(n_995),
.A2(n_1051),
.A3(n_1076),
.B1(n_1087),
.B2(n_1080),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1110),
.B(n_995),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1091),
.A2(n_1080),
.B(n_1051),
.C(n_1117),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1080),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1014),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1116),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1091),
.A2(n_1080),
.B(n_1098),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1091),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1091),
.A2(n_1115),
.B(n_859),
.C(n_640),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1115),
.A2(n_860),
.A3(n_1074),
.B(n_859),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1115),
.A2(n_859),
.B(n_852),
.C(n_991),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1080),
.Y(n_1197)
);

INVxp67_ASAP7_75t_SL g1198 ( 
.A(n_1114),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1115),
.A2(n_859),
.B1(n_852),
.B2(n_647),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1115),
.A2(n_860),
.A3(n_1074),
.B(n_859),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_977),
.A2(n_970),
.B(n_1011),
.Y(n_1201)
);

AOI221xp5_ASAP7_75t_L g1202 ( 
.A1(n_1115),
.A2(n_854),
.B1(n_828),
.B2(n_640),
.C(n_769),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_969),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_979),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_969),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1115),
.B(n_806),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_976),
.B(n_640),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1115),
.A2(n_859),
.B1(n_640),
.B2(n_854),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1211)
);

BUFx4f_ASAP7_75t_SL g1212 ( 
.A(n_975),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_976),
.B(n_640),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_976),
.B(n_640),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_976),
.B(n_640),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_976),
.B(n_640),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1219)
);

OAI22x1_ASAP7_75t_L g1220 ( 
.A1(n_976),
.A2(n_854),
.B1(n_828),
.B2(n_934),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1115),
.A2(n_859),
.B1(n_640),
.B2(n_854),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1115),
.A2(n_859),
.B(n_682),
.Y(n_1222)
);

NAND3xp33_ASAP7_75t_L g1223 ( 
.A(n_1115),
.B(n_640),
.C(n_859),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1115),
.B(n_806),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1053),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1115),
.A2(n_859),
.B(n_640),
.C(n_854),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_974),
.B(n_807),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1115),
.A2(n_859),
.B1(n_852),
.B2(n_647),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1115),
.A2(n_859),
.B(n_852),
.C(n_991),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_976),
.B(n_640),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1050),
.B(n_895),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_969),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1096),
.B(n_945),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_976),
.B(n_640),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1087),
.B(n_995),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_969),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_1089),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_976),
.B(n_640),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1071),
.A2(n_854),
.B1(n_828),
.B2(n_640),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_974),
.B(n_807),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_SL g1250 ( 
.A1(n_1067),
.A2(n_860),
.B(n_1075),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1115),
.A2(n_859),
.B(n_640),
.C(n_854),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1115),
.A2(n_860),
.A3(n_1074),
.B(n_859),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_976),
.B(n_640),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1016),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1050),
.B(n_895),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1017),
.A2(n_1113),
.B(n_1111),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1115),
.A2(n_859),
.B1(n_1030),
.B2(n_934),
.C(n_938),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1262)
);

AOI21xp33_ASAP7_75t_L g1263 ( 
.A1(n_1115),
.A2(n_640),
.B(n_828),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1115),
.A2(n_859),
.B(n_1046),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_971),
.A2(n_633),
.B(n_1052),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1202),
.A2(n_1125),
.B1(n_1248),
.B2(n_1263),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1209),
.B(n_1132),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1191),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1148),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1255),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1158),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1119),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1212),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1151),
.A2(n_1228),
.B1(n_1133),
.B2(n_1210),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1221),
.A2(n_1223),
.B1(n_1245),
.B2(n_1257),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1175),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1131),
.B(n_1213),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1215),
.B(n_1216),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1223),
.A2(n_1245),
.B1(n_1259),
.B2(n_1244),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1226),
.A2(n_1247),
.B1(n_1257),
.B2(n_1259),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1134),
.A2(n_1126),
.B1(n_1149),
.B2(n_1251),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1140),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1226),
.A2(n_1264),
.B1(n_1244),
.B2(n_1247),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1203),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1264),
.A2(n_1129),
.B1(n_1206),
.B2(n_1224),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1190),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1155),
.A2(n_1249),
.B1(n_1229),
.B2(n_1230),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1134),
.A2(n_1194),
.B1(n_1124),
.B2(n_1218),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1198),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1205),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1176),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1183),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1183),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1242),
.Y(n_1294)
);

INVx5_ASAP7_75t_L g1295 ( 
.A(n_1127),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1199),
.A2(n_1230),
.B1(n_1155),
.B2(n_1118),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1232),
.A2(n_1239),
.B1(n_1246),
.B2(n_1253),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1199),
.A2(n_1144),
.B1(n_1152),
.B2(n_1121),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1235),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1241),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1159),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1204),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1220),
.A2(n_1139),
.B1(n_1142),
.B2(n_1160),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1146),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1182),
.A2(n_1234),
.B1(n_1258),
.B2(n_1147),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1152),
.A2(n_1139),
.B1(n_1258),
.B2(n_1234),
.Y(n_1307)
);

CKINVDCx9p33_ASAP7_75t_R g1308 ( 
.A(n_1187),
.Y(n_1308)
);

CKINVDCx6p67_ASAP7_75t_R g1309 ( 
.A(n_1204),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1234),
.A2(n_1258),
.B1(n_1250),
.B2(n_1261),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1168),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1240),
.A2(n_1146),
.B1(n_1227),
.B2(n_1170),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1261),
.A2(n_1142),
.B1(n_1181),
.B2(n_1166),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1173),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1122),
.B(n_1157),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1169),
.A2(n_1165),
.B1(n_1192),
.B2(n_1163),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1180),
.A2(n_1178),
.B(n_1177),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1154),
.A2(n_1128),
.B1(n_1135),
.B2(n_1166),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1193),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1240),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1197),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1195),
.B(n_1252),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1186),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1153),
.A2(n_1156),
.B1(n_1196),
.B2(n_1231),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1186),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1141),
.A2(n_1138),
.B1(n_1150),
.B2(n_1171),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1222),
.A2(n_1252),
.B1(n_1200),
.B2(n_1195),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1197),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1186),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1185),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1167),
.A2(n_1238),
.B1(n_1120),
.B2(n_1265),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1207),
.A2(n_1262),
.B1(n_1208),
.B2(n_1214),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1185),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1195),
.A2(n_1200),
.B1(n_1252),
.B2(n_1174),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1200),
.A2(n_1130),
.B1(n_1243),
.B2(n_1237),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1162),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1189),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1217),
.A2(n_1219),
.B1(n_1179),
.B2(n_1260),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1188),
.A2(n_1201),
.B1(n_1172),
.B2(n_1184),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1145),
.A2(n_1123),
.B1(n_1256),
.B2(n_1254),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1137),
.A2(n_1143),
.B(n_1236),
.Y(n_1341)
);

INVx6_ASAP7_75t_L g1342 ( 
.A(n_1161),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1172),
.A2(n_1161),
.B1(n_1211),
.B2(n_1225),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1172),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1233),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1202),
.A2(n_640),
.B(n_1115),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1202),
.A2(n_1125),
.B1(n_828),
.B2(n_854),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_1183),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1210),
.A2(n_828),
.B1(n_854),
.B2(n_640),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1119),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1119),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1119),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1119),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1210),
.A2(n_828),
.B1(n_854),
.B2(n_640),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1127),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1255),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1209),
.B(n_640),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1136),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1134),
.A2(n_709),
.B1(n_698),
.B2(n_1202),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1202),
.A2(n_1248),
.B1(n_1115),
.B2(n_854),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1136),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1158),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1136),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1136),
.Y(n_1364)
);

OAI21xp33_ASAP7_75t_L g1365 ( 
.A1(n_1202),
.A2(n_854),
.B(n_828),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1119),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1134),
.A2(n_709),
.B1(n_698),
.B2(n_1202),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1202),
.A2(n_1248),
.B1(n_1115),
.B2(n_854),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1119),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1191),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1212),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1210),
.A2(n_828),
.B1(n_854),
.B2(n_640),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1148),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1158),
.Y(n_1374)
);

BUFx8_ASAP7_75t_L g1375 ( 
.A(n_1191),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1158),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1191),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1119),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1209),
.B(n_640),
.Y(n_1379)
);

INVx8_ASAP7_75t_L g1380 ( 
.A(n_1158),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1202),
.A2(n_1125),
.B1(n_828),
.B2(n_854),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1202),
.A2(n_1248),
.B1(n_1115),
.B2(n_854),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1341),
.A2(n_1346),
.B(n_1343),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1284),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1340),
.A2(n_1332),
.B(n_1326),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1336),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1350),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1284),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1311),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1311),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1289),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1289),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1358),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1287),
.B(n_1296),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1291),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1333),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1322),
.B(n_1361),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1340),
.A2(n_1332),
.B(n_1326),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1318),
.A2(n_1317),
.B(n_1303),
.Y(n_1400)
);

INVx5_ASAP7_75t_SL g1401 ( 
.A(n_1308),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1268),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1329),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1290),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1296),
.B(n_1279),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1331),
.A2(n_1318),
.B(n_1345),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1299),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1331),
.A2(n_1339),
.B(n_1275),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1300),
.B(n_1301),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1370),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1316),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1359),
.A2(n_1367),
.B(n_1365),
.C(n_1382),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1303),
.A2(n_1275),
.B(n_1279),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1342),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1360),
.A2(n_1368),
.B(n_1274),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1306),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1308),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1281),
.B(n_1280),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1349),
.A2(n_1354),
.B(n_1372),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1285),
.B(n_1280),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1357),
.B(n_1379),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1269),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1377),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1267),
.B(n_1278),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1334),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1320),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1327),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1271),
.B(n_1295),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1356),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1283),
.A2(n_1285),
.B(n_1266),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1283),
.A2(n_1288),
.B(n_1305),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1347),
.A2(n_1381),
.B1(n_1266),
.B2(n_1359),
.Y(n_1433)
);

AO21x1_ASAP7_75t_L g1434 ( 
.A1(n_1367),
.A2(n_1316),
.B(n_1315),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1347),
.A2(n_1381),
.B(n_1297),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1271),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1351),
.B(n_1353),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1312),
.Y(n_1438)
);

INVxp33_ASAP7_75t_L g1439 ( 
.A(n_1304),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1277),
.B(n_1298),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1373),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1330),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_SL g1443 ( 
.A(n_1273),
.B(n_1371),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1319),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1344),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1313),
.B(n_1310),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1328),
.A2(n_1314),
.B(n_1321),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1324),
.Y(n_1448)
);

INVxp33_ASAP7_75t_L g1449 ( 
.A(n_1272),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1337),
.Y(n_1450)
);

NOR2x1p5_ASAP7_75t_L g1451 ( 
.A(n_1282),
.B(n_1294),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1335),
.A2(n_1307),
.B(n_1338),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1272),
.B(n_1369),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1380),
.A2(n_1362),
.B(n_1309),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1276),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1380),
.B(n_1376),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1405),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1420),
.A2(n_1352),
.B(n_1369),
.C(n_1366),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1426),
.B(n_1355),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1452),
.A2(n_1352),
.B(n_1378),
.C(n_1380),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1384),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1425),
.B(n_1292),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1426),
.B(n_1355),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1410),
.B(n_1428),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1432),
.A2(n_1433),
.B(n_1435),
.C(n_1394),
.Y(n_1465)
);

A2O1A1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1432),
.A2(n_1376),
.B(n_1374),
.C(n_1302),
.Y(n_1466)
);

NAND2x1_ASAP7_75t_L g1467 ( 
.A(n_1391),
.B(n_1376),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1384),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1409),
.B(n_1374),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_SL g1470 ( 
.A1(n_1440),
.A2(n_1286),
.B(n_1375),
.C(n_1374),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1427),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1428),
.B(n_1292),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_SL g1473 ( 
.A(n_1454),
.B(n_1270),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1409),
.A2(n_1385),
.B(n_1398),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1395),
.B(n_1293),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1435),
.A2(n_1348),
.B(n_1375),
.C(n_1394),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1397),
.B(n_1408),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1413),
.B(n_1419),
.C(n_1431),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1447),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1415),
.B(n_1397),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1417),
.B(n_1400),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_L g1482 ( 
.A(n_1419),
.B(n_1406),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1416),
.A2(n_1412),
.B(n_1421),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1404),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1417),
.B(n_1400),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1404),
.B(n_1402),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1400),
.B(n_1399),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1422),
.B(n_1396),
.Y(n_1488)
);

OAI211xp5_ASAP7_75t_L g1489 ( 
.A1(n_1416),
.A2(n_1431),
.B(n_1400),
.C(n_1438),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1437),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1434),
.A2(n_1421),
.B1(n_1446),
.B2(n_1448),
.C(n_1406),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_SL g1492 ( 
.A(n_1403),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1392),
.B(n_1386),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1399),
.B(n_1388),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1392),
.B(n_1386),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1438),
.A2(n_1446),
.B1(n_1431),
.B2(n_1421),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1385),
.A2(n_1398),
.B(n_1407),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1423),
.B(n_1444),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1383),
.A2(n_1434),
.B(n_1407),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1388),
.B(n_1389),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1389),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1445),
.A2(n_1424),
.B1(n_1439),
.B2(n_1418),
.Y(n_1502)
);

NAND2xp33_ASAP7_75t_L g1503 ( 
.A(n_1436),
.B(n_1429),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1390),
.B(n_1445),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1390),
.B(n_1441),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1486),
.B(n_1383),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1484),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1383),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1481),
.B(n_1414),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1461),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1496),
.A2(n_1491),
.B(n_1478),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1486),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1481),
.B(n_1414),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1482),
.A2(n_1421),
.B1(n_1431),
.B2(n_1414),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1485),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1465),
.A2(n_1414),
.B1(n_1401),
.B2(n_1448),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1393),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1477),
.B(n_1485),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1494),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1488),
.B(n_1449),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1457),
.B(n_1498),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1482),
.A2(n_1401),
.B1(n_1442),
.B2(n_1403),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1468),
.Y(n_1523)
);

AOI222xp33_ASAP7_75t_L g1524 ( 
.A1(n_1483),
.A2(n_1401),
.B1(n_1430),
.B2(n_1387),
.C1(n_1442),
.C2(n_1411),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1501),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1500),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1493),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_SL g1529 ( 
.A(n_1471),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1490),
.B(n_1453),
.Y(n_1530)
);

OAI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1462),
.A2(n_1453),
.B1(n_1450),
.B2(n_1411),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1505),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1495),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1510),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1523),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1516),
.A2(n_1458),
.B(n_1460),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1528),
.B(n_1533),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1519),
.B(n_1497),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1510),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1523),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1526),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1522),
.A2(n_1492),
.B1(n_1455),
.B2(n_1502),
.Y(n_1542)
);

AOI211xp5_ASAP7_75t_L g1543 ( 
.A1(n_1511),
.A2(n_1489),
.B(n_1476),
.C(n_1470),
.Y(n_1543)
);

OAI211xp5_ASAP7_75t_L g1544 ( 
.A1(n_1511),
.A2(n_1466),
.B(n_1475),
.C(n_1497),
.Y(n_1544)
);

INVxp33_ASAP7_75t_L g1545 ( 
.A(n_1520),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1508),
.B(n_1499),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1508),
.B(n_1499),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_1495),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1516),
.A2(n_1473),
.B(n_1469),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1508),
.B(n_1464),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1515),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1514),
.A2(n_1401),
.B1(n_1464),
.B2(n_1469),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.B(n_1513),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1514),
.A2(n_1503),
.B1(n_1469),
.B2(n_1472),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1531),
.A2(n_1469),
.B1(n_1471),
.B2(n_1450),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1531),
.A2(n_1436),
.B1(n_1467),
.B2(n_1456),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1559)
);

OAI211xp5_ASAP7_75t_L g1560 ( 
.A1(n_1524),
.A2(n_1504),
.B(n_1463),
.C(n_1459),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1504),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1507),
.Y(n_1563)
);

NAND2x1_ASAP7_75t_SL g1564 ( 
.A(n_1546),
.B(n_1525),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1553),
.B(n_1533),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1557),
.B(n_1558),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1534),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1545),
.B(n_1521),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1553),
.B(n_1506),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1538),
.B(n_1546),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1535),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1540),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1562),
.B(n_1512),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1562),
.B(n_1548),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1540),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1530),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1563),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_R g1582 ( 
.A(n_1536),
.B(n_1455),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1532),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1518),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1518),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1557),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1570),
.B(n_1557),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1569),
.B(n_1548),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1573),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1573),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1570),
.B(n_1557),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1570),
.B(n_1558),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1567),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1573),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1566),
.B(n_1558),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1582),
.B(n_1543),
.C(n_1544),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1574),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1566),
.B(n_1558),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1577),
.B(n_1550),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1577),
.B(n_1550),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1574),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1567),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1574),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1537),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1564),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1564),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1567),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1575),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1578),
.B(n_1537),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1571),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1579),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1579),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1582),
.A2(n_1543),
.B(n_1549),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1579),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1566),
.B(n_1539),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1568),
.B(n_1542),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1568),
.B(n_1541),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1586),
.B(n_1561),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1569),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1588),
.B(n_1572),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1605),
.B(n_1572),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1605),
.B(n_1565),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1623),
.B(n_1576),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1624),
.B(n_1565),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1617),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1623),
.B(n_1576),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1617),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1594),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1608),
.B(n_1566),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1624),
.B(n_1584),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1601),
.B(n_1566),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1601),
.B(n_1566),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1601),
.B(n_1586),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1594),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1620),
.B(n_1586),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1620),
.B(n_1554),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1590),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1607),
.B(n_1584),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1597),
.B(n_1554),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_SL g1650 ( 
.A(n_1597),
.B(n_1542),
.Y(n_1650)
);

NAND4xp25_ASAP7_75t_SL g1651 ( 
.A(n_1607),
.B(n_1524),
.C(n_1560),
.D(n_1569),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1584),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1594),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1590),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1583),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1589),
.B(n_1443),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1591),
.B(n_1585),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1591),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1589),
.B(n_1583),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1594),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1647),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1638),
.B(n_1609),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1630),
.B(n_1612),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_SL g1664 ( 
.A(n_1650),
.B(n_1609),
.C(n_1560),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1650),
.B(n_1589),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1656),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1641),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1641),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1649),
.A2(n_1609),
.B(n_1608),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1632),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1647),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1638),
.B(n_1596),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1646),
.A2(n_1651),
.B(n_1633),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1627),
.A2(n_1608),
.B(n_1555),
.C(n_1556),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1632),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_L g1676 ( 
.A(n_1627),
.B(n_1556),
.C(n_1552),
.Y(n_1676)
);

AOI222xp33_ASAP7_75t_L g1677 ( 
.A1(n_1628),
.A2(n_1552),
.B1(n_1555),
.B2(n_1612),
.C1(n_1616),
.C2(n_1625),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1645),
.A2(n_1596),
.B1(n_1599),
.B2(n_1622),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1628),
.A2(n_1564),
.B1(n_1598),
.B2(n_1621),
.C(n_1595),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1645),
.A2(n_1606),
.B(n_1604),
.C(n_1611),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1629),
.A2(n_1529),
.B1(n_1596),
.B2(n_1599),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1631),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1634),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1639),
.B(n_1612),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1673),
.B(n_1631),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1665),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1661),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1664),
.A2(n_1634),
.B1(n_1639),
.B2(n_1640),
.C(n_1626),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1669),
.A2(n_1626),
.B(n_1640),
.C(n_1636),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1671),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1670),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1670),
.B(n_1654),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1675),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1683),
.B(n_1655),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1662),
.B(n_1655),
.Y(n_1696)
);

AOI222xp33_ASAP7_75t_L g1697 ( 
.A1(n_1666),
.A2(n_1637),
.B1(n_1648),
.B2(n_1652),
.C1(n_1636),
.C2(n_1657),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1677),
.A2(n_1637),
.B(n_1648),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1675),
.Y(n_1699)
);

OAI21xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1678),
.A2(n_1662),
.B(n_1672),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1684),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1680),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1684),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1686),
.A2(n_1674),
.B(n_1681),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1687),
.B(n_1663),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1696),
.B(n_1687),
.Y(n_1707)
);

XNOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1693),
.B(n_1451),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1702),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1667),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1695),
.B(n_1685),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1702),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1689),
.B(n_1667),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1698),
.A2(n_1676),
.B(n_1679),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1715),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1690),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1712),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1707),
.B(n_1700),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1709),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1714),
.B(n_1691),
.C(n_1688),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_L g1723 ( 
.A(n_1714),
.B(n_1697),
.C(n_1694),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1708),
.B(n_1682),
.Y(n_1724)
);

OAI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1713),
.A2(n_1701),
.B(n_1699),
.C(n_1692),
.Y(n_1725)
);

NOR2xp67_ASAP7_75t_L g1726 ( 
.A(n_1716),
.B(n_1710),
.Y(n_1726)
);

OAI321xp33_ASAP7_75t_L g1727 ( 
.A1(n_1717),
.A2(n_1711),
.A3(n_1704),
.B1(n_1668),
.B2(n_1660),
.C(n_1635),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1723),
.A2(n_1719),
.B(n_1722),
.C(n_1725),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1718),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1721),
.A2(n_1668),
.B1(n_1636),
.B2(n_1658),
.C(n_1654),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1720),
.A2(n_1658),
.B(n_1652),
.Y(n_1731)
);

AOI211xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1724),
.A2(n_1642),
.B(n_1657),
.C(n_1643),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1728),
.A2(n_1659),
.B(n_1642),
.C(n_1643),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1727),
.A2(n_1659),
.B(n_1660),
.C(n_1653),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1726),
.A2(n_1596),
.B1(n_1599),
.B2(n_1644),
.Y(n_1735)
);

XNOR2xp5_ASAP7_75t_L g1736 ( 
.A(n_1730),
.B(n_1451),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1731),
.A2(n_1660),
.B1(n_1653),
.B2(n_1644),
.C(n_1635),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1729),
.A2(n_1653),
.B1(n_1644),
.B2(n_1635),
.C(n_1603),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1733),
.A2(n_1732),
.B1(n_1596),
.B2(n_1599),
.Y(n_1739)
);

XNOR2xp5_ASAP7_75t_L g1740 ( 
.A(n_1736),
.B(n_1427),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1734),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1735),
.A2(n_1599),
.B1(n_1592),
.B2(n_1593),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1737),
.B(n_1587),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_SL g1744 ( 
.A(n_1741),
.B(n_1738),
.C(n_1610),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1743),
.B(n_1595),
.Y(n_1745)
);

NOR2x1_ASAP7_75t_L g1746 ( 
.A(n_1740),
.B(n_1427),
.Y(n_1746)
);

OAI211xp5_ASAP7_75t_SL g1747 ( 
.A1(n_1746),
.A2(n_1745),
.B(n_1739),
.C(n_1744),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1742),
.B1(n_1602),
.B2(n_1598),
.Y(n_1748)
);

NAND3xp33_ASAP7_75t_L g1749 ( 
.A(n_1748),
.B(n_1610),
.C(n_1603),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1748),
.Y(n_1750)
);

NAND2x1_ASAP7_75t_SL g1751 ( 
.A(n_1750),
.B(n_1602),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1749),
.A2(n_1613),
.B1(n_1610),
.B2(n_1603),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1751),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1752),
.A2(n_1610),
.B(n_1603),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_L g1755 ( 
.A(n_1753),
.B(n_1615),
.C(n_1613),
.Y(n_1755)
);

AOI32xp33_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1754),
.A3(n_1613),
.B1(n_1615),
.B2(n_1619),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1756),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1613),
.B1(n_1615),
.B2(n_1619),
.C(n_1621),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1615),
.B1(n_1619),
.B2(n_1618),
.Y(n_1759)
);


endmodule