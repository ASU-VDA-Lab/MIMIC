module fake_jpeg_10837_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_52),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_49),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_18),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_57),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_63),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_29),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_1),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_90),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_2),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_73),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_3),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_81),
.Y(n_116)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_13),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_87),
.Y(n_102)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_17),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_45),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_21),
.A2(n_30),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_26),
.B(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_10),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_42),
.B1(n_27),
.B2(n_41),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_99),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_34),
.B1(n_41),
.B2(n_40),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_49),
.A2(n_34),
.B1(n_44),
.B2(n_27),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_44),
.B1(n_22),
.B2(n_45),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_43),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_107),
.C(n_117),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_51),
.B(n_37),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_127),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_64),
.A2(n_37),
.B1(n_36),
.B2(n_32),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_122),
.A2(n_129),
.B1(n_131),
.B2(n_141),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_51),
.B(n_36),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_53),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_47),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_135),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_70),
.B(n_7),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_61),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_74),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_130),
.B1(n_126),
.B2(n_109),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_69),
.B(n_11),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_159),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_64),
.C(n_78),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_171),
.C(n_164),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_95),
.A2(n_88),
.B1(n_83),
.B2(n_76),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_89),
.B1(n_86),
.B2(n_85),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_177),
.B1(n_187),
.B2(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_150),
.B(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_56),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_173),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_181),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_88),
.B1(n_50),
.B2(n_54),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_125),
.B1(n_93),
.B2(n_115),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_157),
.A2(n_168),
.B1(n_189),
.B2(n_162),
.Y(n_213)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_12),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_116),
.B(n_60),
.Y(n_160)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_166),
.Y(n_208)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_96),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_93),
.A2(n_115),
.B1(n_105),
.B2(n_94),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_92),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_170),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_100),
.B(n_134),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_132),
.C(n_104),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_126),
.Y(n_172)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_103),
.B(n_111),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_104),
.A2(n_113),
.B(n_94),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_131),
.A2(n_144),
.B(n_112),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_120),
.B(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_139),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_105),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_149),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_141),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_172),
.B1(n_184),
.B2(n_154),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_169),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_191),
.C(n_203),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_210),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_211),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_170),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_173),
.Y(n_230)
);

AOI22x1_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_177),
.B1(n_150),
.B2(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_207),
.B1(n_214),
.B2(n_160),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_167),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_165),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_152),
.B1(n_151),
.B2(n_166),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_148),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_230),
.C(n_247),
.Y(n_248)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_174),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_231),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_145),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_233),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_156),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_176),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_209),
.B(n_215),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_188),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_207),
.A2(n_183),
.B1(n_188),
.B2(n_197),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_246),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_203),
.B(n_204),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_217),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_249),
.A2(n_258),
.B(n_255),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_252),
.C(n_259),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_218),
.B(n_219),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_206),
.C(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_206),
.C(n_205),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_223),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_192),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_199),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_239),
.C(n_224),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_272),
.B1(n_273),
.B2(n_277),
.Y(n_285)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_274),
.C(n_248),
.Y(n_283)
);

AOI221xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_233),
.B1(n_229),
.B2(n_244),
.C(n_224),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_252),
.B(n_206),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_237),
.C(n_238),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_275),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_240),
.B(n_241),
.C(n_227),
.D(n_209),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_249),
.B(n_261),
.Y(n_291)
);

OA21x2_ASAP7_75t_SL g280 ( 
.A1(n_251),
.A2(n_240),
.B(n_232),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_258),
.B1(n_264),
.B2(n_240),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_286),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_253),
.B1(n_261),
.B2(n_248),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_278),
.B1(n_274),
.B2(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_260),
.C(n_253),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_279),
.B(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_299),
.B(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_284),
.C(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_282),
.B1(n_288),
.B2(n_284),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_267),
.B(n_273),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_303),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_302),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_287),
.B(n_289),
.Y(n_303)
);

AOI211xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_257),
.B(n_266),
.C(n_215),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_299),
.B(n_296),
.C(n_257),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.B1(n_304),
.B2(n_196),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_266),
.A3(n_228),
.B1(n_225),
.B2(n_235),
.C1(n_192),
.C2(n_199),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_194),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_309),
.B(n_235),
.C(n_196),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_194),
.C(n_256),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_314),
.Y(n_317)
);


endmodule