module real_jpeg_13527_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_4),
.A2(n_24),
.B1(n_53),
.B2(n_55),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_4),
.B(n_29),
.C(n_32),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_4),
.B(n_30),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_4),
.B(n_39),
.C(n_42),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_4),
.B(n_50),
.C(n_55),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_36),
.B1(n_53),
.B2(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_45),
.B1(n_53),
.B2(n_55),
.Y(n_89)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_75),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_66),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_15),
.B(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_59),
.B2(n_60),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.C(n_46),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_18),
.A2(n_19),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_18),
.A2(n_19),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_18),
.B(n_82),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_18),
.A2(n_19),
.B1(n_94),
.B2(n_95),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_18),
.A2(n_19),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

AOI211xp5_ASAP7_75t_SL g163 ( 
.A1(n_18),
.A2(n_90),
.B(n_111),
.C(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_18),
.A2(n_19),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_18),
.A2(n_94),
.B(n_118),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_18),
.A2(n_19),
.B1(n_67),
.B2(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_67),
.C(n_71),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_47),
.C(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_83),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_25),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_20),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_24),
.B(n_102),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_24),
.B(n_88),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_32),
.B(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_34),
.A2(n_46),
.B1(n_47),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_73),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_41),
.B(n_44),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_41),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OA22x2_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_41),
.Y(n_199)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_42),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_46),
.A2(n_47),
.B1(n_72),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_58),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_56),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_57),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_56),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_56),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_53),
.B(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_67),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_71),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_72),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_231),
.B(n_248),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_129),
.B(n_230),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_112),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_78),
.B(n_112),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_93),
.C(n_104),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_92),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_80),
.A2(n_81),
.B1(n_106),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_80),
.A2(n_81),
.B1(n_143),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_83),
.B1(n_90),
.B2(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_82),
.B(n_147),
.C(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_82),
.A2(n_83),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_83),
.B(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_83),
.B(n_139),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_83),
.A2(n_139),
.B(n_176),
.C(n_181),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_105),
.B(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_85),
.A2(n_90),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_90),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_107),
.B1(n_139),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_90),
.A2(n_139),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_90),
.A2(n_139),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_90),
.A2(n_139),
.B1(n_193),
.B2(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_90),
.B(n_147),
.C(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_90),
.B(n_183),
.C(n_187),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_103),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_110),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_110),
.B(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_128),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_123),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_117),
.B(n_122),
.C(n_128),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_127),
.A2(n_235),
.B1(n_236),
.B2(n_240),
.Y(n_234)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_149),
.B(n_229),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_131),
.B(n_133),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_141),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_227)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_141),
.A2(n_142),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_148),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_148),
.B1(n_158),
.B2(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_178),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_147),
.A2(n_148),
.B1(n_196),
.B2(n_200),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_147),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_147),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_148),
.B(n_209),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_170),
.B(n_223),
.C(n_228),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_153),
.A2(n_154),
.B1(n_176),
.B2(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_217),
.B(n_222),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_189),
.B(n_216),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_212),
.B(n_215),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_201),
.B(n_211),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_240),
.C(n_241),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_247),
.Y(n_250)
);


endmodule