module real_aes_8890_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g548 ( .A1(n_0), .A2(n_152), .B(n_549), .C(n_552), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_1), .B(n_493), .Y(n_553) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g437 ( .A(n_2), .Y(n_437) );
INVx1_ASAP7_75t_L g186 ( .A(n_3), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_4), .B(n_144), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_5), .A2(n_462), .B(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_6), .A2(n_129), .B(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_7), .A2(n_36), .B1(n_138), .B2(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_8), .B(n_129), .Y(n_155) );
AND2x6_ASAP7_75t_L g153 ( .A(n_9), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_10), .A2(n_153), .B(n_452), .C(n_454), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_11), .B(n_37), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_11), .B(n_37), .Y(n_438) );
INVx1_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
INVx1_ASAP7_75t_L g179 ( .A(n_13), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_14), .B(n_142), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_15), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_16), .B(n_144), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_17), .B(n_130), .Y(n_191) );
AO32x2_ASAP7_75t_L g213 ( .A1(n_18), .A2(n_129), .A3(n_159), .B1(n_170), .B2(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_19), .B(n_138), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_20), .B(n_130), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_21), .A2(n_54), .B1(n_138), .B2(n_216), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g238 ( .A1(n_22), .A2(n_81), .B1(n_138), .B2(n_142), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_23), .B(n_138), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_24), .A2(n_170), .B(n_452), .C(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_25), .A2(n_103), .B1(n_112), .B2(n_756), .Y(n_102) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_26), .A2(n_170), .B(n_452), .C(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_27), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_28), .B(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_29), .A2(n_462), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_30), .B(n_172), .Y(n_210) );
INVx2_ASAP7_75t_L g140 ( .A(n_31), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_32), .A2(n_464), .B(n_472), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_33), .B(n_138), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_34), .B(n_172), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_35), .B(n_224), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_38), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_39), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_40), .A2(n_78), .B1(n_115), .B2(n_116), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_40), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_41), .B(n_144), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_42), .B(n_462), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_43), .A2(n_79), .B1(n_432), .B2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_43), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_44), .A2(n_464), .B(n_466), .C(n_472), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_45), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g550 ( .A(n_46), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_47), .A2(n_90), .B1(n_216), .B2(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g467 ( .A(n_48), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_49), .B(n_138), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_50), .B(n_138), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_51), .B(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_51), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_52), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_53), .B(n_150), .Y(n_149) );
AOI22xp33_ASAP7_75t_SL g195 ( .A1(n_55), .A2(n_59), .B1(n_138), .B2(n_142), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_56), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_57), .B(n_138), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_58), .B(n_138), .Y(n_221) );
INVx1_ASAP7_75t_L g154 ( .A(n_60), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_61), .B(n_462), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_62), .B(n_493), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_63), .A2(n_150), .B(n_182), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_64), .B(n_138), .Y(n_187) );
INVx1_ASAP7_75t_L g133 ( .A(n_65), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_66), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_67), .B(n_144), .Y(n_503) );
AO32x2_ASAP7_75t_L g234 ( .A1(n_68), .A2(n_129), .A3(n_170), .B1(n_235), .B2(n_239), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_69), .B(n_145), .Y(n_455) );
INVx1_ASAP7_75t_L g165 ( .A(n_70), .Y(n_165) );
INVx1_ASAP7_75t_L g205 ( .A(n_71), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_72), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_73), .B(n_469), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_74), .A2(n_452), .B(n_472), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_75), .B(n_142), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_76), .Y(n_488) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_78), .Y(n_115) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_79), .A2(n_121), .B1(n_431), .B2(n_432), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_79), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_80), .B(n_468), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_82), .B(n_216), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_83), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_84), .B(n_142), .Y(n_209) );
INVx2_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_86), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_87), .B(n_169), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_88), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
OR2x2_ASAP7_75t_L g435 ( .A(n_89), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g749 ( .A(n_89), .B(n_735), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_91), .A2(n_101), .B1(n_142), .B2(n_143), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_92), .B(n_462), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_93), .Y(n_732) );
INVx1_ASAP7_75t_L g502 ( .A(n_94), .Y(n_502) );
INVxp67_ASAP7_75t_L g491 ( .A(n_95), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_96), .B(n_142), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_97), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g448 ( .A(n_98), .Y(n_448) );
INVx1_ASAP7_75t_L g526 ( .A(n_99), .Y(n_526) );
AND2x2_ASAP7_75t_L g474 ( .A(n_100), .B(n_172), .Y(n_474) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g756 ( .A(n_105), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g725 ( .A(n_108), .B(n_436), .Y(n_725) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_108), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO221x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_736), .B1(n_739), .B2(n_750), .C(n_752), .Y(n_112) );
OAI222xp33_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_117), .B1(n_726), .B2(n_727), .C1(n_732), .C2(n_733), .Y(n_113) );
INVx1_ASAP7_75t_L g726 ( .A(n_114), .Y(n_726) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_433), .B1(n_439), .B2(n_723), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_120), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
INVx2_ASAP7_75t_L g431 ( .A(n_121), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_121), .A2(n_431), .B1(n_742), .B2(n_743), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_355), .Y(n_121) );
AND2x2_ASAP7_75t_SL g122 ( .A(n_123), .B(n_313), .Y(n_122) );
NOR4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_253), .C(n_289), .D(n_303), .Y(n_123) );
OAI221xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_197), .B1(n_229), .B2(n_240), .C(n_244), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_125), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_173), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_156), .Y(n_127) );
AND2x2_ASAP7_75t_L g250 ( .A(n_128), .B(n_157), .Y(n_250) );
INVx3_ASAP7_75t_L g258 ( .A(n_128), .Y(n_258) );
AND2x2_ASAP7_75t_L g312 ( .A(n_128), .B(n_176), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_128), .B(n_175), .Y(n_348) );
AND2x2_ASAP7_75t_L g406 ( .A(n_128), .B(n_268), .Y(n_406) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_135), .B(n_155), .Y(n_128) );
INVx4_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_129), .A2(n_479), .B(n_480), .Y(n_478) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_129), .Y(n_485) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g159 ( .A(n_130), .Y(n_159) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_131), .B(n_132), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_147), .B(n_153), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_144), .Y(n_136) );
INVx3_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_138), .Y(n_528) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g216 ( .A(n_139), .Y(n_216) );
BUFx3_ASAP7_75t_L g237 ( .A(n_139), .Y(n_237) );
AND2x6_ASAP7_75t_L g452 ( .A(n_139), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g143 ( .A(n_140), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
INVx2_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_144), .A2(n_162), .B(n_163), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_SL g203 ( .A1(n_144), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_144), .B(n_491), .Y(n_490) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_145), .A2(n_169), .B1(n_236), .B2(n_238), .Y(n_235) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
INVx1_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
AND2x2_ASAP7_75t_L g450 ( .A(n_146), .B(n_151), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_146), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_152), .Y(n_147) );
INVx2_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_152), .A2(n_166), .B(n_186), .C(n_187), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_152), .A2(n_169), .B1(n_194), .B2(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_152), .A2(n_169), .B1(n_215), .B2(n_217), .Y(n_214) );
BUFx3_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_153), .A2(n_178), .B(n_185), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_153), .A2(n_203), .B(n_207), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_153), .A2(n_220), .B(n_225), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_153), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g462 ( .A(n_153), .B(n_450), .Y(n_462) );
INVx4_ASAP7_75t_SL g473 ( .A(n_153), .Y(n_473) );
AND2x2_ASAP7_75t_L g241 ( .A(n_156), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g255 ( .A(n_156), .B(n_176), .Y(n_255) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_157), .B(n_176), .Y(n_270) );
AND2x2_ASAP7_75t_L g282 ( .A(n_157), .B(n_258), .Y(n_282) );
OR2x2_ASAP7_75t_L g284 ( .A(n_157), .B(n_242), .Y(n_284) );
AND2x2_ASAP7_75t_L g319 ( .A(n_157), .B(n_242), .Y(n_319) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_157), .Y(n_364) );
INVx1_ASAP7_75t_L g372 ( .A(n_157), .Y(n_372) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_171), .Y(n_157) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_158), .A2(n_177), .B(n_188), .Y(n_176) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_159), .B(n_458), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_170), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_168), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_166), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_168), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g551 ( .A(n_169), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_170), .B(n_193), .C(n_196), .Y(n_192) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_172), .A2(n_202), .B(n_210), .Y(n_201) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_172), .A2(n_219), .B(n_228), .Y(n_218) );
INVx2_ASAP7_75t_L g239 ( .A(n_172), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_172), .A2(n_461), .B(n_463), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_172), .A2(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g519 ( .A(n_172), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_173), .A2(n_290), .B1(n_294), .B2(n_298), .C(n_299), .Y(n_289) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g249 ( .A(n_174), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_189), .Y(n_174) );
INVx2_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
AND2x2_ASAP7_75t_L g301 ( .A(n_175), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_175), .B(n_258), .Y(n_320) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g383 ( .A(n_176), .B(n_258), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .C(n_182), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_180), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_180), .A2(n_482), .B(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_182), .A2(n_526), .B(n_527), .C(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_183), .A2(n_208), .B(n_209), .Y(n_207) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g469 ( .A(n_184), .Y(n_469) );
AND2x2_ASAP7_75t_L g305 ( .A(n_189), .B(n_250), .Y(n_305) );
OAI322xp33_ASAP7_75t_L g373 ( .A1(n_189), .A2(n_329), .A3(n_374), .B1(n_376), .B2(n_379), .C1(n_381), .C2(n_385), .Y(n_373) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_190), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g269 ( .A(n_190), .Y(n_269) );
AND2x2_ASAP7_75t_L g378 ( .A(n_190), .B(n_258), .Y(n_378) );
AND2x2_ASAP7_75t_L g410 ( .A(n_190), .B(n_282), .Y(n_410) );
OR2x2_ASAP7_75t_L g413 ( .A(n_190), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g243 ( .A(n_191), .Y(n_243) );
AO21x1_ASAP7_75t_L g242 ( .A1(n_193), .A2(n_196), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_196), .A2(n_447), .B(n_457), .Y(n_446) );
INVx3_ASAP7_75t_L g493 ( .A(n_196), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_196), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_196), .A2(n_523), .B(n_530), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_196), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_211), .Y(n_198) );
INVx1_ASAP7_75t_L g426 ( .A(n_199), .Y(n_426) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g231 ( .A(n_200), .B(n_218), .Y(n_231) );
INVx2_ASAP7_75t_L g266 ( .A(n_200), .Y(n_266) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g288 ( .A(n_201), .Y(n_288) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_201), .Y(n_296) );
OR2x2_ASAP7_75t_L g420 ( .A(n_201), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g245 ( .A(n_211), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g285 ( .A(n_211), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g337 ( .A(n_211), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_218), .Y(n_211) );
AND2x2_ASAP7_75t_L g232 ( .A(n_212), .B(n_233), .Y(n_232) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_212), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g346 ( .A(n_212), .B(n_234), .Y(n_346) );
OR2x2_ASAP7_75t_L g354 ( .A(n_212), .B(n_288), .Y(n_354) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx2_ASAP7_75t_L g263 ( .A(n_213), .Y(n_263) );
AND2x2_ASAP7_75t_L g273 ( .A(n_213), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g297 ( .A(n_213), .B(n_218), .Y(n_297) );
AND2x2_ASAP7_75t_L g361 ( .A(n_213), .B(n_234), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_218), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_218), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g274 ( .A(n_218), .Y(n_274) );
INVx1_ASAP7_75t_L g279 ( .A(n_218), .Y(n_279) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_218), .Y(n_369) );
INVx1_ASAP7_75t_L g421 ( .A(n_218), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g398 ( .A(n_230), .B(n_307), .Y(n_398) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g325 ( .A(n_232), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g424 ( .A(n_232), .B(n_359), .Y(n_424) );
INVx1_ASAP7_75t_L g246 ( .A(n_233), .Y(n_246) );
AND2x2_ASAP7_75t_L g272 ( .A(n_233), .B(n_266), .Y(n_272) );
BUFx2_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_234), .Y(n_252) );
INVx1_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_237), .Y(n_471) );
INVx2_ASAP7_75t_L g552 ( .A(n_237), .Y(n_552) );
INVx1_ASAP7_75t_L g516 ( .A(n_239), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_240), .B(n_247), .Y(n_400) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AOI32xp33_ASAP7_75t_L g244 ( .A1(n_241), .A2(n_245), .A3(n_247), .B1(n_249), .B2(n_251), .Y(n_244) );
AND2x2_ASAP7_75t_L g384 ( .A(n_241), .B(n_257), .Y(n_384) );
AND2x2_ASAP7_75t_L g422 ( .A(n_241), .B(n_320), .Y(n_422) );
INVx1_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_246), .B(n_308), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_247), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_247), .B(n_250), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_247), .B(n_319), .Y(n_401) );
OR2x2_ASAP7_75t_L g415 ( .A(n_247), .B(n_284), .Y(n_415) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g342 ( .A(n_248), .B(n_250), .Y(n_342) );
OR2x2_ASAP7_75t_L g351 ( .A(n_248), .B(n_338), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_250), .B(n_301), .Y(n_323) );
INVx2_ASAP7_75t_L g338 ( .A(n_252), .Y(n_338) );
OR2x2_ASAP7_75t_L g353 ( .A(n_252), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g368 ( .A(n_252), .B(n_369), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_252), .A2(n_345), .B(n_426), .C(n_427), .Y(n_425) );
OAI321xp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_259), .A3(n_264), .B1(n_267), .B2(n_271), .C(n_275), .Y(n_253) );
INVx1_ASAP7_75t_L g366 ( .A(n_254), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g377 ( .A(n_255), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g329 ( .A(n_257), .Y(n_329) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_258), .B(n_372), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_259), .A2(n_397), .B1(n_399), .B2(n_401), .C(n_402), .Y(n_396) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x2_ASAP7_75t_L g334 ( .A(n_261), .B(n_308), .Y(n_334) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_262), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g307 ( .A(n_263), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_264), .A2(n_305), .B(n_350), .C(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g316 ( .A(n_266), .B(n_273), .Y(n_316) );
BUFx2_ASAP7_75t_L g326 ( .A(n_266), .Y(n_326) );
INVx1_ASAP7_75t_L g341 ( .A(n_266), .Y(n_341) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OR2x2_ASAP7_75t_L g347 ( .A(n_269), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g430 ( .A(n_269), .Y(n_430) );
INVx1_ASAP7_75t_L g423 ( .A(n_270), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x2_ASAP7_75t_L g276 ( .A(n_272), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g380 ( .A(n_272), .B(n_297), .Y(n_380) );
INVx1_ASAP7_75t_L g309 ( .A(n_273), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B1(n_283), .B2(n_285), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_277), .B(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g345 ( .A(n_278), .B(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_279), .B(n_288), .Y(n_308) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g300 ( .A(n_282), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g310 ( .A(n_284), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_287), .A2(n_405), .B1(n_407), .B2(n_408), .C(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g293 ( .A(n_288), .Y(n_293) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_288), .Y(n_359) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_291), .B(n_410), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_292), .A2(n_297), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_295), .B(n_305), .Y(n_402) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g371 ( .A(n_296), .Y(n_371) );
AND2x2_ASAP7_75t_L g330 ( .A(n_297), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g419 ( .A(n_297), .Y(n_419) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
INVx1_ASAP7_75t_L g390 ( .A(n_301), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_306), .B1(n_309), .B2(n_310), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_307), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g375 ( .A(n_308), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_308), .B(n_346), .Y(n_412) );
OR2x2_ASAP7_75t_L g385 ( .A(n_309), .B(n_338), .Y(n_385) );
INVx1_ASAP7_75t_L g324 ( .A(n_310), .Y(n_324) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_312), .B(n_363), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_332), .C(n_343), .Y(n_313) );
OAI211xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_321), .C(n_327), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_316), .A2(n_387), .B1(n_391), .B2(n_394), .C(n_396), .Y(n_386) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g328 ( .A(n_319), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g382 ( .A(n_319), .B(n_383), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g367 ( .A1(n_320), .A2(n_368), .B(n_370), .C(n_372), .Y(n_367) );
INVx2_ASAP7_75t_L g414 ( .A(n_320), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g393 ( .A(n_326), .B(n_346), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
OAI21xp5_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_335), .B(n_336), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI21xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B(n_342), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_337), .B(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_342), .B(n_429), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_349), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g370 ( .A(n_346), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND4x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_386), .C(n_403), .D(n_425), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_373), .Y(n_356) );
OAI211xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_362), .B(n_365), .C(n_367), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_361), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_372), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
INVx2_ASAP7_75t_SL g395 ( .A(n_383), .Y(n_395) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g408 ( .A(n_393), .Y(n_408) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_SL g403 ( .A(n_404), .B(n_411), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_413), .B1(n_415), .B2(n_416), .C(n_417), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g729 ( .A(n_434), .Y(n_729) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g735 ( .A(n_436), .Y(n_735) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx2_ASAP7_75t_L g730 ( .A(n_439), .Y(n_730) );
OR3x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_621), .C(n_686), .Y(n_439) );
NAND4xp25_ASAP7_75t_SL g440 ( .A(n_441), .B(n_562), .C(n_588), .D(n_611), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_494), .B1(n_532), .B2(n_539), .C(n_554), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_443), .A2(n_555), .B1(n_579), .B2(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_475), .Y(n_443) );
INVx1_ASAP7_75t_SL g615 ( .A(n_444), .Y(n_615) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_459), .Y(n_444) );
OR2x2_ASAP7_75t_L g537 ( .A(n_445), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g557 ( .A(n_445), .B(n_476), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_445), .B(n_484), .Y(n_570) );
AND2x2_ASAP7_75t_L g587 ( .A(n_445), .B(n_459), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_445), .B(n_535), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_445), .B(n_586), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_445), .B(n_475), .Y(n_708) );
AOI211xp5_ASAP7_75t_SL g719 ( .A1(n_445), .A2(n_625), .B(n_720), .C(n_721), .Y(n_719) );
INVx5_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_446), .B(n_476), .Y(n_591) );
AND2x2_ASAP7_75t_L g594 ( .A(n_446), .B(n_477), .Y(n_594) );
OR2x2_ASAP7_75t_L g639 ( .A(n_446), .B(n_476), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_446), .B(n_484), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_451), .Y(n_447) );
INVx5_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
INVx5_ASAP7_75t_SL g538 ( .A(n_459), .Y(n_538) );
AND2x2_ASAP7_75t_L g556 ( .A(n_459), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_459), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g642 ( .A(n_459), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g674 ( .A(n_459), .B(n_484), .Y(n_674) );
OR2x2_ASAP7_75t_L g680 ( .A(n_459), .B(n_570), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_459), .B(n_630), .Y(n_689) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
BUFx2_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_465), .A2(n_473), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g546 ( .A1(n_465), .A2(n_473), .B(n_547), .C(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .C(n_471), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_468), .A2(n_471), .B(n_502), .C(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_484), .Y(n_475) );
AND2x2_ASAP7_75t_L g571 ( .A(n_476), .B(n_538), .Y(n_571) );
INVx1_ASAP7_75t_SL g584 ( .A(n_476), .Y(n_584) );
OR2x2_ASAP7_75t_L g619 ( .A(n_476), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g625 ( .A(n_476), .B(n_484), .Y(n_625) );
AND2x2_ASAP7_75t_L g683 ( .A(n_476), .B(n_535), .Y(n_683) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_477), .B(n_538), .Y(n_610) );
INVx3_ASAP7_75t_L g535 ( .A(n_484), .Y(n_535) );
OR2x2_ASAP7_75t_L g576 ( .A(n_484), .B(n_538), .Y(n_576) );
AND2x2_ASAP7_75t_L g586 ( .A(n_484), .B(n_584), .Y(n_586) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_484), .Y(n_634) );
AND2x2_ASAP7_75t_L g643 ( .A(n_484), .B(n_557), .Y(n_643) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_492), .Y(n_484) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_493), .A2(n_545), .B(n_553), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_494), .A2(n_660), .B1(n_662), .B2(n_664), .C(n_667), .Y(n_659) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
AND2x2_ASAP7_75t_L g633 ( .A(n_496), .B(n_614), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_496), .B(n_692), .Y(n_696) );
OR2x2_ASAP7_75t_L g717 ( .A(n_496), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_496), .B(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx5_ASAP7_75t_L g564 ( .A(n_497), .Y(n_564) );
AND2x2_ASAP7_75t_L g641 ( .A(n_497), .B(n_508), .Y(n_641) );
AND2x2_ASAP7_75t_L g702 ( .A(n_497), .B(n_581), .Y(n_702) );
AND2x2_ASAP7_75t_L g715 ( .A(n_497), .B(n_535), .Y(n_715) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_520), .Y(n_506) );
AND2x4_ASAP7_75t_L g542 ( .A(n_507), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g560 ( .A(n_507), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
AND2x2_ASAP7_75t_L g636 ( .A(n_507), .B(n_614), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_507), .B(n_564), .Y(n_646) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_507), .Y(n_654) );
AND2x2_ASAP7_75t_L g666 ( .A(n_507), .B(n_544), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_507), .B(n_598), .Y(n_670) );
AND2x2_ASAP7_75t_L g707 ( .A(n_507), .B(n_702), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_507), .B(n_581), .Y(n_718) );
OR2x2_ASAP7_75t_L g720 ( .A(n_507), .B(n_656), .Y(n_720) );
INVx5_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g606 ( .A(n_508), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g616 ( .A(n_508), .B(n_561), .Y(n_616) );
AND2x2_ASAP7_75t_L g628 ( .A(n_508), .B(n_544), .Y(n_628) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_508), .Y(n_658) );
AND2x4_ASAP7_75t_L g692 ( .A(n_508), .B(n_543), .Y(n_692) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_512), .B(n_516), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
BUFx2_ASAP7_75t_L g541 ( .A(n_520), .Y(n_541) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
AND2x2_ASAP7_75t_L g614 ( .A(n_521), .B(n_544), .Y(n_614) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g561 ( .A(n_522), .B(n_544), .Y(n_561) );
BUFx2_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_534), .B(n_615), .Y(n_694) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_535), .B(n_557), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_535), .B(n_538), .Y(n_596) );
AND2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_587), .Y(n_651) );
AOI221xp5_ASAP7_75t_SL g588 ( .A1(n_536), .A2(n_589), .B1(n_597), .B2(n_599), .C(n_603), .Y(n_588) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g583 ( .A(n_537), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g624 ( .A(n_537), .B(n_625), .Y(n_624) );
OAI321xp33_ASAP7_75t_L g631 ( .A1(n_537), .A2(n_590), .A3(n_632), .B1(n_634), .B2(n_635), .C(n_637), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_538), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_541), .B(n_692), .Y(n_710) );
AND2x2_ASAP7_75t_L g597 ( .A(n_542), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_542), .B(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
AND2x2_ASAP7_75t_L g580 ( .A(n_543), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_543), .B(n_655), .Y(n_685) );
INVx1_ASAP7_75t_L g722 ( .A(n_543), .Y(n_722) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B(n_559), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_556), .A2(n_666), .B(n_715), .C(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_557), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_557), .B(n_595), .Y(n_661) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g604 ( .A(n_561), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_561), .B(n_564), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_561), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_561), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_577), .B2(n_582), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g578 ( .A(n_564), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g601 ( .A(n_564), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g613 ( .A(n_564), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_564), .B(n_607), .Y(n_649) );
OR2x2_ASAP7_75t_L g656 ( .A(n_564), .B(n_581), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_564), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g706 ( .A(n_564), .B(n_692), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B1(n_572), .B2(n_574), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g612 ( .A(n_567), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_570), .A2(n_585), .B1(n_653), .B2(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g700 ( .A(n_571), .Y(n_700) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_575), .A2(n_612), .B1(n_615), .B2(n_616), .C(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g590 ( .A(n_576), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_580), .B(n_646), .Y(n_678) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_581), .Y(n_598) );
INVx1_ASAP7_75t_L g602 ( .A(n_581), .Y(n_602) );
NAND2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
AND2x2_ASAP7_75t_L g629 ( .A(n_587), .B(n_630), .Y(n_629) );
NAND2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g673 ( .A(n_594), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_597), .A2(n_623), .B1(n_626), .B2(n_629), .C(n_631), .Y(n_622) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_601), .B(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_608), .Y(n_603) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx16_ASAP7_75t_R g705 ( .A(n_608), .Y(n_705) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g647 ( .A(n_610), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g668 ( .A(n_613), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_613), .B(n_673), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_616), .B(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .C(n_659), .D(n_672), .Y(n_621) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g630 ( .A(n_625), .Y(n_630) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g663 ( .A(n_634), .B(n_639), .Y(n_663) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_644), .C(n_652), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_642), .A2(n_684), .B(n_712), .C(n_719), .Y(n_711) );
INVx1_ASAP7_75t_SL g671 ( .A(n_643), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g675 ( .A(n_649), .Y(n_675) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_655), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_655), .B(n_666), .Y(n_699) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g676 ( .A(n_666), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_671), .Y(n_667) );
INVxp33_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .A3(n_676), .B1(n_677), .B2(n_679), .C1(n_681), .C2(n_684), .Y(n_672) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_704), .C(n_711), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B1(n_693), .B2(n_695), .C(n_697), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g703 ( .A(n_692), .Y(n_703) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .C(n_709), .Y(n_704) );
NAND2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g731 ( .A(n_724), .Y(n_731) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g751 ( .A(n_737), .Y(n_751) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_745), .C(n_748), .Y(n_739) );
INVx1_ASAP7_75t_L g747 ( .A(n_741), .Y(n_747) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g755 ( .A(n_749), .Y(n_755) );
BUFx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
endmodule