module fake_jpeg_28871_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_22),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_35),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_5),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_13),
.B1(n_15),
.B2(n_23),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_12),
.B(n_17),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.C(n_39),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_20),
.B1(n_12),
.B2(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_13),
.B1(n_16),
.B2(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_50),
.B1(n_47),
.B2(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_16),
.B1(n_1),
.B2(n_10),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_65),
.B(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_16),
.A3(n_52),
.B1(n_39),
.B2(n_43),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_70),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_51),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.C(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_46),
.C(n_42),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

XNOR2x1_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_71),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.C(n_77),
.D(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_59),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_79),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_82),
.C(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_92),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_77),
.B(n_58),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_84),
.B(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_96),
.B1(n_66),
.B2(n_88),
.Y(n_97)
);

AOI321xp33_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_81),
.A3(n_61),
.B1(n_60),
.B2(n_51),
.C(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_98),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_99),
.B(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_81),
.C(n_42),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_81),
.Y(n_104)
);


endmodule