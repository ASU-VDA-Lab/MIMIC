module fake_jpeg_5686_n_326 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_51),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_52),
.B1(n_32),
.B2(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_53),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_3),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_5),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_60),
.B1(n_61),
.B2(n_42),
.Y(n_110)
);

NOR4xp25_ASAP7_75t_SL g63 ( 
.A(n_27),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_36),
.B1(n_29),
.B2(n_38),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_67),
.B(n_72),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_17),
.B1(n_36),
.B2(n_28),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_102),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_17),
.B1(n_21),
.B2(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_17),
.B1(n_36),
.B2(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_82),
.B1(n_84),
.B2(n_93),
.Y(n_121)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_78),
.Y(n_117)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_85),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_38),
.B1(n_30),
.B2(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_30),
.B1(n_37),
.B2(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_37),
.B1(n_33),
.B2(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_37),
.B1(n_33),
.B2(n_25),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_43),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_44),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_103),
.B1(n_64),
.B2(n_9),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_107),
.Y(n_140)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_10),
.Y(n_142)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_111),
.A2(n_78),
.B1(n_66),
.B2(n_81),
.Y(n_164)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_120),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_48),
.C(n_58),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_144),
.C(n_119),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_67),
.B(n_76),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_118),
.Y(n_178)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_55),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_79),
.B1(n_101),
.B2(n_85),
.Y(n_158)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_69),
.B(n_6),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_122),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_139),
.Y(n_174)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_127),
.Y(n_153)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_136),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_97),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_16),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_77),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_79),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_144),
.B1(n_101),
.B2(n_106),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_75),
.B(n_16),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_14),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_75),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_159),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_80),
.B(n_92),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_149),
.A2(n_170),
.B(n_143),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_156),
.A2(n_129),
.B1(n_135),
.B2(n_131),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_127),
.B1(n_135),
.B2(n_136),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_89),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_146),
.B1(n_125),
.B2(n_118),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_74),
.B1(n_109),
.B2(n_70),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_86),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_86),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_171),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_169),
.B(n_174),
.Y(n_204)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_125),
.C(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_114),
.B1(n_124),
.B2(n_117),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_178),
.A2(n_141),
.B(n_143),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_172),
.B(n_157),
.Y(n_228)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_136),
.B1(n_120),
.B2(n_111),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_194),
.B1(n_206),
.B2(n_169),
.Y(n_218)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_193),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_143),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_201),
.A2(n_185),
.B1(n_213),
.B2(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_129),
.B1(n_131),
.B2(n_178),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_166),
.B1(n_165),
.B2(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_156),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_212),
.Y(n_238)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_147),
.B(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_182),
.C(n_155),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_220),
.C(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_204),
.C(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_229),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_171),
.B1(n_150),
.B2(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_228),
.A2(n_234),
.B(n_226),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_205),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_157),
.B1(n_181),
.B2(n_188),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_183),
.B(n_197),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_194),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_191),
.C(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_184),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_199),
.B1(n_184),
.B2(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_243),
.C(n_227),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_240),
.B(n_211),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_251),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_185),
.B(n_198),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_187),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_257),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_207),
.B(n_192),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_254),
.B1(n_244),
.B2(n_251),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_189),
.B(n_193),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_239),
.B(n_222),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_220),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_190),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_275),
.B1(n_252),
.B2(n_245),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_238),
.B1(n_217),
.B2(n_231),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_259),
.B1(n_249),
.B2(n_246),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_233),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_282)
);

OAI322xp33_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_219),
.A3(n_216),
.B1(n_218),
.B2(n_221),
.C1(n_238),
.C2(n_235),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_243),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_225),
.B1(n_236),
.B2(n_224),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_224),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_242),
.C(n_248),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_289),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_292),
.B1(n_276),
.B2(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_256),
.B1(n_262),
.B2(n_254),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_279),
.A2(n_262),
.B1(n_245),
.B2(n_258),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_288),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_278),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_302),
.C(n_258),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_300),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_269),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_268),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_287),
.B(n_291),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_305),
.B(n_308),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_272),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_311),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_280),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_286),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_299),
.B(n_292),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.C(n_294),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_295),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_300),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_270),
.B(n_255),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_270),
.Y(n_320)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_320),
.A3(n_322),
.B1(n_312),
.B2(n_315),
.C1(n_303),
.C2(n_290),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_247),
.B(n_253),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_325),
.Y(n_326)
);


endmodule