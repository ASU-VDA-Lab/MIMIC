module fake_jpeg_30152_n_429 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_429);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx10_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_46),
.B(n_83),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_48),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_0),
.CON(n_53),
.SN(n_53)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_76),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_67),
.Y(n_94)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_26),
.B(n_3),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_85),
.Y(n_120)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_87),
.Y(n_129)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_71),
.Y(n_132)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_89),
.B(n_20),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_91),
.B(n_139),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_40),
.B1(n_39),
.B2(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_95),
.A2(n_110),
.B1(n_112),
.B2(n_29),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_32),
.B1(n_36),
.B2(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_97),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_116),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_32),
.B1(n_36),
.B2(n_20),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_63),
.B1(n_61),
.B2(n_70),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_52),
.B(n_34),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_68),
.A2(n_36),
.B1(n_32),
.B2(n_33),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_131),
.B1(n_86),
.B2(n_77),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_34),
.B(n_33),
.C(n_35),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_87),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_36),
.B1(n_35),
.B2(n_20),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_8),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_3),
.C(n_5),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_42),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_85),
.B(n_42),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_42),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_29),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_145),
.B(n_148),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_147),
.A2(n_156),
.B1(n_109),
.B2(n_142),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_66),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_179),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_108),
.B(n_55),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_152),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_84),
.B1(n_59),
.B2(n_73),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_158),
.A2(n_140),
.B1(n_143),
.B2(n_115),
.Y(n_210)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_81),
.C(n_72),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_181),
.Y(n_208)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_106),
.A2(n_69),
.B1(n_50),
.B2(n_29),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_171),
.B1(n_190),
.B2(n_122),
.Y(n_196)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_29),
.B1(n_5),
.B2(n_6),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_118),
.B1(n_116),
.B2(n_113),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_172),
.A2(n_176),
.B1(n_99),
.B2(n_143),
.Y(n_213)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_94),
.A2(n_29),
.B1(n_9),
.B2(n_10),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_177),
.A2(n_187),
.B1(n_194),
.B2(n_99),
.Y(n_232)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_195),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_105),
.Y(n_182)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_101),
.B(n_8),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_183),
.B(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_97),
.B(n_8),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_9),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_94),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_92),
.B(n_9),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_11),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_181),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_11),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_161),
.Y(n_202)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_192),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_129),
.A2(n_96),
.A3(n_130),
.B1(n_144),
.B2(n_135),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_99),
.B(n_117),
.C(n_111),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_94),
.A2(n_12),
.B1(n_130),
.B2(n_138),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_196),
.B(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_202),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_153),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_223),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_210),
.A2(n_140),
.B1(n_155),
.B2(n_142),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_152),
.A2(n_113),
.B1(n_126),
.B2(n_124),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_168),
.B1(n_184),
.B2(n_174),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_218),
.B1(n_190),
.B2(n_189),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_147),
.A2(n_124),
.B1(n_126),
.B2(n_109),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_156),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_135),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_144),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_236),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_156),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_145),
.B(n_105),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_237),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_161),
.B(n_137),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_164),
.C(n_181),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_239),
.A2(n_273),
.B(n_241),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_186),
.B1(n_193),
.B2(n_163),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_157),
.C(n_162),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_257),
.C(n_220),
.Y(n_290)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_255),
.B1(n_262),
.B2(n_234),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_180),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_245),
.B(n_252),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_259),
.B1(n_261),
.B2(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_149),
.B(n_191),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_236),
.B(n_208),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_185),
.C(n_189),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_166),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_156),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_253),
.B(n_254),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_197),
.C(n_200),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_196),
.A2(n_212),
.B1(n_197),
.B2(n_214),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_202),
.B(n_172),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_269),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_178),
.B1(n_169),
.B2(n_195),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_192),
.B1(n_160),
.B2(n_173),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_198),
.B(n_182),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_198),
.B(n_150),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_204),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_175),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_159),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_220),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_228),
.A2(n_154),
.B1(n_90),
.B2(n_111),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_231),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_281),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_214),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_213),
.B(n_218),
.C(n_206),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_270),
.B(n_264),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_245),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_283),
.B(n_290),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_304),
.B1(n_265),
.B2(n_261),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_289),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_238),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_225),
.B1(n_209),
.B2(n_233),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_209),
.B1(n_233),
.B2(n_203),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_241),
.B(n_204),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_256),
.A2(n_117),
.B(n_215),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_304),
.B(n_287),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_269),
.B(n_215),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_243),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_242),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_268),
.Y(n_299)
);

AND2x2_ASAP7_75t_SL g320 ( 
.A(n_299),
.B(n_248),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_242),
.B(n_90),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_257),
.C(n_249),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_260),
.A2(n_203),
.B1(n_229),
.B2(n_117),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_308),
.B1(n_289),
.B2(n_274),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_286),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_254),
.B1(n_267),
.B2(n_271),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_314),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_246),
.B1(n_252),
.B2(n_262),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_310),
.A2(n_326),
.B1(n_328),
.B2(n_279),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_316),
.C(n_330),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_285),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_276),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_249),
.C(n_248),
.Y(n_316)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_250),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_322),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_323),
.Y(n_351)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_332),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_325),
.A2(n_294),
.B(n_301),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_278),
.A2(n_244),
.B1(n_247),
.B2(n_266),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_272),
.B1(n_239),
.B2(n_229),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_239),
.C(n_12),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_280),
.C(n_295),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_291),
.C(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_282),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_333),
.B(n_348),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_329),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_335),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_338),
.B(n_339),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_337),
.A2(n_346),
.B1(n_318),
.B2(n_320),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_300),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_274),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_340),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_301),
.B1(n_277),
.B2(n_300),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_341),
.A2(n_352),
.B1(n_310),
.B2(n_319),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_347),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_275),
.C(n_299),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_354),
.C(n_356),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_299),
.B(n_292),
.Y(n_347)
);

A2O1A1Ixp33_ASAP7_75t_SL g352 ( 
.A1(n_313),
.A2(n_279),
.B(n_305),
.C(n_288),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_305),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_311),
.Y(n_355)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_355),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_302),
.C(n_279),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_374),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_360),
.A2(n_361),
.B1(n_347),
.B2(n_343),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_318),
.B1(n_327),
.B2(n_320),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_334),
.C(n_356),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_366),
.C(n_370),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_312),
.C(n_307),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_373),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_345),
.C(n_316),
.Y(n_370)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_339),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_341),
.A2(n_326),
.B1(n_327),
.B2(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_306),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_367),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_379),
.Y(n_392)
);

FAx1_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_339),
.CI(n_336),
.CON(n_379),
.SN(n_379)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_388),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_360),
.A2(n_343),
.B1(n_344),
.B2(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_383),
.B(n_387),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_348),
.C(n_338),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_389),
.C(n_367),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_336),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_330),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_324),
.C(n_350),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

OAI221xp5_ASAP7_75t_L g393 ( 
.A1(n_385),
.A2(n_371),
.B1(n_364),
.B2(n_362),
.C(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_393),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_395),
.B(n_402),
.Y(n_408)
);

AO221x1_ASAP7_75t_L g399 ( 
.A1(n_391),
.A2(n_352),
.B1(n_374),
.B2(n_362),
.C(n_358),
.Y(n_399)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_399),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_389),
.C(n_386),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_378),
.C(n_388),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_384),
.A2(n_377),
.B(n_363),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_407),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_384),
.B(n_380),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_404),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_409),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_398),
.A2(n_373),
.B1(n_379),
.B2(n_382),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_381),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_401),
.B(n_379),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_410),
.B(n_392),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_392),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_414),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_395),
.C(n_394),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_416),
.A2(n_406),
.B(n_403),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_394),
.Y(n_418)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_418),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_409),
.B(n_404),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_SL g424 ( 
.A(n_419),
.B(n_420),
.C(n_413),
.Y(n_424)
);

NAND4xp25_ASAP7_75t_L g423 ( 
.A(n_421),
.B(n_412),
.C(n_405),
.D(n_415),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_423),
.A2(n_424),
.B(n_411),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_425),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_387),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_426),
.B1(n_352),
.B2(n_279),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_352),
.Y(n_429)
);


endmodule