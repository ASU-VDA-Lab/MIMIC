module fake_jpeg_11425_n_549 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_549);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_549;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_1),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_87),
.Y(n_117)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_65),
.B(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_28),
.B(n_9),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_84),
.Y(n_110)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_28),
.A2(n_7),
.B(n_16),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_27),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_31),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_27),
.B1(n_38),
.B2(n_24),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_6),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_27),
.B(n_17),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_42),
.Y(n_114)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_100),
.Y(n_148)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_17),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_50),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_54),
.C(n_52),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_105),
.A2(n_24),
.B(n_36),
.C(n_38),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_112),
.B(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_113),
.B(n_143),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_114),
.B(n_124),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_24),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_19),
.B1(n_32),
.B2(n_44),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_156),
.B1(n_32),
.B2(n_19),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_39),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_129),
.B(n_130),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_72),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_47),
.B1(n_40),
.B2(n_37),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_132),
.A2(n_32),
.B(n_36),
.Y(n_199)
);

BUFx16f_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_134),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_141),
.A2(n_36),
.B1(n_29),
.B2(n_2),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_48),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_48),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_161),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_83),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_88),
.B1(n_59),
.B2(n_60),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_44),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_56),
.A2(n_42),
.B1(n_40),
.B2(n_19),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_57),
.B(n_50),
.Y(n_161)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_50),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_175),
.Y(n_227)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_169),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_200),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_171),
.A2(n_194),
.B1(n_107),
.B2(n_163),
.Y(n_236)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_173),
.A2(n_174),
.B1(n_190),
.B2(n_203),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_105),
.A2(n_104),
.B1(n_97),
.B2(n_95),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_41),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_41),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_191),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_23),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_182),
.B(n_136),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_94),
.B1(n_91),
.B2(n_90),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_183),
.A2(n_202),
.B1(n_222),
.B2(n_223),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_29),
.B(n_14),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_221),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_186),
.Y(n_277)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_187),
.Y(n_274)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_64),
.B1(n_80),
.B2(n_78),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_41),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_148),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_194),
.B(n_218),
.Y(n_269)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_199),
.A2(n_184),
.B(n_210),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_116),
.A2(n_82),
.B1(n_70),
.B2(n_23),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_132),
.A2(n_25),
.B1(n_40),
.B2(n_42),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_120),
.B(n_0),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_211),
.Y(n_245)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_142),
.B(n_25),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_215),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_151),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_142),
.B(n_38),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_219),
.Y(n_230)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_138),
.A2(n_29),
.B1(n_10),
.B2(n_11),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_139),
.A2(n_29),
.B1(n_10),
.B2(n_11),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_151),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_225),
.Y(n_270)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_192),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_234),
.B(n_0),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_168),
.B(n_149),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_271),
.C(n_211),
.Y(n_280)
);

AOI22x1_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_122),
.B1(n_165),
.B2(n_135),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_247),
.A2(n_266),
.B(n_5),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_175),
.A2(n_111),
.B(n_149),
.C(n_108),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_207),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_167),
.A2(n_163),
.B1(n_118),
.B2(n_135),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_204),
.B1(n_188),
.B2(n_181),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_252),
.A2(n_6),
.B(n_16),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_178),
.B(n_165),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_255),
.B(n_259),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_187),
.A2(n_158),
.B1(n_140),
.B2(n_108),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_177),
.B(n_128),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_257),
.B(n_216),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_191),
.B(n_128),
.Y(n_259)
);

AOI22x1_ASAP7_75t_SL g266 ( 
.A1(n_199),
.A2(n_152),
.B1(n_155),
.B2(n_164),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_184),
.A2(n_118),
.B1(n_160),
.B2(n_152),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_273),
.B1(n_275),
.B2(n_247),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_206),
.B(n_158),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_215),
.A2(n_160),
.B1(n_107),
.B2(n_155),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_164),
.B1(n_157),
.B2(n_11),
.Y(n_275)
);

AO22x1_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_211),
.B1(n_221),
.B2(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_278),
.B(n_289),
.Y(n_338)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_180),
.A3(n_185),
.B1(n_201),
.B2(n_211),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_279),
.A2(n_304),
.B(n_306),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_280),
.B(n_313),
.Y(n_355)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_282),
.A2(n_301),
.B1(n_320),
.B2(n_258),
.Y(n_349)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_214),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_284),
.B(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_265),
.Y(n_285)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_285),
.A2(n_287),
.B(n_311),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_231),
.B(n_196),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_288),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_209),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_SL g290 ( 
.A(n_251),
.B(n_213),
.C(n_212),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_300),
.C(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_232),
.Y(n_293)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_298),
.A2(n_302),
.B1(n_1),
.B2(n_2),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_225),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_308),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_227),
.C(n_252),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_235),
.B1(n_226),
.B2(n_227),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_240),
.A2(n_249),
.B1(n_263),
.B2(n_245),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_230),
.B(n_197),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_307),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_245),
.A2(n_172),
.B1(n_208),
.B2(n_198),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g306 ( 
.A1(n_235),
.A2(n_195),
.B(n_166),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_245),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_176),
.Y(n_308)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_169),
.C(n_157),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_240),
.A2(n_193),
.B1(n_179),
.B2(n_216),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_243),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_314),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_261),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_228),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_238),
.B(n_6),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_321),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_318),
.A2(n_324),
.B(n_250),
.Y(n_333)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_273),
.A2(n_268),
.B1(n_275),
.B2(n_248),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_262),
.B(n_5),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_262),
.A2(n_0),
.B(n_1),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_322),
.A2(n_325),
.B(n_258),
.Y(n_346)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_323),
.A2(n_260),
.B1(n_254),
.B2(n_229),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_264),
.A2(n_6),
.B1(n_14),
.B2(n_12),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_331),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_264),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_334),
.C(n_335),
.Y(n_379)
);

OAI32xp33_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_267),
.A3(n_274),
.B1(n_228),
.B2(n_265),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_342),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_322),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_242),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_267),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_306),
.A2(n_250),
.B(n_277),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_336),
.A2(n_337),
.B(n_346),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_306),
.A2(n_308),
.B(n_307),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_354),
.C(n_366),
.Y(n_389)
);

AO22x1_ASAP7_75t_SL g342 ( 
.A1(n_278),
.A2(n_302),
.B1(n_282),
.B2(n_320),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_301),
.A2(n_239),
.B1(n_274),
.B2(n_276),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_357),
.B1(n_365),
.B2(n_317),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_1),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_306),
.A2(n_239),
.B1(n_229),
.B2(n_276),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_260),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_284),
.A2(n_254),
.B1(n_2),
.B2(n_3),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_290),
.A2(n_11),
.B(n_12),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_361),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_312),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_339),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_17),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_348),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_369),
.Y(n_410)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_374),
.A2(n_383),
.B1(n_393),
.B2(n_394),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_349),
.A2(n_297),
.B1(n_304),
.B2(n_278),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_376),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_338),
.A2(n_297),
.B1(n_278),
.B2(n_291),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_330),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_385),
.Y(n_423)
);

OA22x2_ASAP7_75t_L g380 ( 
.A1(n_351),
.A2(n_325),
.B1(n_298),
.B2(n_281),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_380),
.B(n_391),
.Y(n_436)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_382),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_352),
.A2(n_317),
.B1(n_279),
.B2(n_285),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_313),
.C(n_318),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_395),
.C(n_355),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_358),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_339),
.Y(n_386)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_314),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_392),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_338),
.A2(n_283),
.B1(n_323),
.B2(n_309),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_342),
.A2(n_324),
.B1(n_296),
.B2(n_294),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_293),
.C(n_305),
.Y(n_395)
);

AO22x2_ASAP7_75t_L g396 ( 
.A1(n_342),
.A2(n_292),
.B1(n_295),
.B2(n_319),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_396),
.A2(n_364),
.B1(n_362),
.B2(n_353),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_356),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_397),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_367),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_398),
.A2(n_399),
.B1(n_404),
.B2(n_332),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_343),
.A2(n_296),
.B1(n_2),
.B2(n_3),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_359),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_401),
.A2(n_361),
.B(n_346),
.Y(n_416)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_402),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_403),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_365),
.A2(n_4),
.B1(n_363),
.B2(n_329),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_327),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_412),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_425),
.C(n_426),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_379),
.B(n_355),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_413),
.A2(n_427),
.B1(n_375),
.B2(n_394),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_388),
.A2(n_337),
.B(n_329),
.Y(n_415)
);

XOR2x2_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_421),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_416),
.B(n_400),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_389),
.B(n_340),
.Y(n_421)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_334),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_363),
.C(n_366),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_372),
.A2(n_328),
.B1(n_336),
.B2(n_333),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_391),
.C(n_377),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_430),
.C(n_431),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_376),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_388),
.B(n_368),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_371),
.A2(n_332),
.B(n_368),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_432),
.A2(n_400),
.B(n_401),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_383),
.B(n_372),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_380),
.C(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_369),
.Y(n_438)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_438),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_404),
.B1(n_371),
.B2(n_374),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_439),
.A2(n_449),
.B1(n_460),
.B2(n_434),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_451),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_441),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_410),
.Y(n_442)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_443),
.A2(n_444),
.B1(n_445),
.B2(n_452),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_410),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_413),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_414),
.A2(n_393),
.B1(n_396),
.B2(n_380),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_422),
.Y(n_450)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_396),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_419),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_390),
.Y(n_455)
);

AOI31xp33_ASAP7_75t_L g468 ( 
.A1(n_455),
.A2(n_438),
.A3(n_442),
.B(n_444),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_418),
.A2(n_396),
.B1(n_380),
.B2(n_387),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_456),
.A2(n_458),
.B1(n_461),
.B2(n_463),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_381),
.C(n_370),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_459),
.C(n_426),
.Y(n_472)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_405),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_412),
.B(n_411),
.C(n_425),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_433),
.A2(n_396),
.B1(n_399),
.B2(n_373),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_405),
.Y(n_461)
);

NOR2x1_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_357),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_409),
.B(n_428),
.C(n_419),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_423),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_421),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_465),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_429),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_427),
.B1(n_436),
.B2(n_435),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_467),
.A2(n_475),
.B1(n_479),
.B2(n_443),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_468),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_436),
.B(n_415),
.C(n_432),
.Y(n_471)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_478),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_430),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_476),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_416),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_417),
.C(n_428),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_484),
.C(n_448),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_446),
.A2(n_449),
.B1(n_460),
.B2(n_445),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_483),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_409),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_417),
.C(n_434),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_486),
.Y(n_513)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_487),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_488),
.A2(n_495),
.B(n_437),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_483),
.B(n_437),
.C(n_453),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_489),
.B(n_490),
.Y(n_512)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_469),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_437),
.C(n_446),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_472),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_420),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_497),
.A2(n_498),
.B1(n_499),
.B2(n_501),
.Y(n_505)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_482),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_474),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_507),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_481),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_510),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_465),
.C(n_476),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_515),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_479),
.Y(n_510)
);

OAI321xp33_ASAP7_75t_L g511 ( 
.A1(n_492),
.A2(n_452),
.A3(n_450),
.B1(n_440),
.B2(n_461),
.C(n_458),
.Y(n_511)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_511),
.Y(n_523)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_514),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_500),
.A2(n_467),
.B1(n_480),
.B2(n_456),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_517),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_464),
.C(n_469),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_471),
.C(n_441),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_510),
.C(n_496),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_513),
.A2(n_492),
.B1(n_486),
.B2(n_494),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_519),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_520),
.B(n_521),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_502),
.C(n_491),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_493),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_512),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_513),
.A2(n_462),
.B1(n_502),
.B2(n_463),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_514),
.C(n_517),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_531),
.A2(n_532),
.B(n_535),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_527),
.B(n_509),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_505),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_520),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_523),
.B(n_506),
.Y(n_535)
);

MAJx2_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_521),
.C(n_508),
.Y(n_540)
);

O2A1O1Ixp33_ASAP7_75t_SL g541 ( 
.A1(n_537),
.A2(n_538),
.B(n_540),
.C(n_533),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_530),
.A2(n_524),
.B(n_528),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_541),
.A2(n_542),
.B(n_543),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_539),
.A2(n_533),
.B(n_519),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_539),
.A2(n_529),
.B(n_526),
.Y(n_543)
);

OAI311xp33_ASAP7_75t_L g545 ( 
.A1(n_542),
.A2(n_462),
.A3(n_522),
.B1(n_407),
.C1(n_392),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_407),
.B(n_347),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_544),
.B(n_347),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_547),
.B(n_345),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_353),
.Y(n_549)
);


endmodule