module fake_jpeg_19824_n_263 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_29),
.Y(n_68)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_23),
.B1(n_33),
.B2(n_20),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_49),
.B1(n_65),
.B2(n_18),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_23),
.B1(n_33),
.B2(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_58),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_61),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_21),
.C(n_18),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_21),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_35),
.B(n_25),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_70),
.B(n_39),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_22),
.B1(n_29),
.B2(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_26),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_73),
.B(n_79),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_74),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_79),
.B1(n_87),
.B2(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_91),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_19),
.B1(n_43),
.B2(n_36),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_21),
.B(n_38),
.C(n_17),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_104),
.B(n_35),
.C(n_25),
.Y(n_121)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_38),
.B1(n_56),
.B2(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_52),
.Y(n_131)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_17),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_17),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_52),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_16),
.C(n_15),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_19),
.B1(n_43),
.B2(n_50),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_43),
.A3(n_50),
.B1(n_19),
.B2(n_17),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_98),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_76),
.B1(n_71),
.B2(n_94),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_97),
.B(n_72),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_42),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_120),
.C(n_131),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_25),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_28),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_35),
.C(n_25),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_44),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_82),
.B1(n_85),
.B2(n_89),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_114),
.B1(n_116),
.B2(n_125),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_92),
.B1(n_80),
.B2(n_100),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_144),
.B1(n_149),
.B2(n_127),
.Y(n_182)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_140),
.B(n_141),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_76),
.B(n_72),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_156),
.B(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_148),
.Y(n_177)
);

AND2x4_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_42),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_145),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_41),
.B1(n_44),
.B2(n_42),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_16),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_81),
.B1(n_77),
.B2(n_41),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_32),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_41),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_1),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_R g163 ( 
.A(n_154),
.B(n_111),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_35),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_141),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_35),
.B1(n_25),
.B2(n_32),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_28),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_115),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_28),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_146),
.C(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_165),
.B1(n_182),
.B2(n_141),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_184),
.C(n_172),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_108),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_183),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_128),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_145),
.B1(n_143),
.B2(n_125),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_116),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_124),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_139),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_152),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_192),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_143),
.B1(n_135),
.B2(n_136),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_193),
.B1(n_166),
.B2(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_173),
.B1(n_182),
.B2(n_181),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_137),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_202),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_169),
.B1(n_165),
.B2(n_174),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_201),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_154),
.A3(n_149),
.B1(n_156),
.B2(n_26),
.C1(n_124),
.C2(n_74),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_1),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_177),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_177),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_220),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_212),
.B1(n_190),
.B2(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_215),
.B1(n_202),
.B2(n_192),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_166),
.B1(n_163),
.B2(n_170),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_204),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_166),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

OA21x2_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_2),
.B(n_3),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_5),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_3),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_228),
.B1(n_220),
.B2(n_209),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_224),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_194),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_196),
.B(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_226),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_201),
.B1(n_186),
.B2(n_198),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_208),
.B1(n_6),
.B2(n_7),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_219),
.B(n_215),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_231),
.B(n_7),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_208),
.B(n_216),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_221),
.B(n_223),
.C(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.C(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_5),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_236),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_6),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_241),
.C(n_240),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_251),
.B(n_7),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_235),
.B(n_234),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_233),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_246),
.C(n_9),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

A2O1A1O1Ixp25_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_9),
.B(n_10),
.C(n_12),
.D(n_244),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_257),
.C(n_258),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_259),
.B(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_10),
.Y(n_263)
);


endmodule