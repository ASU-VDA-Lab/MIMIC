module real_jpeg_21666_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_0),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_0),
.A2(n_25),
.B1(n_46),
.B2(n_47),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_1),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_35),
.B1(n_86),
.B2(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_5),
.A2(n_28),
.B1(n_31),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_6),
.B(n_78),
.Y(n_140)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_13),
.B(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_13),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_13),
.A2(n_24),
.B(n_42),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_84),
.B1(n_86),
.B2(n_114),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_13),
.A2(n_31),
.B(n_55),
.C(n_63),
.D(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_31),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_13),
.B(n_27),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_91),
.B(n_140),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_23),
.B(n_36),
.C(n_70),
.D(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_120),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_18),
.B(n_79),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_53),
.C(n_66),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_19),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_38),
.B2(n_52),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_39),
.C(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_32),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_22),
.A2(n_26),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_27),
.B(n_29),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_26),
.B(n_34),
.Y(n_168)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_28),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_37),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_29),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_40),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_41),
.A2(n_43),
.B(n_86),
.C(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_43),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_45),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_47),
.B1(n_56),
.B2(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_46),
.B(n_56),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_46),
.B(n_157),
.Y(n_156)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_47),
.A2(n_57),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_53),
.A2(n_66),
.B1(n_67),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_53),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_60),
.B(n_62),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_54),
.A2(n_60),
.B1(n_64),
.B2(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_55),
.B(n_103),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_64),
.A2(n_102),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_64),
.B(n_84),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_68),
.B(n_72),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_74),
.A2(n_77),
.B(n_145),
.Y(n_153)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_76),
.B(n_84),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_98),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_91),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_109),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_174),
.B(n_179),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_161),
.B(n_173),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_141),
.B(n_160),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.C(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_150),
.B(n_159),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_148),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_154),
.B(n_158),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_153),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_171),
.B2(n_172),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_175),
.B(n_176),
.Y(n_179)
);


endmodule