module fake_jpeg_11786_n_293 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_67),
.Y(n_94)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_74),
.Y(n_96)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_79),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_24),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_81),
.Y(n_105)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_83),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_25),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_109),
.B1(n_124),
.B2(n_127),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_46),
.B1(n_28),
.B2(n_25),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_89),
.A2(n_124),
.B1(n_127),
.B2(n_110),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_29),
.C(n_43),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_131),
.C(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_111),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_44),
.B1(n_28),
.B2(n_40),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_43),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_122),
.Y(n_146)
);

AND2x4_ASAP7_75t_SL g115 ( 
.A(n_70),
.B(n_79),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_40),
.B1(n_38),
.B2(n_33),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_128),
.B1(n_131),
.B2(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_38),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_52),
.A2(n_33),
.B1(n_27),
.B2(n_5),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_53),
.A2(n_27),
.B1(n_3),
.B2(n_5),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_9),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_60),
.A2(n_12),
.B1(n_2),
.B2(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_133),
.B1(n_110),
.B2(n_94),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_2),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_100),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_10),
.B1(n_12),
.B2(n_83),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_54),
.B(n_85),
.C(n_76),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_153),
.B1(n_127),
.B2(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_157),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_115),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_151),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_121),
.B1(n_92),
.B2(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_155),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_115),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_159),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_97),
.B(n_133),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_162),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_97),
.B(n_123),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_167),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_136),
.B1(n_150),
.B2(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_94),
.B(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_172),
.Y(n_199)
);

NOR2x1_ASAP7_75t_R g189 ( 
.A(n_169),
.B(n_175),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_118),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_145),
.B1(n_141),
.B2(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_195),
.B1(n_177),
.B2(n_186),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_138),
.B1(n_151),
.B2(n_147),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_148),
.C(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_198),
.C(n_207),
.Y(n_210)
);

AOI22x1_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_135),
.B1(n_152),
.B2(n_157),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_173),
.B1(n_163),
.B2(n_140),
.Y(n_195)
);

AOI22x1_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_142),
.B1(n_159),
.B2(n_171),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_144),
.B1(n_138),
.B2(n_143),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_144),
.A2(n_138),
.B1(n_143),
.B2(n_150),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_148),
.C(n_151),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_227),
.B1(n_195),
.B2(n_192),
.Y(n_239)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_198),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_193),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_188),
.B(n_190),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_229),
.B(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_185),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_206),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_228),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_183),
.B(n_199),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_226),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_182),
.A2(n_194),
.B1(n_180),
.B2(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_199),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_194),
.B(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_235),
.B(n_241),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_189),
.B(n_203),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_245),
.B1(n_215),
.B2(n_217),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_184),
.B(n_176),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_209),
.A2(n_176),
.B1(n_184),
.B2(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_212),
.B1(n_227),
.B2(n_221),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_223),
.C(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_253),
.C(n_258),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_215),
.B1(n_217),
.B2(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_256),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_210),
.C(n_228),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_226),
.B1(n_229),
.B2(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_211),
.B1(n_214),
.B2(n_232),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_216),
.C(n_213),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OA21x2_ASAP7_75t_SL g266 ( 
.A1(n_250),
.A2(n_243),
.B(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_269),
.C(n_254),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_233),
.C(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_272),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_259),
.B(n_257),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_276),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_268),
.A2(n_257),
.B1(n_249),
.B2(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_267),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_264),
.B(n_273),
.Y(n_284)
);

NAND4xp25_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_236),
.C(n_276),
.D(n_272),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_284),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

OAI21x1_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_262),
.B(n_263),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_286),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_246),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_289),
.B(n_264),
.CI(n_275),
.CON(n_290),
.SN(n_290)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_291),
.C(n_288),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_281),
.Y(n_293)
);


endmodule