module fake_jpeg_19897_n_184 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_6),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_21),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_32),
.B1(n_26),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_47),
.B1(n_57),
.B2(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_32),
.B1(n_39),
.B2(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_32),
.B1(n_25),
.B2(n_30),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_27),
.C(n_33),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_29),
.B(n_14),
.C(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_64),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_29),
.B(n_42),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_67),
.B(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_24),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_76),
.B1(n_35),
.B2(n_33),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_71),
.B1(n_35),
.B2(n_30),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_52),
.B(n_37),
.C(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_33),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_33),
.B1(n_25),
.B2(n_44),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_15),
.B(n_17),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_44),
.B(n_25),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_78),
.B(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_24),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_65),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_85),
.B1(n_67),
.B2(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_89),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_91),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_50),
.B1(n_48),
.B2(n_28),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_17),
.B(n_15),
.C(n_14),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_77),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_28),
.B1(n_20),
.B2(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_69),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_36),
.B(n_27),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_92),
.B(n_74),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_104),
.C(n_107),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_108),
.B(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_113),
.B1(n_88),
.B2(n_94),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_67),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_109),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_78),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_123),
.Y(n_137)
);

OA21x2_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_100),
.B(n_112),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_122),
.C(n_1),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_98),
.B1(n_113),
.B2(n_106),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_90),
.B1(n_82),
.B2(n_85),
.C(n_69),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_97),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_129),
.C(n_12),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_62),
.B1(n_13),
.B2(n_19),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_68),
.C(n_12),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_109),
.B(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_136),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2x1_ASAP7_75t_R g135 ( 
.A(n_120),
.B(n_108),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_140),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_0),
.B(n_1),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_11),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_12),
.B1(n_19),
.B2(n_13),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_128),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_129),
.C(n_119),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_127),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_121),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_150),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_131),
.C(n_135),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_114),
.C(n_116),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_134),
.B1(n_152),
.B2(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_155),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_131),
.B(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_159),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_126),
.C(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_126),
.C(n_115),
.Y(n_161)
);

NAND4xp25_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_151),
.C(n_19),
.D(n_4),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_10),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_168),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_171),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_8),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_168),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_177),
.C(n_8),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_167),
.B(n_9),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_173),
.B1(n_169),
.B2(n_10),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_175),
.C(n_9),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_9),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_181),
.Y(n_184)
);


endmodule