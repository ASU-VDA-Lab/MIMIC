module fake_jpeg_23180_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_SL g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_0),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx12_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_1),
.A2(n_3),
.B1(n_2),
.B2(n_4),
.Y(n_13)
);

INVx5_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_24),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_13),
.B1(n_7),
.B2(n_14),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_19),
.A2(n_22),
.B1(n_16),
.B2(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_8),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_7),
.B1(n_15),
.B2(n_12),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_30),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_25),
.C(n_32),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_40),
.Y(n_46)
);

AOI31xp67_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_27),
.A3(n_28),
.B(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_44),
.B2(n_36),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_42),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B(n_27),
.Y(n_51)
);


endmodule