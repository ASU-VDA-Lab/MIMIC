module real_jpeg_6030_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_288;
wire n_78;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_0),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_1),
.Y(n_364)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_1),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g461 ( 
.A(n_1),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_2),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_43),
.B1(n_67),
.B2(n_71),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_3),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_3),
.A2(n_71),
.B1(n_231),
.B2(n_314),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_3),
.A2(n_71),
.B1(n_291),
.B2(n_391),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_3),
.A2(n_71),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_4),
.Y(n_333)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_4),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_5),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_5),
.A2(n_76),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_5),
.A2(n_76),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_5),
.A2(n_76),
.B1(n_441),
.B2(n_443),
.Y(n_440)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_6),
.Y(n_538)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_7),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_7),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_9),
.A2(n_131),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_9),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_9),
.A2(n_256),
.B1(n_281),
.B2(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_9),
.A2(n_281),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g457 ( 
.A1(n_9),
.A2(n_281),
.B1(n_458),
.B2(n_460),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_10),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_42),
.B1(n_54),
.B2(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_12),
.A2(n_57),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_12),
.A2(n_57),
.B1(n_204),
.B2(n_223),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_12),
.A2(n_57),
.B1(n_288),
.B2(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_13),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_13),
.A2(n_167),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_13),
.A2(n_29),
.B1(n_167),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_13),
.A2(n_167),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_14),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_14),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_14),
.A2(n_138),
.B1(n_188),
.B2(n_255),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_14),
.A2(n_188),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_14),
.A2(n_73),
.B1(n_188),
.B2(n_409),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_15),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_15),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_15),
.A2(n_182),
.B1(n_211),
.B2(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_15),
.A2(n_85),
.B1(n_211),
.B2(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_15),
.A2(n_55),
.B1(n_74),
.B2(n_211),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_16),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_16),
.A2(n_50),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_16),
.A2(n_50),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_16),
.A2(n_50),
.B1(n_133),
.B2(n_223),
.Y(n_388)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_18),
.A2(n_141),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_18),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_18),
.B(n_175),
.C(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_18),
.B(n_93),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_18),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_18),
.B(n_136),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_18),
.B(n_269),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_537),
.B(n_539),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_51),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B(n_40),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_24),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_24),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_28),
.Y(n_266)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_28),
.Y(n_273)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_30),
.Y(n_403)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_34),
.A2(n_359),
.B(n_360),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_34),
.B(n_362),
.Y(n_462)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_49),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_51),
.B(n_62),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_58),
.B1(n_66),
.B2(n_72),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_52),
.A2(n_53),
.B1(n_58),
.B2(n_72),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_52),
.A2(n_361),
.B(n_408),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_52),
.A2(n_58),
.B1(n_408),
.B2(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_52),
.A2(n_58),
.B1(n_66),
.B2(n_509),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_SL g359 ( 
.A1(n_54),
.A2(n_160),
.B(n_340),
.Y(n_359)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_58),
.B(n_160),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_58),
.A2(n_429),
.B(n_462),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_146),
.B(n_536),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_142),
.C(n_143),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_63),
.A2(n_64),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.C(n_113),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_65),
.B(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_77),
.A2(n_113),
.B1(n_114),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_77),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_77)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_78),
.A2(n_107),
.B1(n_305),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_78),
.A2(n_107),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_78),
.A2(n_101),
.B1(n_107),
.B2(n_513),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_93),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_80),
.A2(n_268),
.A3(n_285),
.B1(n_288),
.B2(n_290),
.Y(n_284)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_85),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_87),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_89),
.Y(n_294)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_92),
.Y(n_445)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_93),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

AOI22x1_ASAP7_75t_L g430 ( 
.A1(n_93),
.A2(n_144),
.B1(n_309),
.B2(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_93),
.A2(n_144),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_97),
.Y(n_214)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_97),
.Y(n_259)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_102),
.Y(n_371)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_107),
.B(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_107),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_113),
.A2(n_114),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_113),
.B(n_508),
.C(n_511),
.Y(n_519)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_135),
.B(n_137),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_156),
.B(n_161),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_115),
.A2(n_135),
.B1(n_208),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_115),
.A2(n_161),
.B(n_254),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_115),
.A2(n_135),
.B1(n_373),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_116),
.B(n_162),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_116),
.A2(n_136),
.B1(n_390),
.B2(n_393),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_116),
.A2(n_136),
.B1(n_393),
.B2(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_116),
.A2(n_136),
.B1(n_414),
.B2(n_448),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_128),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_127),
.Y(n_292)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_128),
.A2(n_208),
.B(n_215),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_135),
.A2(n_215),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_137),
.Y(n_448)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_140),
.Y(n_374)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_140),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_142),
.B(n_143),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_144),
.A2(n_262),
.B(n_270),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_144),
.B(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_144),
.A2(n_270),
.B(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_530),
.B(n_535),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_501),
.B(n_527),
.Y(n_147)
);

OAI311xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_377),
.A3(n_477),
.B1(n_495),
.C1(n_496),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_319),
.B(n_376),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_296),
.B(n_318),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_248),
.B(n_295),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_218),
.B(n_247),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_179),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_154),
.B(n_179),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_170),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_155),
.A2(n_170),
.B1(n_171),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_159),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_160),
.A2(n_192),
.B(n_198),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_160),
.A2(n_263),
.B(n_267),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_160),
.B(n_331),
.Y(n_340)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_166),
.Y(n_417)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_205),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_180),
.B(n_206),
.C(n_217),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_192),
.B(n_198),
.Y(n_180)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_186),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_192),
.A2(n_343),
.B1(n_344),
.B2(n_347),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_192),
.A2(n_383),
.B1(n_384),
.B2(n_388),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_192),
.A2(n_386),
.B(n_388),
.Y(n_418)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_202),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_236),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_193),
.A2(n_277),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_193),
.A2(n_348),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_201),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_201),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_216),
.B2(n_217),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_240),
.B(n_246),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_228),
.B(n_239),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_224),
.Y(n_352)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_238),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_238),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_237),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_233),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_276),
.B(n_282),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_244),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_250),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_274),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_260),
.B2(n_261),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_260),
.C(n_274),
.Y(n_297)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_258),
.Y(n_392)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_263),
.Y(n_405)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_266),
.Y(n_328)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

INVx4_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_298),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_317),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_302),
.C(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_311),
.C(n_312),
.Y(n_353)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_320),
.B(n_321),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_356),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_322)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_341),
.B2(n_342),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_325),
.B(n_341),
.Y(n_473)
);

OAI32xp33_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_329),
.A3(n_332),
.B1(n_334),
.B2(n_340),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_353),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_353),
.B(n_354),
.C(n_356),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_366),
.B2(n_375),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_357),
.B(n_367),
.C(n_372),
.Y(n_486)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_366),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_372),
.Y(n_366)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_368),
.Y(n_475)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_370),
.Y(n_442)
);

INVx11_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_463),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_SL g496 ( 
.A1(n_378),
.A2(n_463),
.B(n_497),
.C(n_500),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_432),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_379),
.B(n_432),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_411),
.C(n_420),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g476 ( 
.A(n_380),
.B(n_411),
.CI(n_420),
.CON(n_476),
.SN(n_476)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_399),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_400),
.C(n_407),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_389),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_382),
.B(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_SL g396 ( 
.A(n_397),
.Y(n_396)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_407),
.Y(n_399)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_409),
.Y(n_459)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_418),
.B2(n_419),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_418),
.Y(n_452)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_418),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_419),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_418),
.A2(n_452),
.B(n_455),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_427),
.C(n_430),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_421),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_424),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_422),
.B(n_424),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_427),
.A2(n_428),
.B1(n_430),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_433),
.B(n_436),
.C(n_450),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_450),
.B2(n_451),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_446),
.B(n_449),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_447),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_440),
.Y(n_513)
);

INVx4_ASAP7_75t_SL g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_449),
.B(n_504),
.C(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_462),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_476),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_476),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_469),
.C(n_470),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_465),
.A2(n_466),
.B1(n_469),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_488),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.C(n_474),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_471),
.A2(n_472),
.B1(n_474),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_474),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_476),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_490),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_498),
.B(n_499),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_487),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_487),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_484),
.C(n_486),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_493),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_485),
.B1(n_486),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_486),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_492),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_516),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_515),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_515),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_508),
.B1(n_510),
.B2(n_514),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_507),
.A2(n_508),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_518),
.C(n_522),
.Y(n_534)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_510),
.Y(n_514)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_516),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_517),
.B(n_526),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_526),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx8_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx13_ASAP7_75t_L g540 ( 
.A(n_538),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);


endmodule