module fake_jpeg_19855_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_27),
.B1(n_15),
.B2(n_19),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_18),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_27),
.B1(n_20),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_45),
.B1(n_26),
.B2(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_15),
.B1(n_19),
.B2(n_25),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_22),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_39),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_20),
.B1(n_24),
.B2(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_17),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_36),
.B1(n_35),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_39),
.B1(n_44),
.B2(n_20),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_36),
.C(n_35),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.C(n_2),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_24),
.C(n_17),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_45),
.B(n_41),
.C(n_39),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_72),
.B(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_44),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_63),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_81),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_60),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_3),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_79),
.B(n_72),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_49),
.C(n_59),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_104),
.B(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_73),
.B1(n_66),
.B2(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_92),
.B1(n_86),
.B2(n_91),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_85),
.C(n_92),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_70),
.A3(n_81),
.B1(n_11),
.B2(n_8),
.C1(n_9),
.C2(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_75),
.B(n_67),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_8),
.C(n_9),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_92),
.B1(n_93),
.B2(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp67_ASAP7_75t_SL g114 ( 
.A(n_111),
.B(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_99),
.B(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_103),
.B(n_97),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_60),
.B(n_64),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_106),
.B1(n_109),
.B2(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_4),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_106),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_114),
.C(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_123),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_121),
.B(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_5),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_5),
.B(n_6),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_5),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_128),
.B(n_132),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_7),
.Y(n_135)
);


endmodule