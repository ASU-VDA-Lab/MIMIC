module fake_jpeg_778_n_384 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_384);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_384;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_49),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_55),
.B(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_56),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_7),
.C(n_13),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_78),
.C(n_97),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_6),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_69),
.B(n_72),
.Y(n_141)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_76),
.Y(n_142)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_74),
.Y(n_117)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_26),
.B(n_8),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_37),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g152 ( 
.A(n_79),
.Y(n_152)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_26),
.B(n_8),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_16),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_92),
.Y(n_115)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_16),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_45),
.B(n_11),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_11),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_18),
.B1(n_41),
.B2(n_40),
.Y(n_120)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_41),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_54),
.A2(n_44),
.B1(n_27),
.B2(n_46),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_110),
.A2(n_126),
.B1(n_152),
.B2(n_140),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_30),
.B1(n_23),
.B2(n_42),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_118),
.A2(n_139),
.B1(n_153),
.B2(n_156),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_120),
.A2(n_125),
.B1(n_128),
.B2(n_135),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_65),
.B1(n_52),
.B2(n_66),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_46),
.B1(n_23),
.B2(n_30),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_84),
.B1(n_80),
.B2(n_59),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_133),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_52),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_132),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_41),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_65),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_12),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_137),
.A2(n_146),
.B1(n_148),
.B2(n_150),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_12),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_63),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_5),
.B1(n_79),
.B2(n_91),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_91),
.A2(n_99),
.B1(n_61),
.B2(n_75),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_77),
.B1(n_101),
.B2(n_60),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_49),
.A2(n_93),
.B1(n_87),
.B2(n_100),
.Y(n_153)
);

OR2x2_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_119),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_51),
.A2(n_53),
.B1(n_57),
.B2(n_64),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_67),
.A2(n_19),
.B1(n_38),
.B2(n_35),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_103),
.B(n_58),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_166),
.B(n_167),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_58),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_169),
.B(n_178),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_112),
.CI(n_150),
.CON(n_170),
.SN(n_170)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_170),
.B(n_177),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_111),
.B(n_113),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_174),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_132),
.C(n_112),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

BUFx4f_ASAP7_75t_SL g211 ( 
.A(n_175),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_147),
.B(n_114),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_176),
.A2(n_195),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_123),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_105),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_107),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_184),
.Y(n_239)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_192),
.B1(n_193),
.B2(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_106),
.B(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_117),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_191),
.Y(n_217)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_111),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_189),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_108),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_136),
.A2(n_160),
.B1(n_140),
.B2(n_104),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_134),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_196),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_119),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_144),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_120),
.B1(n_153),
.B2(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_207),
.B1(n_183),
.B2(n_199),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_113),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_209),
.B1(n_124),
.B2(n_199),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_157),
.B1(n_154),
.B2(n_109),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_135),
.A2(n_137),
.B1(n_163),
.B2(n_148),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_183),
.B1(n_190),
.B2(n_166),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_146),
.B(n_109),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_130),
.A2(n_110),
.B1(n_126),
.B2(n_82),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_124),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_219),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_218),
.B1(n_205),
.B2(n_174),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_233),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_165),
.A2(n_169),
.B1(n_178),
.B2(n_179),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_203),
.B1(n_168),
.B2(n_165),
.Y(n_219)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_200),
.B1(n_206),
.B2(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_231),
.B1(n_198),
.B2(n_202),
.Y(n_263)
);

CKINVDCx12_ASAP7_75t_R g230 ( 
.A(n_201),
.Y(n_230)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_170),
.B(n_176),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_246),
.Y(n_270)
);

AO22x1_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_173),
.B1(n_195),
.B2(n_191),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_220),
.B(n_186),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_195),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_196),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_255),
.Y(n_274)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_239),
.B(n_181),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_171),
.B(n_187),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_261),
.B(n_264),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_177),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_167),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_201),
.B(n_180),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_251),
.B(n_246),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_226),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_188),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_262),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_175),
.B(n_182),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_209),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_225),
.B1(n_210),
.B2(n_223),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_214),
.B(n_237),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_221),
.C(n_215),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_267),
.C(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_221),
.C(n_223),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_219),
.B(n_213),
.C(n_221),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_285),
.B(n_261),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_277),
.B1(n_279),
.B2(n_258),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_219),
.B1(n_240),
.B2(n_212),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_241),
.A2(n_219),
.B1(n_227),
.B2(n_208),
.Y(n_279)
);

XOR2x1_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_227),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_251),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_260),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_220),
.B1(n_236),
.B2(n_216),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_245),
.B1(n_249),
.B2(n_254),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_297),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_244),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_295),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_293),
.B1(n_298),
.B2(n_302),
.Y(n_318)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_250),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_270),
.B(n_248),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_248),
.C(n_259),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_307),
.C(n_275),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_301),
.B(n_273),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_258),
.B1(n_243),
.B2(n_255),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_258),
.B1(n_243),
.B2(n_262),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_282),
.B1(n_274),
.B2(n_270),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_261),
.C(n_243),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_308),
.A2(n_321),
.B(n_269),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_319),
.C(n_301),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_273),
.B1(n_277),
.B2(n_286),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_323),
.B1(n_325),
.B2(n_307),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_281),
.C(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_284),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_284),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_286),
.B1(n_269),
.B2(n_272),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_285),
.B1(n_271),
.B2(n_287),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_291),
.B1(n_294),
.B2(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_297),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_327),
.B(n_330),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_342)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_299),
.C(n_281),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_333),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_314),
.C(n_309),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_304),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_319),
.B(n_269),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_335),
.B(n_336),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_320),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_325),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_323),
.A2(n_305),
.B1(n_283),
.B2(n_303),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_340),
.B(n_308),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_334),
.A2(n_318),
.B1(n_312),
.B2(n_316),
.Y(n_345)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_345),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_326),
.A2(n_321),
.B1(n_317),
.B2(n_310),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_338),
.B1(n_339),
.B2(n_326),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_314),
.C(n_311),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_349),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_308),
.C(n_317),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_351),
.Y(n_365)
);

BUFx4f_ASAP7_75t_SL g351 ( 
.A(n_344),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_341),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_343),
.B(n_328),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_355),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_344),
.B(n_333),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_342),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_351),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_348),
.A2(n_331),
.B(n_339),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_357),
.A2(n_340),
.B(n_324),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_353),
.A2(n_346),
.B1(n_351),
.B2(n_349),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_359),
.B(n_362),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_361),
.Y(n_372)
);

NOR2x1_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_341),
.Y(n_361)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_364),
.A2(n_257),
.B1(n_211),
.B2(n_242),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_366),
.Y(n_370)
);

AO221x1_ASAP7_75t_L g367 ( 
.A1(n_362),
.A2(n_324),
.B1(n_322),
.B2(n_278),
.C(n_242),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_367),
.A2(n_257),
.B1(n_211),
.B2(n_242),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_322),
.C(n_278),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_369),
.B(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_371),
.B(n_363),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_SL g380 ( 
.A(n_373),
.B(n_377),
.C(n_253),
.Y(n_380)
);

AO22x1_ASAP7_75t_L g374 ( 
.A1(n_370),
.A2(n_365),
.B1(n_359),
.B2(n_361),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_374),
.A2(n_368),
.B1(n_369),
.B2(n_257),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_376),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_222),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_378),
.A2(n_380),
.B(n_253),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_382),
.Y(n_383)
);

BUFx24_ASAP7_75t_SL g382 ( 
.A(n_379),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_211),
.Y(n_384)
);


endmodule