module fake_jpeg_6886_n_165 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_33),
.B1(n_24),
.B2(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_39),
.B(n_3),
.Y(n_69)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_20),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_47),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_24),
.B1(n_15),
.B2(n_4),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_51),
.B1(n_65),
.B2(n_68),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_19),
.C(n_27),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_34),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_23),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_19),
.B1(n_27),
.B2(n_22),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_30),
.B1(n_25),
.B2(n_14),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_16),
.B1(n_25),
.B2(n_22),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_14),
.B1(n_20),
.B2(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_69),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_29),
.B1(n_26),
.B2(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_68),
.B1(n_51),
.B2(n_65),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_6),
.B(n_42),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_40),
.B1(n_36),
.B2(n_41),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_66),
.B1(n_64),
.B2(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_87),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_66),
.B(n_57),
.Y(n_98)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_41),
.Y(n_85)
);

OR2x4_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_9),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_94),
.B1(n_73),
.B2(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_47),
.B1(n_62),
.B2(n_70),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_81),
.B(n_74),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_101),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_48),
.B(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_112),
.B1(n_73),
.B2(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_88),
.B1(n_75),
.B2(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_121),
.B(n_109),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_128),
.B1(n_104),
.B2(n_101),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_107),
.B1(n_96),
.B2(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_92),
.B(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_99),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_126),
.B(n_127),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_134),
.B(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_107),
.C(n_92),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_136),
.C(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_101),
.B(n_108),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_101),
.B(n_106),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_108),
.C(n_90),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_117),
.B(n_116),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_139),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_122),
.B1(n_124),
.B2(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_118),
.B1(n_125),
.B2(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_84),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_139),
.C(n_106),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_143),
.C(n_151),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_140),
.C(n_142),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_144),
.B(n_152),
.C(n_141),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_160),
.B(n_161),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_149),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_158),
.A3(n_155),
.B1(n_87),
.B2(n_80),
.C(n_90),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_95),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_162),
.Y(n_165)
);


endmodule