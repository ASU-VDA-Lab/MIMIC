module fake_aes_5444_n_27 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
AND2x6_ASAP7_75t_L g15 ( .A(n_9), .B(n_0), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_16), .B(n_0), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_12), .B(n_2), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_14), .B(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OA21x2_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_11), .B(n_17), .Y(n_22) );
AOI31xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_15), .A3(n_7), .B(n_8), .Y(n_23) );
NOR2x1p5_ASAP7_75t_L g24 ( .A(n_23), .B(n_15), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_24), .B(n_5), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
endmodule