module fake_jpeg_18024_n_183 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_6),
.B(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NOR2x1_ASAP7_75t_R g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_33),
.B1(n_21),
.B2(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_33),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_20),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_28),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_53),
.C(n_55),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_89),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_41),
.B(n_46),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_76),
.B(n_94),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_41),
.CI(n_30),
.CON(n_69),
.SN(n_69)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_88),
.Y(n_102)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_75),
.B1(n_83),
.B2(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_62),
.B1(n_58),
.B2(n_45),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_87),
.B1(n_95),
.B2(n_23),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_29),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_26),
.B1(n_37),
.B2(n_23),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_37),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_37),
.C(n_34),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_2),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_54),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_29),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_26),
.B(n_23),
.C(n_17),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_76),
.B1(n_24),
.B2(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_106),
.B1(n_109),
.B2(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_24),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_114),
.CI(n_117),
.CON(n_122),
.SN(n_122)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_17),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_17),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_88),
.C(n_89),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_135),
.C(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_94),
.B1(n_87),
.B2(n_67),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_94),
.B1(n_78),
.B2(n_72),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_100),
.B1(n_117),
.B2(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_94),
.B1(n_78),
.B2(n_70),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_73),
.B(n_69),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_133),
.B(n_111),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_84),
.B(n_72),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_99),
.B(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_99),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_81),
.B(n_83),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_81),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_137),
.B1(n_96),
.B2(n_98),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_71),
.B1(n_74),
.B2(n_29),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.C(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_115),
.C(n_107),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_145),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_115),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_129),
.C(n_130),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_128),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_96),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_112),
.C(n_103),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_135),
.C(n_123),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_144),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_139),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_136),
.C(n_137),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_157),
.B1(n_4),
.B2(n_5),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_145),
.CI(n_141),
.CON(n_164),
.SN(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_150),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_169),
.B(n_157),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_151),
.Y(n_169)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.C(n_165),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_162),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_170),
.B1(n_164),
.B2(n_167),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_15),
.B1(n_14),
.B2(n_7),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_176),
.A2(n_4),
.B(n_6),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_177),
.B(n_180),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_10),
.Y(n_183)
);


endmodule