module fake_jpeg_13854_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_43;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_4),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_7),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_15),
.B1(n_7),
.B2(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_21),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_20),
.B(n_17),
.Y(n_36)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_36),
.B1(n_26),
.B2(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_19),
.C(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AO221x1_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_31),
.B2(n_25),
.C(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_27),
.B1(n_30),
.B2(n_25),
.Y(n_40)
);

OAI321xp33_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_31),
.A3(n_35),
.B1(n_16),
.B2(n_17),
.C(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_29),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_28),
.C(n_29),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_34),
.B(n_29),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_29),
.C(n_34),
.Y(n_50)
);


endmodule