module real_jpeg_22100_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_244;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_0),
.A2(n_10),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_0),
.A2(n_35),
.B1(n_66),
.B2(n_71),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_0),
.A2(n_35),
.B1(n_38),
.B2(n_43),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_1),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_44),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_10),
.B1(n_28),
.B2(n_44),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_69),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_10),
.B(n_14),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_38),
.B1(n_43),
.B2(n_122),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_80),
.B1(n_99),
.B2(n_195),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_168),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_53),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_53),
.B(n_219),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_66),
.B1(n_71),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_4),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_107),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_10),
.B1(n_28),
.B2(n_107),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_38),
.B1(n_43),
.B2(n_107),
.Y(n_210)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_65),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_7),
.A2(n_66),
.B1(n_71),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_7),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_133),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_7),
.A2(n_38),
.B1(n_43),
.B2(n_133),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_10),
.B1(n_28),
.B2(n_133),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_28),
.Y(n_30)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_9),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_9),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_72),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_9),
.A2(n_10),
.B1(n_28),
.B2(n_72),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_9),
.A2(n_38),
.B1(n_43),
.B2(n_72),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_10),
.A2(n_11),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_14),
.B1(n_28),
.B2(n_41),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_13),
.B1(n_28),
.B2(n_46),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_29),
.B1(n_38),
.B2(n_43),
.Y(n_84)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_13),
.A2(n_38),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_38),
.Y(n_39)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_136),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_19),
.B(n_109),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_76),
.B2(n_77),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_25),
.A2(n_33),
.B(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_27),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_28),
.B(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_30),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_30),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_30),
.A2(n_34),
.B(n_98),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_31),
.A2(n_80),
.B(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_33),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_33),
.A2(n_80),
.B1(n_179),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_37),
.A2(n_45),
.B(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_37),
.A2(n_83),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_37),
.A2(n_40),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_37),
.A2(n_40),
.B1(n_190),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_37),
.A2(n_40),
.B1(n_210),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_37),
.A2(n_226),
.B(n_241),
.Y(n_240)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_38),
.A2(n_51),
.A3(n_54),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_40),
.A2(n_42),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_40),
.B(n_122),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_41),
.A2(n_43),
.B(n_122),
.C(n_186),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_43),
.B(n_50),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_61),
.B1(n_62),
.B2(n_75),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_55),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_50),
.B(n_53),
.C(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_102),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_49),
.A2(n_57),
.B1(n_127),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_49),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_49),
.A2(n_57),
.B1(n_167),
.B2(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_53),
.Y(n_58)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_53),
.B(n_65),
.Y(n_120)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_54),
.A2(n_68),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_126),
.B(n_128),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_56),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_70),
.B(n_73),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_70),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_63),
.A2(n_106),
.B1(n_108),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_64),
.A2(n_69),
.B1(n_121),
.B2(n_132),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_66),
.B(n_122),
.CON(n_121),
.SN(n_121)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_86),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_80),
.A2(n_96),
.B1(n_99),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_85),
.B(n_146),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_100),
.C(n_104),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_89),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_99),
.B(n_122),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_110),
.Y(n_255)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_116),
.A2(n_117),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.C(n_129),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_129),
.B1(n_130),
.B2(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_170),
.B(n_250),
.C(n_256),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_155),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_138),
.B(n_155),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_151),
.B2(n_154),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_141),
.B(n_142),
.C(n_154),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_150),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_165),
.B(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_249),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_244),
.B(n_248),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_231),
.B(n_243),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_213),
.B(n_230),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_202),
.B(n_212),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_191),
.B(n_201),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_183),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_196),
.B(n_200),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_204),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_209),
.C(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_215),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_221),
.B1(n_228),
.B2(n_229),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_240),
.C(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2x2_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);


endmodule