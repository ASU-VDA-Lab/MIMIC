module fake_jpeg_11748_n_67 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_21),
.A2(n_11),
.B1(n_9),
.B2(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_28),
.Y(n_32)
);

CKINVDCx12_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_4),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_9),
.A3(n_10),
.B1(n_15),
.B2(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_15),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_11),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_26),
.C(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_14),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_43),
.B(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_24),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_39),
.C(n_40),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_9),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_51),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_6),
.C(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_33),
.B1(n_30),
.B2(n_7),
.Y(n_53)
);

OAI321xp33_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_41),
.A3(n_43),
.B1(n_45),
.B2(n_30),
.C(n_5),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_50),
.CI(n_53),
.CON(n_59),
.SN(n_59)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_6),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_55),
.B(n_49),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_54),
.B1(n_50),
.B2(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_54),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_66),
.A2(n_63),
.B(n_65),
.Y(n_67)
);


endmodule