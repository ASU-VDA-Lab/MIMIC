module fake_jpeg_3631_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_58),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_83),
.Y(n_116)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_30),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_82),
.B(n_94),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_0),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_45),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_95),
.Y(n_123)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_23),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_91),
.B(n_46),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_1),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_19),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_102),
.Y(n_142)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_19),
.B(n_3),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_24),
.B1(n_48),
.B2(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_104),
.A2(n_106),
.B1(n_109),
.B2(n_118),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_46),
.B1(n_45),
.B2(n_24),
.Y(n_106)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_83),
.CON(n_107),
.SN(n_107)
);

NAND2x1_ASAP7_75t_SL g170 ( 
.A(n_107),
.B(n_134),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_101),
.B1(n_91),
.B2(n_46),
.Y(n_109)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_24),
.B1(n_46),
.B2(n_48),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_97),
.B1(n_72),
.B2(n_73),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_53),
.A2(n_21),
.B1(n_50),
.B2(n_44),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_21),
.B(n_50),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_119),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_46),
.B1(n_51),
.B2(n_27),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_66),
.A2(n_20),
.B1(n_44),
.B2(n_43),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_129),
.A2(n_136),
.B1(n_139),
.B2(n_152),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_68),
.A2(n_51),
.B1(n_20),
.B2(n_43),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_71),
.A2(n_40),
.B1(n_34),
.B2(n_33),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_147),
.B(n_70),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_87),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_28),
.C(n_27),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_16),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_159),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_92),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_166),
.B(n_172),
.Y(n_238)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_98),
.B1(n_103),
.B2(n_76),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_169),
.A2(n_217),
.B1(n_223),
.B2(n_144),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_76),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_179),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_89),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_173),
.B(n_176),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_174),
.Y(n_235)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g247 ( 
.A(n_175),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_81),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_189),
.Y(n_240)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_105),
.B(n_63),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_180),
.Y(n_258)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_63),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_54),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_54),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_110),
.B(n_52),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_104),
.A2(n_52),
.B1(n_73),
.B2(n_70),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_113),
.B1(n_117),
.B2(n_151),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_77),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_190),
.B(n_194),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_114),
.B(n_3),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_192),
.B(n_210),
.Y(n_255)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_3),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_107),
.B(n_4),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_195),
.B(n_200),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_201),
.Y(n_267)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_5),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_202),
.B(n_208),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_159),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_203),
.A2(n_222),
.B1(n_14),
.B2(n_16),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_114),
.B(n_128),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_211),
.B(n_213),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_130),
.B(n_5),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_220),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_138),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_111),
.B(n_6),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_111),
.B(n_6),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_216),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_115),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_115),
.Y(n_218)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_121),
.B(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_160),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_131),
.C(n_124),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_236),
.C(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_126),
.B1(n_106),
.B2(n_121),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_246),
.B1(n_273),
.B2(n_184),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_170),
.C(n_167),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_251),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_131),
.B(n_117),
.C(n_124),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_244),
.B(n_164),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_120),
.C(n_133),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_192),
.A2(n_151),
.B1(n_153),
.B2(n_120),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_174),
.A2(n_144),
.B(n_153),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_249),
.A2(n_244),
.B(n_251),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_209),
.A2(n_113),
.B1(n_117),
.B2(n_16),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_256),
.A2(n_204),
.B1(n_214),
.B2(n_219),
.Y(n_322)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_257),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_170),
.B(n_14),
.C(n_15),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_260),
.C(n_212),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_14),
.C(n_15),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_174),
.A2(n_14),
.B(n_15),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_217),
.B(n_208),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_199),
.A2(n_201),
.B1(n_208),
.B2(n_164),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_173),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_277),
.B(n_282),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_278),
.A2(n_284),
.B(n_308),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_280),
.A2(n_281),
.B1(n_289),
.B2(n_298),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_255),
.A2(n_239),
.B1(n_224),
.B2(n_273),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_240),
.B(n_195),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_285),
.B(n_291),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_294),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_220),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_288),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_182),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_239),
.A2(n_199),
.B1(n_164),
.B2(n_183),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_179),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_311),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_262),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_305),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_224),
.A2(n_164),
.B1(n_185),
.B2(n_222),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_231),
.A2(n_218),
.B1(n_165),
.B2(n_175),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_322),
.B1(n_248),
.B2(n_258),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_301),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_198),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_316),
.C(n_235),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_234),
.A2(n_168),
.B1(n_181),
.B2(n_200),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_303),
.A2(n_248),
.B1(n_258),
.B2(n_272),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

OAI22x1_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_207),
.B1(n_205),
.B2(n_197),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_178),
.B(n_180),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_228),
.B(n_235),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_309),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_228),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_314),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_231),
.B(n_211),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_176),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_320),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_226),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_315),
.A2(n_278),
.B(n_296),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_229),
.B(n_187),
.C(n_193),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_319),
.Y(n_349)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_241),
.B(n_186),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_314),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_363),
.C(n_313),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_280),
.A2(n_256),
.B1(n_249),
.B2(n_254),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_324),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_302),
.B(n_259),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_362),
.Y(n_375)
);

AO22x1_ASAP7_75t_SL g331 ( 
.A1(n_281),
.A2(n_246),
.B1(n_263),
.B2(n_225),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_298),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_284),
.A2(n_254),
.B1(n_247),
.B2(n_232),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_304),
.A2(n_247),
.B1(n_232),
.B2(n_268),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_304),
.A2(n_268),
.B1(n_230),
.B2(n_263),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_340),
.A2(n_358),
.B(n_360),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_304),
.A2(n_230),
.B1(n_233),
.B2(n_227),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_343),
.A2(n_361),
.B1(n_345),
.B2(n_352),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_308),
.Y(n_345)
);

INVx13_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

AO21x2_ASAP7_75t_L g354 ( 
.A1(n_289),
.A2(n_227),
.B(n_272),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g379 ( 
.A1(n_354),
.A2(n_318),
.B1(n_295),
.B2(n_309),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_355),
.A2(n_356),
.B1(n_299),
.B2(n_312),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_308),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_347),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_315),
.A2(n_260),
.B(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_293),
.A2(n_287),
.B1(n_288),
.B2(n_290),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_279),
.B(n_311),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_279),
.B(n_316),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_412)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_387),
.C(n_399),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_344),
.A2(n_319),
.B(n_291),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_334),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_333),
.A2(n_303),
.B1(n_297),
.B2(n_276),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_374),
.A2(n_385),
.B1(n_324),
.B2(n_354),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_322),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_344),
.A2(n_283),
.B(n_306),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_380),
.Y(n_418)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_329),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_347),
.A2(n_285),
.B(n_294),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_384),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_333),
.A2(n_320),
.B1(n_292),
.B2(n_307),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_286),
.C(n_321),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_391),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_300),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_360),
.Y(n_405)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_394),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_330),
.A2(n_312),
.B1(n_364),
.B2(n_354),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_327),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_397),
.A2(n_398),
.B1(n_400),
.B2(n_394),
.Y(n_419)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_323),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_399),
.C(n_368),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_409),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_403),
.A2(n_370),
.B1(n_398),
.B2(n_367),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_405),
.B(n_371),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_375),
.B(n_325),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_411),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_361),
.C(n_334),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_382),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_342),
.C(n_358),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_425),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_400),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_422),
.Y(n_440)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_419),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_365),
.A2(n_354),
.B1(n_342),
.B2(n_355),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_421),
.B1(n_384),
.B2(n_390),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_372),
.A2(n_354),
.B1(n_331),
.B2(n_352),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_331),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_351),
.C(n_339),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_386),
.B(n_335),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_379),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_351),
.C(n_339),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_430),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_374),
.C(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_391),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_376),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_383),
.B1(n_377),
.B2(n_370),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_416),
.A2(n_383),
.B(n_377),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_435),
.A2(n_447),
.B(n_444),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_444),
.C(n_446),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_424),
.A2(n_336),
.B1(n_337),
.B2(n_343),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_438),
.A2(n_441),
.B1(n_326),
.B2(n_329),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_346),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_452),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_376),
.Y(n_443)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_445),
.A2(n_408),
.B1(n_420),
.B2(n_422),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_379),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_416),
.A2(n_379),
.B(n_381),
.Y(n_447)
);

NAND3xp33_ASAP7_75t_SL g468 ( 
.A(n_447),
.B(n_435),
.C(n_451),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_389),
.B(n_393),
.C(n_329),
.Y(n_451)
);

A2O1A1O1Ixp25_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_401),
.B(n_404),
.C(n_423),
.D(n_426),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_428),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_421),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_430),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_425),
.Y(n_455)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_456),
.B(n_457),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_409),
.B(n_326),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_407),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_460),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_407),
.C(n_413),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_459),
.B(n_472),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_405),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_464),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_412),
.Y(n_467)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_406),
.C(n_427),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_432),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_477),
.B1(n_445),
.B2(n_453),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_454),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_431),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_449),
.Y(n_489)
);

NAND4xp25_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_466),
.C(n_462),
.D(n_478),
.Y(n_495)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_483),
.Y(n_498)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_485),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_458),
.B(n_455),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_487),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_461),
.B(n_449),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_491),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_440),
.C(n_436),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_492),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_463),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_440),
.C(n_436),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_454),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_495),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_465),
.A2(n_434),
.B1(n_454),
.B2(n_467),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_494),
.A2(n_464),
.B1(n_479),
.B2(n_470),
.Y(n_497)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_497),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_496),
.A2(n_474),
.B(n_471),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_499),
.A2(n_510),
.B(n_497),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_460),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_503),
.Y(n_513)
);

INVx6_ASAP7_75t_L g502 ( 
.A(n_495),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_510),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_469),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_469),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_504),
.B(n_503),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_472),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_482),
.B(n_490),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_481),
.A2(n_484),
.B1(n_491),
.B2(n_483),
.Y(n_510)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_512),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_488),
.C(n_480),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_517),
.Y(n_523)
);

FAx1_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_493),
.CI(n_494),
.CON(n_515),
.SN(n_515)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_515),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_505),
.C(n_500),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_518),
.A2(n_519),
.B(n_521),
.Y(n_525)
);

AOI21xp33_ASAP7_75t_L g519 ( 
.A1(n_499),
.A2(n_500),
.B(n_508),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_507),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_521),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_504),
.C(n_514),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_513),
.C(n_518),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_525),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_516),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_528),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_513),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_529),
.B(n_531),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_532),
.A2(n_527),
.B(n_526),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_530),
.B(n_515),
.C(n_524),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_535),
.B(n_524),
.Y(n_536)
);

AOI21x1_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_533),
.B(n_515),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_529),
.Y(n_538)
);


endmodule