module fake_jpeg_5684_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

OR2x4_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_25),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_16),
.B1(n_27),
.B2(n_19),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_38),
.B1(n_28),
.B2(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_16),
.B1(n_17),
.B2(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_16),
.B1(n_28),
.B2(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_53),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_62),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_65),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_33),
.B(n_17),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_48),
.B(n_21),
.Y(n_83)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_51),
.B(n_53),
.C(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_74),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_58),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_31),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_80),
.C(n_73),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_44),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_68),
.B(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_26),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_61),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_84),
.C(n_41),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

AO221x1_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_107),
.B1(n_77),
.B2(n_99),
.C(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_78),
.B1(n_80),
.B2(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_109),
.C(n_110),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_48),
.C(n_65),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_61),
.C(n_62),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_117),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_29),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_22),
.B(n_20),
.C(n_24),
.D(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_90),
.B(n_87),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_107),
.B(n_102),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_24),
.C(n_20),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_91),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_115),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_88),
.B(n_29),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_128),
.B(n_22),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_127),
.Y(n_134)
);

INVxp33_ASAP7_75t_SL g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_46),
.B1(n_77),
.B2(n_35),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_3),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_141),
.B1(n_129),
.B2(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_142),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_122),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_140),
.C(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_20),
.B(n_54),
.C(n_49),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_54),
.C(n_49),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_49),
.B1(n_22),
.B2(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_4),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_139),
.C(n_5),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_150),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_22),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_124),
.B1(n_5),
.B2(n_6),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_160),
.B(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_150),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_146),
.B1(n_136),
.B2(n_137),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_156),
.B1(n_161),
.B2(n_6),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_R g159 ( 
.A(n_153),
.B(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_10),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_167),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_12),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_4),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_161),
.B(n_7),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_172),
.B(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_7),
.B(n_8),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_7),
.C(n_8),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);


endmodule