module fake_netlist_6_3454_n_5843 (n_992, n_1671, n_1, n_801, n_1613, n_1234, n_1458, n_1199, n_1674, n_741, n_1027, n_1351, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_212, n_700, n_50, n_1307, n_1038, n_578, n_1581, n_1003, n_365, n_168, n_1237, n_1061, n_1357, n_77, n_783, n_798, n_188, n_1575, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_677, n_805, n_1151, n_396, n_350, n_78, n_1380, n_442, n_480, n_142, n_1402, n_1009, n_62, n_1160, n_883, n_1238, n_1032, n_1247, n_1547, n_1553, n_893, n_1099, n_1264, n_1192, n_471, n_424, n_1555, n_1415, n_1370, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_1285, n_1371, n_200, n_447, n_1172, n_852, n_71, n_229, n_1590, n_1532, n_1393, n_1517, n_1078, n_250, n_544, n_1140, n_1444, n_1670, n_1603, n_1579, n_35, n_1263, n_836, n_375, n_522, n_1261, n_945, n_1649, n_1511, n_1143, n_1422, n_1232, n_1572, n_616, n_658, n_1119, n_428, n_1433, n_1620, n_1541, n_1300, n_641, n_822, n_693, n_1313, n_1056, n_758, n_516, n_1455, n_1163, n_1180, n_943, n_1550, n_491, n_1591, n_42, n_772, n_1344, n_666, n_371, n_940, n_770, n_567, n_405, n_213, n_538, n_1106, n_886, n_1471, n_343, n_953, n_1094, n_1345, n_494, n_539, n_493, n_155, n_45, n_454, n_1421, n_638, n_1404, n_1211, n_381, n_887, n_1660, n_112, n_1280, n_713, n_1400, n_126, n_1467, n_58, n_976, n_224, n_48, n_1445, n_1526, n_1560, n_734, n_1088, n_196, n_1231, n_917, n_574, n_9, n_907, n_6, n_1446, n_14, n_659, n_407, n_913, n_1658, n_808, n_867, n_1230, n_473, n_1193, n_1054, n_559, n_1333, n_44, n_1648, n_163, n_1644, n_1558, n_281, n_551, n_699, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_1641, n_577, n_166, n_619, n_1367, n_1336, n_521, n_572, n_395, n_813, n_1481, n_323, n_606, n_1441, n_818, n_1123, n_1309, n_92, n_513, n_645, n_1381, n_331, n_916, n_483, n_102, n_608, n_261, n_630, n_32, n_541, n_512, n_121, n_433, n_792, n_476, n_2, n_1328, n_219, n_264, n_263, n_1162, n_860, n_1530, n_788, n_939, n_1543, n_821, n_938, n_1302, n_1068, n_1599, n_329, n_982, n_549, n_1075, n_408, n_932, n_61, n_237, n_243, n_979, n_905, n_1680, n_117, n_175, n_322, n_993, n_689, n_354, n_1330, n_1413, n_1605, n_134, n_1278, n_547, n_558, n_1064, n_1396, n_634, n_136, n_966, n_764, n_1663, n_692, n_733, n_1233, n_1289, n_487, n_241, n_30, n_1107, n_1014, n_1290, n_882, n_1354, n_586, n_423, n_318, n_1111, n_715, n_1251, n_1265, n_88, n_530, n_1563, n_277, n_618, n_1297, n_1662, n_1312, n_199, n_1167, n_1359, n_674, n_871, n_922, n_268, n_1335, n_210, n_1069, n_5, n_1664, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_1175, n_328, n_1386, n_429, n_1012, n_195, n_780, n_675, n_903, n_1540, n_1504, n_286, n_254, n_1655, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_1654, n_816, n_1157, n_1462, n_1188, n_877, n_604, n_825, n_728, n_1063, n_1588, n_26, n_55, n_267, n_1124, n_1624, n_515, n_598, n_696, n_1515, n_961, n_437, n_1082, n_1317, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_950, n_388, n_190, n_484, n_170, n_891, n_1412, n_949, n_1630, n_678, n_283, n_91, n_507, n_968, n_909, n_1369, n_881, n_1008, n_760, n_1546, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_1296, n_304, n_694, n_1294, n_1420, n_125, n_1634, n_297, n_595, n_627, n_524, n_1465, n_342, n_1044, n_1391, n_449, n_131, n_1523, n_1208, n_1164, n_1295, n_1627, n_1072, n_1527, n_1495, n_1438, n_495, n_815, n_1100, n_585, n_1487, n_840, n_874, n_1128, n_382, n_673, n_1071, n_1067, n_1565, n_1493, n_898, n_255, n_284, n_865, n_925, n_1101, n_15, n_1026, n_38, n_289, n_1364, n_615, n_1249, n_59, n_1293, n_1127, n_1512, n_1451, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_685, n_353, n_605, n_1514, n_826, n_1646, n_872, n_1139, n_86, n_104, n_718, n_1018, n_1521, n_1366, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_1308, n_1376, n_1513, n_413, n_791, n_510, n_837, n_79, n_1488, n_948, n_704, n_977, n_1005, n_536, n_622, n_147, n_1469, n_581, n_765, n_432, n_987, n_1492, n_1340, n_631, n_720, n_153, n_842, n_1432, n_156, n_145, n_843, n_656, n_989, n_1277, n_797, n_1473, n_1246, n_899, n_189, n_738, n_1304, n_1035, n_294, n_499, n_1426, n_705, n_11, n_1004, n_1176, n_1529, n_1022, n_614, n_529, n_425, n_684, n_1431, n_1615, n_1474, n_1571, n_1577, n_1181, n_37, n_486, n_947, n_1117, n_1087, n_1448, n_648, n_657, n_1049, n_1666, n_1505, n_803, n_290, n_118, n_926, n_927, n_919, n_478, n_929, n_107, n_1228, n_417, n_446, n_89, n_1568, n_1490, n_777, n_1299, n_272, n_526, n_1183, n_1436, n_1384, n_69, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_1665, n_18, n_154, n_1383, n_1178, n_98, n_1424, n_1073, n_1000, n_796, n_252, n_1195, n_1626, n_1507, n_184, n_552, n_1358, n_1388, n_216, n_912, n_1519, n_745, n_1284, n_1604, n_1142, n_716, n_1475, n_623, n_1048, n_1201, n_1398, n_884, n_1395, n_731, n_1502, n_1659, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_1368, n_66, n_1418, n_958, n_292, n_1250, n_100, n_1137, n_880, n_889, n_150, n_1478, n_589, n_1310, n_819, n_1363, n_1334, n_767, n_1314, n_600, n_964, n_831, n_477, n_954, n_864, n_1110, n_1410, n_399, n_1440, n_124, n_1382, n_1534, n_1564, n_211, n_1483, n_1372, n_231, n_40, n_1457, n_505, n_319, n_1339, n_537, n_1427, n_311, n_1466, n_10, n_403, n_1080, n_723, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1220, n_556, n_162, n_1602, n_1136, n_128, n_1125, n_970, n_642, n_995, n_276, n_1159, n_1092, n_441, n_221, n_1060, n_444, n_146, n_1252, n_1223, n_303, n_511, n_193, n_1286, n_1053, n_416, n_520, n_418, n_1093, n_113, n_1533, n_1597, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_1618, n_217, n_518, n_1531, n_1185, n_453, n_215, n_914, n_759, n_426, n_317, n_1653, n_1679, n_1625, n_90, n_54, n_1453, n_488, n_497, n_773, n_920, n_99, n_1374, n_1315, n_1647, n_13, n_1224, n_1614, n_1459, n_1135, n_1169, n_1179, n_401, n_324, n_1617, n_335, n_1470, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_1091, n_1580, n_1425, n_36, n_1267, n_1281, n_983, n_427, n_1520, n_496, n_906, n_1390, n_688, n_1077, n_1419, n_351, n_259, n_177, n_1636, n_1437, n_1645, n_385, n_1439, n_1323, n_858, n_1331, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_379, n_778, n_1668, n_1134, n_410, n_1129, n_554, n_602, n_1594, n_664, n_171, n_169, n_1429, n_1610, n_435, n_793, n_326, n_587, n_1593, n_580, n_762, n_1030, n_1202, n_465, n_1635, n_1079, n_341, n_828, n_607, n_316, n_419, n_28, n_1551, n_1103, n_144, n_1203, n_820, n_951, n_106, n_725, n_952, n_999, n_358, n_1254, n_160, n_186, n_0, n_368, n_575, n_994, n_1508, n_732, n_974, n_392, n_724, n_1020, n_1042, n_628, n_1273, n_1434, n_1573, n_557, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_1661, n_1275, n_485, n_1549, n_67, n_443, n_1510, n_892, n_768, n_421, n_1468, n_238, n_1095, n_1595, n_202, n_597, n_280, n_1270, n_1187, n_610, n_1403, n_1669, n_1024, n_198, n_179, n_248, n_517, n_1667, n_667, n_1206, n_621, n_1037, n_1397, n_1279, n_1115, n_750, n_901, n_1499, n_468, n_923, n_504, n_1409, n_1639, n_1623, n_183, n_1015, n_1503, n_466, n_1057, n_603, n_991, n_1657, n_235, n_1126, n_340, n_710, n_1108, n_1182, n_1298, n_39, n_73, n_1611, n_785, n_746, n_609, n_1601, n_101, n_167, n_1356, n_1589, n_127, n_1497, n_1168, n_1216, n_133, n_1320, n_96, n_1430, n_1316, n_1287, n_1452, n_1622, n_1586, n_302, n_380, n_1535, n_137, n_1596, n_20, n_1190, n_397, n_122, n_34, n_1262, n_218, n_1213, n_70, n_1350, n_1673, n_172, n_1443, n_1272, n_239, n_97, n_782, n_1539, n_490, n_220, n_809, n_1043, n_1608, n_986, n_80, n_1472, n_1081, n_402, n_352, n_800, n_1084, n_1171, n_460, n_1361, n_1491, n_662, n_374, n_1152, n_450, n_921, n_1346, n_711, n_1642, n_579, n_1352, n_937, n_370, n_650, n_1046, n_1145, n_330, n_1121, n_1102, n_972, n_1405, n_258, n_1406, n_456, n_1332, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_1569, n_936, n_1288, n_1186, n_1062, n_885, n_896, n_83, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_105, n_227, n_204, n_482, n_934, n_1637, n_1407, n_420, n_1341, n_394, n_1456, n_1489, n_164, n_23, n_942, n_1524, n_543, n_1496, n_1271, n_1545, n_1355, n_1225, n_1544, n_1485, n_325, n_1640, n_804, n_464, n_533, n_806, n_879, n_959, n_584, n_244, n_1343, n_1522, n_76, n_548, n_94, n_282, n_1676, n_833, n_1567, n_523, n_1319, n_707, n_345, n_799, n_1548, n_1155, n_139, n_41, n_273, n_1633, n_787, n_1416, n_1528, n_1146, n_159, n_1086, n_1066, n_157, n_1282, n_550, n_275, n_652, n_560, n_1484, n_1241, n_1321, n_1672, n_569, n_737, n_1318, n_1235, n_1229, n_306, n_1292, n_1373, n_21, n_346, n_3, n_1029, n_1447, n_790, n_138, n_1498, n_1210, n_49, n_299, n_1248, n_1556, n_902, n_333, n_1047, n_1385, n_431, n_24, n_459, n_1269, n_502, n_672, n_1257, n_285, n_1375, n_85, n_655, n_706, n_1045, n_1650, n_786, n_1236, n_1559, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1325, n_1002, n_545, n_489, n_251, n_1019, n_636, n_729, n_110, n_151, n_876, n_774, n_1337, n_660, n_438, n_1477, n_1360, n_1200, n_479, n_1607, n_1353, n_1454, n_869, n_1154, n_1113, n_1600, n_646, n_528, n_391, n_1098, n_1329, n_817, n_262, n_187, n_897, n_846, n_841, n_1476, n_1001, n_508, n_1050, n_1411, n_1463, n_1177, n_332, n_1150, n_1562, n_398, n_1191, n_566, n_1023, n_1076, n_1118, n_194, n_57, n_1007, n_1378, n_855, n_1592, n_1631, n_52, n_591, n_1377, n_256, n_853, n_440, n_695, n_1542, n_875, n_209, n_367, n_680, n_1678, n_661, n_278, n_1256, n_671, n_7, n_933, n_740, n_703, n_978, n_384, n_1291, n_1217, n_751, n_749, n_310, n_1628, n_1324, n_1399, n_1435, n_969, n_988, n_1065, n_84, n_1401, n_1255, n_568, n_1516, n_143, n_1536, n_180, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_1327, n_1326, n_739, n_400, n_955, n_337, n_1379, n_214, n_246, n_1338, n_1097, n_935, n_781, n_789, n_1554, n_1130, n_181, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_1583, n_555, n_389, n_814, n_1643, n_669, n_176, n_114, n_300, n_222, n_747, n_74, n_1389, n_1105, n_721, n_1461, n_742, n_535, n_691, n_372, n_111, n_314, n_1408, n_378, n_1196, n_377, n_1598, n_863, n_601, n_338, n_1283, n_918, n_748, n_506, n_1114, n_56, n_763, n_1147, n_360, n_1506, n_119, n_1652, n_957, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1303, n_1205, n_1258, n_1392, n_174, n_1173, n_525, n_1677, n_1116, n_611, n_1570, n_1219, n_8, n_1174, n_1016, n_1347, n_795, n_1501, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_1083, n_109, n_445, n_1561, n_930, n_888, n_1112, n_234, n_910, n_1656, n_1460, n_911, n_82, n_1464, n_27, n_236, n_653, n_1414, n_752, n_908, n_944, n_576, n_1028, n_472, n_270, n_414, n_563, n_1011, n_1566, n_1215, n_25, n_93, n_839, n_708, n_668, n_626, n_990, n_1500, n_779, n_1537, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_1509, n_103, n_1109, n_185, n_712, n_348, n_1276, n_376, n_390, n_1148, n_31, n_334, n_1161, n_1085, n_232, n_46, n_1239, n_771, n_1584, n_470, n_475, n_924, n_298, n_1582, n_492, n_1149, n_265, n_1184, n_228, n_719, n_1525, n_455, n_1585, n_363, n_1090, n_592, n_1518, n_829, n_1156, n_1362, n_393, n_984, n_503, n_1450, n_1638, n_132, n_868, n_570, n_859, n_406, n_735, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_1482, n_981, n_714, n_1349, n_291, n_1144, n_357, n_985, n_481, n_997, n_1301, n_802, n_561, n_33, n_980, n_1306, n_1651, n_1198, n_1609, n_436, n_116, n_409, n_1244, n_1574, n_240, n_756, n_1619, n_1606, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_1552, n_583, n_249, n_201, n_1039, n_1442, n_1034, n_1480, n_1158, n_754, n_941, n_975, n_1031, n_115, n_1305, n_553, n_43, n_849, n_753, n_467, n_269, n_359, n_973, n_1479, n_1055, n_1675, n_582, n_861, n_857, n_967, n_571, n_271, n_404, n_158, n_206, n_679, n_633, n_1170, n_665, n_1629, n_588, n_225, n_1260, n_308, n_309, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_812, n_1131, n_534, n_1578, n_1006, n_373, n_87, n_1632, n_257, n_1557, n_730, n_1311, n_1494, n_670, n_203, n_207, n_1089, n_1587, n_1365, n_1417, n_205, n_1242, n_681, n_1226, n_1274, n_1486, n_412, n_640, n_1322, n_81, n_965, n_1428, n_1616, n_1576, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_135, n_165, n_540, n_1423, n_457, n_364, n_629, n_1621, n_900, n_1449, n_531, n_827, n_60, n_361, n_1025, n_336, n_12, n_1013, n_1259, n_192, n_1538, n_51, n_649, n_1612, n_1240, n_5843);

input n_992;
input n_1671;
input n_1;
input n_801;
input n_1613;
input n_1234;
input n_1458;
input n_1199;
input n_1674;
input n_741;
input n_1027;
input n_1351;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_212;
input n_700;
input n_50;
input n_1307;
input n_1038;
input n_578;
input n_1581;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_1357;
input n_77;
input n_783;
input n_798;
input n_188;
input n_1575;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_677;
input n_805;
input n_1151;
input n_396;
input n_350;
input n_78;
input n_1380;
input n_442;
input n_480;
input n_142;
input n_1402;
input n_1009;
input n_62;
input n_1160;
input n_883;
input n_1238;
input n_1032;
input n_1247;
input n_1547;
input n_1553;
input n_893;
input n_1099;
input n_1264;
input n_1192;
input n_471;
input n_424;
input n_1555;
input n_1415;
input n_1370;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_200;
input n_447;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1590;
input n_1532;
input n_1393;
input n_1517;
input n_1078;
input n_250;
input n_544;
input n_1140;
input n_1444;
input n_1670;
input n_1603;
input n_1579;
input n_35;
input n_1263;
input n_836;
input n_375;
input n_522;
input n_1261;
input n_945;
input n_1649;
input n_1511;
input n_1143;
input n_1422;
input n_1232;
input n_1572;
input n_616;
input n_658;
input n_1119;
input n_428;
input n_1433;
input n_1620;
input n_1541;
input n_1300;
input n_641;
input n_822;
input n_693;
input n_1313;
input n_1056;
input n_758;
input n_516;
input n_1455;
input n_1163;
input n_1180;
input n_943;
input n_1550;
input n_491;
input n_1591;
input n_42;
input n_772;
input n_1344;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_405;
input n_213;
input n_538;
input n_1106;
input n_886;
input n_1471;
input n_343;
input n_953;
input n_1094;
input n_1345;
input n_494;
input n_539;
input n_493;
input n_155;
input n_45;
input n_454;
input n_1421;
input n_638;
input n_1404;
input n_1211;
input n_381;
input n_887;
input n_1660;
input n_112;
input n_1280;
input n_713;
input n_1400;
input n_126;
input n_1467;
input n_58;
input n_976;
input n_224;
input n_48;
input n_1445;
input n_1526;
input n_1560;
input n_734;
input n_1088;
input n_196;
input n_1231;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_1446;
input n_14;
input n_659;
input n_407;
input n_913;
input n_1658;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1054;
input n_559;
input n_1333;
input n_44;
input n_1648;
input n_163;
input n_1644;
input n_1558;
input n_281;
input n_551;
input n_699;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_1641;
input n_577;
input n_166;
input n_619;
input n_1367;
input n_1336;
input n_521;
input n_572;
input n_395;
input n_813;
input n_1481;
input n_323;
input n_606;
input n_1441;
input n_818;
input n_1123;
input n_1309;
input n_92;
input n_513;
input n_645;
input n_1381;
input n_331;
input n_916;
input n_483;
input n_102;
input n_608;
input n_261;
input n_630;
input n_32;
input n_541;
input n_512;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_1328;
input n_219;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_1530;
input n_788;
input n_939;
input n_1543;
input n_821;
input n_938;
input n_1302;
input n_1068;
input n_1599;
input n_329;
input n_982;
input n_549;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_243;
input n_979;
input n_905;
input n_1680;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_354;
input n_1330;
input n_1413;
input n_1605;
input n_134;
input n_1278;
input n_547;
input n_558;
input n_1064;
input n_1396;
input n_634;
input n_136;
input n_966;
input n_764;
input n_1663;
input n_692;
input n_733;
input n_1233;
input n_1289;
input n_487;
input n_241;
input n_30;
input n_1107;
input n_1014;
input n_1290;
input n_882;
input n_1354;
input n_586;
input n_423;
input n_318;
input n_1111;
input n_715;
input n_1251;
input n_1265;
input n_88;
input n_530;
input n_1563;
input n_277;
input n_618;
input n_1297;
input n_1662;
input n_1312;
input n_199;
input n_1167;
input n_1359;
input n_674;
input n_871;
input n_922;
input n_268;
input n_1335;
input n_210;
input n_1069;
input n_5;
input n_1664;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_1175;
input n_328;
input n_1386;
input n_429;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_1540;
input n_1504;
input n_286;
input n_254;
input n_1655;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_1654;
input n_816;
input n_1157;
input n_1462;
input n_1188;
input n_877;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_1588;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_1624;
input n_515;
input n_598;
input n_696;
input n_1515;
input n_961;
input n_437;
input n_1082;
input n_1317;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_950;
input n_388;
input n_190;
input n_484;
input n_170;
input n_891;
input n_1412;
input n_949;
input n_1630;
input n_678;
input n_283;
input n_91;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_881;
input n_1008;
input n_760;
input n_1546;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_1296;
input n_304;
input n_694;
input n_1294;
input n_1420;
input n_125;
input n_1634;
input n_297;
input n_595;
input n_627;
input n_524;
input n_1465;
input n_342;
input n_1044;
input n_1391;
input n_449;
input n_131;
input n_1523;
input n_1208;
input n_1164;
input n_1295;
input n_1627;
input n_1072;
input n_1527;
input n_1495;
input n_1438;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_1487;
input n_840;
input n_874;
input n_1128;
input n_382;
input n_673;
input n_1071;
input n_1067;
input n_1565;
input n_1493;
input n_898;
input n_255;
input n_284;
input n_865;
input n_925;
input n_1101;
input n_15;
input n_1026;
input n_38;
input n_289;
input n_1364;
input n_615;
input n_1249;
input n_59;
input n_1293;
input n_1127;
input n_1512;
input n_1451;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_605;
input n_1514;
input n_826;
input n_1646;
input n_872;
input n_1139;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_1521;
input n_1366;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_1376;
input n_1513;
input n_413;
input n_791;
input n_510;
input n_837;
input n_79;
input n_1488;
input n_948;
input n_704;
input n_977;
input n_1005;
input n_536;
input n_622;
input n_147;
input n_1469;
input n_581;
input n_765;
input n_432;
input n_987;
input n_1492;
input n_1340;
input n_631;
input n_720;
input n_153;
input n_842;
input n_1432;
input n_156;
input n_145;
input n_843;
input n_656;
input n_989;
input n_1277;
input n_797;
input n_1473;
input n_1246;
input n_899;
input n_189;
input n_738;
input n_1304;
input n_1035;
input n_294;
input n_499;
input n_1426;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_1529;
input n_1022;
input n_614;
input n_529;
input n_425;
input n_684;
input n_1431;
input n_1615;
input n_1474;
input n_1571;
input n_1577;
input n_1181;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_1448;
input n_648;
input n_657;
input n_1049;
input n_1666;
input n_1505;
input n_803;
input n_290;
input n_118;
input n_926;
input n_927;
input n_919;
input n_478;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_1568;
input n_1490;
input n_777;
input n_1299;
input n_272;
input n_526;
input n_1183;
input n_1436;
input n_1384;
input n_69;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_1665;
input n_18;
input n_154;
input n_1383;
input n_1178;
input n_98;
input n_1424;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_1626;
input n_1507;
input n_184;
input n_552;
input n_1358;
input n_1388;
input n_216;
input n_912;
input n_1519;
input n_745;
input n_1284;
input n_1604;
input n_1142;
input n_716;
input n_1475;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1395;
input n_731;
input n_1502;
input n_1659;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_1368;
input n_66;
input n_1418;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_880;
input n_889;
input n_150;
input n_1478;
input n_589;
input n_1310;
input n_819;
input n_1363;
input n_1334;
input n_767;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_1410;
input n_399;
input n_1440;
input n_124;
input n_1382;
input n_1534;
input n_1564;
input n_211;
input n_1483;
input n_1372;
input n_231;
input n_40;
input n_1457;
input n_505;
input n_319;
input n_1339;
input n_537;
input n_1427;
input n_311;
input n_1466;
input n_10;
input n_403;
input n_1080;
input n_723;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1220;
input n_556;
input n_162;
input n_1602;
input n_1136;
input n_128;
input n_1125;
input n_970;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_441;
input n_221;
input n_1060;
input n_444;
input n_146;
input n_1252;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1286;
input n_1053;
input n_416;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_1533;
input n_1597;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_1618;
input n_217;
input n_518;
input n_1531;
input n_1185;
input n_453;
input n_215;
input n_914;
input n_759;
input n_426;
input n_317;
input n_1653;
input n_1679;
input n_1625;
input n_90;
input n_54;
input n_1453;
input n_488;
input n_497;
input n_773;
input n_920;
input n_99;
input n_1374;
input n_1315;
input n_1647;
input n_13;
input n_1224;
input n_1614;
input n_1459;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_1617;
input n_335;
input n_1470;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_1091;
input n_1580;
input n_1425;
input n_36;
input n_1267;
input n_1281;
input n_983;
input n_427;
input n_1520;
input n_496;
input n_906;
input n_1390;
input n_688;
input n_1077;
input n_1419;
input n_351;
input n_259;
input n_177;
input n_1636;
input n_1437;
input n_1645;
input n_385;
input n_1439;
input n_1323;
input n_858;
input n_1331;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_379;
input n_778;
input n_1668;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_1594;
input n_664;
input n_171;
input n_169;
input n_1429;
input n_1610;
input n_435;
input n_793;
input n_326;
input n_587;
input n_1593;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_465;
input n_1635;
input n_1079;
input n_341;
input n_828;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1551;
input n_1103;
input n_144;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_1508;
input n_732;
input n_974;
input n_392;
input n_724;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_1434;
input n_1573;
input n_557;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_1661;
input n_1275;
input n_485;
input n_1549;
input n_67;
input n_443;
input n_1510;
input n_892;
input n_768;
input n_421;
input n_1468;
input n_238;
input n_1095;
input n_1595;
input n_202;
input n_597;
input n_280;
input n_1270;
input n_1187;
input n_610;
input n_1403;
input n_1669;
input n_1024;
input n_198;
input n_179;
input n_248;
input n_517;
input n_1667;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1397;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_1499;
input n_468;
input n_923;
input n_504;
input n_1409;
input n_1639;
input n_1623;
input n_183;
input n_1015;
input n_1503;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_1657;
input n_235;
input n_1126;
input n_340;
input n_710;
input n_1108;
input n_1182;
input n_1298;
input n_39;
input n_73;
input n_1611;
input n_785;
input n_746;
input n_609;
input n_1601;
input n_101;
input n_167;
input n_1356;
input n_1589;
input n_127;
input n_1497;
input n_1168;
input n_1216;
input n_133;
input n_1320;
input n_96;
input n_1430;
input n_1316;
input n_1287;
input n_1452;
input n_1622;
input n_1586;
input n_302;
input n_380;
input n_1535;
input n_137;
input n_1596;
input n_20;
input n_1190;
input n_397;
input n_122;
input n_34;
input n_1262;
input n_218;
input n_1213;
input n_70;
input n_1350;
input n_1673;
input n_172;
input n_1443;
input n_1272;
input n_239;
input n_97;
input n_782;
input n_1539;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_1608;
input n_986;
input n_80;
input n_1472;
input n_1081;
input n_402;
input n_352;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_1361;
input n_1491;
input n_662;
input n_374;
input n_1152;
input n_450;
input n_921;
input n_1346;
input n_711;
input n_1642;
input n_579;
input n_1352;
input n_937;
input n_370;
input n_650;
input n_1046;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_972;
input n_1405;
input n_258;
input n_1406;
input n_456;
input n_1332;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_1569;
input n_936;
input n_1288;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_105;
input n_227;
input n_204;
input n_482;
input n_934;
input n_1637;
input n_1407;
input n_420;
input n_1341;
input n_394;
input n_1456;
input n_1489;
input n_164;
input n_23;
input n_942;
input n_1524;
input n_543;
input n_1496;
input n_1271;
input n_1545;
input n_1355;
input n_1225;
input n_1544;
input n_1485;
input n_325;
input n_1640;
input n_804;
input n_464;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_244;
input n_1343;
input n_1522;
input n_76;
input n_548;
input n_94;
input n_282;
input n_1676;
input n_833;
input n_1567;
input n_523;
input n_1319;
input n_707;
input n_345;
input n_799;
input n_1548;
input n_1155;
input n_139;
input n_41;
input n_273;
input n_1633;
input n_787;
input n_1416;
input n_1528;
input n_1146;
input n_159;
input n_1086;
input n_1066;
input n_157;
input n_1282;
input n_550;
input n_275;
input n_652;
input n_560;
input n_1484;
input n_1241;
input n_1321;
input n_1672;
input n_569;
input n_737;
input n_1318;
input n_1235;
input n_1229;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_1447;
input n_790;
input n_138;
input n_1498;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_1556;
input n_902;
input n_333;
input n_1047;
input n_1385;
input n_431;
input n_24;
input n_459;
input n_1269;
input n_502;
input n_672;
input n_1257;
input n_285;
input n_1375;
input n_85;
input n_655;
input n_706;
input n_1045;
input n_1650;
input n_786;
input n_1236;
input n_1559;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1325;
input n_1002;
input n_545;
input n_489;
input n_251;
input n_1019;
input n_636;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_1337;
input n_660;
input n_438;
input n_1477;
input n_1360;
input n_1200;
input n_479;
input n_1607;
input n_1353;
input n_1454;
input n_869;
input n_1154;
input n_1113;
input n_1600;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_1329;
input n_817;
input n_262;
input n_187;
input n_897;
input n_846;
input n_841;
input n_1476;
input n_1001;
input n_508;
input n_1050;
input n_1411;
input n_1463;
input n_1177;
input n_332;
input n_1150;
input n_1562;
input n_398;
input n_1191;
input n_566;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_1378;
input n_855;
input n_1592;
input n_1631;
input n_52;
input n_591;
input n_1377;
input n_256;
input n_853;
input n_440;
input n_695;
input n_1542;
input n_875;
input n_209;
input n_367;
input n_680;
input n_1678;
input n_661;
input n_278;
input n_1256;
input n_671;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1291;
input n_1217;
input n_751;
input n_749;
input n_310;
input n_1628;
input n_1324;
input n_1399;
input n_1435;
input n_969;
input n_988;
input n_1065;
input n_84;
input n_1401;
input n_1255;
input n_568;
input n_1516;
input n_143;
input n_1536;
input n_180;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_1379;
input n_214;
input n_246;
input n_1338;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1554;
input n_1130;
input n_181;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_1583;
input n_555;
input n_389;
input n_814;
input n_1643;
input n_669;
input n_176;
input n_114;
input n_300;
input n_222;
input n_747;
input n_74;
input n_1389;
input n_1105;
input n_721;
input n_1461;
input n_742;
input n_535;
input n_691;
input n_372;
input n_111;
input n_314;
input n_1408;
input n_378;
input n_1196;
input n_377;
input n_1598;
input n_863;
input n_601;
input n_338;
input n_1283;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1147;
input n_360;
input n_1506;
input n_119;
input n_1652;
input n_957;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1303;
input n_1205;
input n_1258;
input n_1392;
input n_174;
input n_1173;
input n_525;
input n_1677;
input n_1116;
input n_611;
input n_1570;
input n_1219;
input n_8;
input n_1174;
input n_1016;
input n_1347;
input n_795;
input n_1501;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_1083;
input n_109;
input n_445;
input n_1561;
input n_930;
input n_888;
input n_1112;
input n_234;
input n_910;
input n_1656;
input n_1460;
input n_911;
input n_82;
input n_1464;
input n_27;
input n_236;
input n_653;
input n_1414;
input n_752;
input n_908;
input n_944;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_414;
input n_563;
input n_1011;
input n_1566;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_668;
input n_626;
input n_990;
input n_1500;
input n_779;
input n_1537;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_1509;
input n_103;
input n_1109;
input n_185;
input n_712;
input n_348;
input n_1276;
input n_376;
input n_390;
input n_1148;
input n_31;
input n_334;
input n_1161;
input n_1085;
input n_232;
input n_46;
input n_1239;
input n_771;
input n_1584;
input n_470;
input n_475;
input n_924;
input n_298;
input n_1582;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_1525;
input n_455;
input n_1585;
input n_363;
input n_1090;
input n_592;
input n_1518;
input n_829;
input n_1156;
input n_1362;
input n_393;
input n_984;
input n_503;
input n_1450;
input n_1638;
input n_132;
input n_868;
input n_570;
input n_859;
input n_406;
input n_735;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_1482;
input n_981;
input n_714;
input n_1349;
input n_291;
input n_1144;
input n_357;
input n_985;
input n_481;
input n_997;
input n_1301;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1306;
input n_1651;
input n_1198;
input n_1609;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_1574;
input n_240;
input n_756;
input n_1619;
input n_1606;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_1552;
input n_583;
input n_249;
input n_201;
input n_1039;
input n_1442;
input n_1034;
input n_1480;
input n_1158;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_1305;
input n_553;
input n_43;
input n_849;
input n_753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1479;
input n_1055;
input n_1675;
input n_582;
input n_861;
input n_857;
input n_967;
input n_571;
input n_271;
input n_404;
input n_158;
input n_206;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_1629;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_812;
input n_1131;
input n_534;
input n_1578;
input n_1006;
input n_373;
input n_87;
input n_1632;
input n_257;
input n_1557;
input n_730;
input n_1311;
input n_1494;
input n_670;
input n_203;
input n_207;
input n_1089;
input n_1587;
input n_1365;
input n_1417;
input n_205;
input n_1242;
input n_681;
input n_1226;
input n_1274;
input n_1486;
input n_412;
input n_640;
input n_1322;
input n_81;
input n_965;
input n_1428;
input n_1616;
input n_1576;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_135;
input n_165;
input n_540;
input n_1423;
input n_457;
input n_364;
input n_629;
input n_1621;
input n_900;
input n_1449;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_336;
input n_12;
input n_1013;
input n_1259;
input n_192;
input n_1538;
input n_51;
input n_649;
input n_1612;
input n_1240;

output n_5843;

wire n_5643;
wire n_2542;
wire n_2817;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_5315;
wire n_5254;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_3089;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_4829;
wire n_5393;
wire n_3222;
wire n_4699;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_2179;
wire n_5055;
wire n_3376;
wire n_4868;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_3564;
wire n_1844;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_5838;
wire n_5725;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_5598;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_5819;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_4814;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_4262;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_5638;
wire n_4110;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_5680;
wire n_4102;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_5504;
wire n_5522;
wire n_5828;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_5063;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_2641;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_5667;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_5281;
wire n_2092;
wire n_1750;
wire n_2514;
wire n_5314;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_5795;
wire n_4473;
wire n_5552;
wire n_5226;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_4394;
wire n_2279;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_3696;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_3614;
wire n_5183;
wire n_2145;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_5787;
wire n_3179;
wire n_3400;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_4345;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_5636;
wire n_2239;
wire n_4310;
wire n_5212;
wire n_2689;
wire n_5286;
wire n_2191;
wire n_4528;
wire n_5811;
wire n_4914;
wire n_4939;
wire n_3418;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_3631;
wire n_5599;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_5035;
wire n_3390;
wire n_3656;
wire n_3025;
wire n_2137;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_3006;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_5394;
wire n_4592;
wire n_2199;
wire n_2661;
wire n_5359;
wire n_1955;
wire n_1791;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_5741;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_3591;
wire n_2788;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_5176;
wire n_4428;
wire n_3323;
wire n_2274;
wire n_5761;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_2822;
wire n_4180;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_3299;
wire n_5688;
wire n_5740;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_5534;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_5023;
wire n_2656;
wire n_4952;
wire n_2375;
wire n_1934;
wire n_5660;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_4761;
wire n_2884;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_3797;
wire n_2024;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_4230;
wire n_2637;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_4189;
wire n_3817;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_5618;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_4380;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_3594;
wire n_5689;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_3210;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_5731;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_4601;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_5754;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_2798;
wire n_2852;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_3375;
wire n_3899;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_4512;
wire n_4081;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_5577;
wire n_5124;
wire n_3951;
wire n_3569;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_3027;
wire n_4083;
wire n_1810;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_5779;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_4027;
wire n_3154;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_4095;
wire n_2881;
wire n_1702;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_1944;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_3176;
wire n_5541;
wire n_5568;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_3697;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_5696;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_3936;
wire n_2723;
wire n_5485;
wire n_5823;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_4062;
wire n_3902;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_3101;
wire n_1981;
wire n_4233;
wire n_3374;
wire n_2640;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_3017;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_3795;
wire n_3852;
wire n_5289;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1862;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_5303;
wire n_3266;
wire n_3574;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_4504;
wire n_3844;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_4819;
wire n_5248;
wire n_1708;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_3946;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_3275;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_5788;
wire n_1902;
wire n_1842;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_3750;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_3532;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_5762;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_5519;
wire n_4047;
wire n_5753;
wire n_3413;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5808;
wire n_5436;
wire n_5139;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5822;
wire n_5195;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_4277;
wire n_4526;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_5792;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_3725;
wire n_3933;
wire n_5554;
wire n_2311;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_4066;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_4340;
wire n_5790;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_5757;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_1987;
wire n_2271;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_5484;
wire n_2954;
wire n_2728;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_3159;
wire n_4701;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_1913;
wire n_4934;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_2604;
wire n_2407;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_4114;
wire n_2948;
wire n_2119;
wire n_1992;
wire n_5686;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_3654;
wire n_2848;
wire n_1849;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_3324;
wire n_2338;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_2144;
wire n_4487;
wire n_4866;
wire n_4889;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_5773;
wire n_5482;
wire n_3393;
wire n_3451;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2892;
wire n_2132;
wire n_4120;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_5676;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1951;
wire n_4362;
wire n_3311;
wire n_3913;
wire n_5121;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_4404;
wire n_5589;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_2724;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_5807;
wire n_4448;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_2315;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_5273;
wire n_4844;
wire n_4438;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_2803;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_5706;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_5621;
wire n_5608;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_3250;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_3414;
wire n_4870;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_2598;
wire n_1916;
wire n_1683;
wire n_4304;
wire n_4558;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_4016;
wire n_5508;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_3730;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_5050;
wire n_2740;
wire n_4808;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_4192;
wire n_4109;
wire n_4824;
wire n_2808;
wire n_2037;
wire n_4567;
wire n_5150;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5585;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_5348;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_2970;
wire n_2167;
wire n_2342;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_2258;
wire n_5503;
wire n_2390;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_2734;
wire n_1782;
wire n_5600;
wire n_5755;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_3381;
wire n_3208;
wire n_2195;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_5749;
wire n_1925;
wire n_4407;
wire n_3517;
wire n_4045;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_4143;
wire n_4170;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_2588;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_5170;
wire n_2827;
wire n_3515;
wire n_2951;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1879;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_3629;
wire n_5400;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_4783;
wire n_4910;
wire n_3083;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_5623;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_5693;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_2463;
wire n_3363;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_5647;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_5803;
wire n_2112;
wire n_2430;
wire n_5285;
wire n_2721;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_4521;
wire n_3204;
wire n_5715;
wire n_4920;
wire n_5395;
wire n_5709;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_4861;
wire n_5799;
wire n_4064;
wire n_4926;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_5266;
wire n_5580;
wire n_4828;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_2726;
wire n_4303;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_4768;
wire n_3717;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_1856;
wire n_2077;
wire n_5691;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_5615;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_5468;
wire n_4730;
wire n_5399;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_5713;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_5550;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_5509;
wire n_5382;
wire n_5659;
wire n_3619;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1867;
wire n_2630;
wire n_2470;
wire n_4446;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_2256;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_5796;
wire n_2806;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_3624;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_5492;
wire n_2378;
wire n_2655;
wire n_4600;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_3568;
wire n_3850;
wire n_5770;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_4745;
wire n_5642;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_4792;
wire n_3842;
wire n_2031;
wire n_4878;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_3599;
wire n_5543;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_4773;
wire n_5654;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_4427;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_5692;
wire n_4800;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_3252;
wire n_3253;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_5080;
wire n_3128;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_5690;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_5801;
wire n_3037;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_3053;
wire n_1808;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_5125;
wire n_2650;
wire n_5652;
wire n_5499;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_4280;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_4097;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_5455;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_4419;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_3848;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_2745;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_4830;
wire n_4706;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_2783;
wire n_3188;
wire n_3243;
wire n_2462;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_2270;
wire n_5049;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_5592;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_5278;
wire n_5157;
wire n_3314;
wire n_2100;
wire n_3525;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_1905;
wire n_3466;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_3636;
wire n_2327;
wire n_5516;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_3637;
wire n_4574;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_3236;
wire n_2755;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_5570;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_3249;
wire n_2722;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_5486;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1692;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3501;
wire n_3475;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_2699;
wire n_1828;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_5804;
wire n_3134;
wire n_3115;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5682;
wire n_5387;
wire n_5557;
wire n_2458;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_3307;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_5681;
wire n_4901;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_4040;
wire n_2406;
wire n_2141;
wire n_5316;
wire n_5703;
wire n_3930;
wire n_4943;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_2172;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_4530;
wire n_2021;
wire n_4942;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_2417;
wire n_5093;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1872;
wire n_5040;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_5746;
wire n_2045;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1929;
wire n_2369;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_5432;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_5842;
wire n_5814;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_5777;
wire n_4225;
wire n_2565;
wire n_5495;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_5064;
wire n_5610;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_3473;
wire n_1994;
wire n_2566;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_5559;
wire n_2438;
wire n_2914;
wire n_5786;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_4106;
wire n_5737;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_5768;
wire n_3553;
wire n_2465;
wire n_2275;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_5700;
wire n_3699;
wire n_4913;
wire n_2312;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_2042;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1770;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_4089;
wire n_5478;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_3264;
wire n_2010;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_4865;
wire n_2043;
wire n_5832;
wire n_3206;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_5812;
wire n_2540;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_5368;
wire n_4263;
wire n_1819;
wire n_3555;
wire n_3155;
wire n_3110;
wire n_1888;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1958;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_3387;
wire n_5782;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_2183;
wire n_3002;
wire n_4809;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_3301;
wire n_4241;
wire n_1853;
wire n_2324;
wire n_5563;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_2847;
wire n_2557;
wire n_2405;
wire n_4050;
wire n_2647;
wire n_2336;
wire n_5717;
wire n_2521;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1985;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_3626;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_4555;
wire n_5650;
wire n_4969;
wire n_5105;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_3998;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_5022;
wire n_5670;
wire n_3296;
wire n_5276;
wire n_2551;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_3822;
wire n_4163;
wire n_5535;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_3319;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_4372;
wire n_5640;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_2123;
wire n_1697;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_2941;
wire n_5108;
wire n_4032;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_3092;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_3419;
wire n_4478;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_4673;
wire n_2519;
wire n_3415;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_2663;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_2165;
wire n_5547;
wire n_2750;
wire n_2775;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_2684;
wire n_3146;
wire n_3953;
wire n_4588;
wire n_4653;
wire n_4435;
wire n_5604;
wire n_1756;
wire n_5411;
wire n_4019;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_3616;
wire n_5815;
wire n_4191;
wire n_5695;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_2148;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5669;
wire n_5772;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_5603;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_5712;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_2372;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_3546;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_4573;
wire n_5398;
wire n_2589;
wire n_4535;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_3196;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_5270;
wire n_2063;
wire n_5005;
wire n_2475;
wire n_5181;
wire n_3144;
wire n_3244;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_3640;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_5775;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_4867;
wire n_5061;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_2648;
wire n_3212;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1806;
wire n_2023;
wire n_2720;
wire n_2204;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_3956;
wire n_4001;
wire n_2627;
wire n_4422;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_5735;
wire n_2278;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_5752;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_5189;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_2220;
wire n_2577;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_2373;
wire n_3628;
wire n_5454;
wire n_4734;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_2704;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1830;
wire n_2351;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_2536;
wire n_3915;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_2759;
wire n_2361;
wire n_2266;
wire n_4876;
wire n_5813;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_1794;
wire n_4493;
wire n_4924;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_4953;
wire n_2944;
wire n_2348;
wire n_3831;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_3589;
wire n_2066;
wire n_3391;
wire n_1800;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_5236;
wire n_5012;
wire n_3787;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_4173;
wire n_3135;
wire n_5651;
wire n_4630;
wire n_5645;
wire n_3990;
wire n_5766;
wire n_2109;
wire n_2796;
wire n_2507;
wire n_5671;
wire n_4534;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_4494;
wire n_5412;
wire n_2380;
wire n_4786;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_4282;
wire n_3493;
wire n_3774;
wire n_5733;
wire n_2910;
wire n_3268;
wire n_1785;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_2287;
wire n_5791;
wire n_5727;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_5657;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_3334;
wire n_5602;
wire n_5097;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2203;
wire n_2255;
wire n_5246;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_5666;
wire n_4059;
wire n_4121;
wire n_3290;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_5546;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_2600;
wire n_5626;
wire n_3508;
wire n_4353;
wire n_4787;
wire n_5633;
wire n_5664;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_2440;
wire n_3521;
wire n_2681;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_2909;
wire n_5369;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_3945;
wire n_5817;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_4804;
wire n_5619;
wire n_3965;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_5776;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_4703;
wire n_2419;
wire n_5683;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1430),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_673),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_436),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1575),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1276),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_767),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1239),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1468),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_910),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1541),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1502),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1448),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1137),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1235),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_894),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1569),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_519),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1554),
.Y(n_1698)
);

CKINVDCx16_ASAP7_75t_R g1699 ( 
.A(n_914),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1668),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1507),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_137),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_28),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1197),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_643),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_116),
.Y(n_1706)
);

INVxp33_ASAP7_75t_R g1707 ( 
.A(n_304),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1511),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_244),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_133),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1358),
.Y(n_1711)
);

BUFx5_ASAP7_75t_L g1712 ( 
.A(n_120),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1446),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_734),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_763),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_964),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_191),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_213),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_147),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_568),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_92),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1295),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_18),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_422),
.Y(n_1724)
);

BUFx5_ASAP7_75t_L g1725 ( 
.A(n_970),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1135),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1546),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1234),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1458),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_576),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1488),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_485),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1198),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1592),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_696),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1517),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1164),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1463),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1527),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1474),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_741),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1451),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1425),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1097),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1227),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1622),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_939),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1470),
.Y(n_1748)
);

BUFx10_ASAP7_75t_L g1749 ( 
.A(n_641),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1253),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_83),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1279),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_902),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1483),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_101),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1584),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_752),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_647),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1455),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_945),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_175),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1108),
.Y(n_1762)
);

BUFx10_ASAP7_75t_L g1763 ( 
.A(n_892),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_1381),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_120),
.Y(n_1765)
);

CKINVDCx16_ASAP7_75t_R g1766 ( 
.A(n_620),
.Y(n_1766)
);

BUFx10_ASAP7_75t_L g1767 ( 
.A(n_1504),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1440),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_400),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_509),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1241),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1544),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_848),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1491),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1616),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_505),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_54),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1420),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1579),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1069),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_314),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1260),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_212),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1133),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_102),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1443),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1004),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_129),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_312),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1375),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_217),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1154),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1189),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1666),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1496),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1438),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_91),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1432),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_554),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1228),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_882),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1123),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1515),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1503),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_784),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1578),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_638),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_386),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_695),
.Y(n_1809)
);

BUFx10_ASAP7_75t_L g1810 ( 
.A(n_1557),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1570),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1044),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1098),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1470),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_610),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_364),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1456),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1550),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_812),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_161),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1201),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_642),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1224),
.Y(n_1823)
);

CKINVDCx14_ASAP7_75t_R g1824 ( 
.A(n_1009),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1519),
.Y(n_1825)
);

INVxp33_ASAP7_75t_SL g1826 ( 
.A(n_1324),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1065),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1650),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1442),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1526),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_1106),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_520),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1385),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_431),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1583),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_373),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1132),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_357),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1453),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1313),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1392),
.Y(n_1841)
);

BUFx5_ASAP7_75t_L g1842 ( 
.A(n_532),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_862),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1585),
.Y(n_1844)
);

BUFx5_ASAP7_75t_L g1845 ( 
.A(n_442),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_794),
.Y(n_1846)
);

INVx4_ASAP7_75t_R g1847 ( 
.A(n_697),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1431),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1450),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_600),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_495),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_98),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_120),
.Y(n_1853)
);

CKINVDCx20_ASAP7_75t_R g1854 ( 
.A(n_188),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_213),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1296),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_516),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1600),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1375),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_960),
.Y(n_1860)
);

CKINVDCx20_ASAP7_75t_R g1861 ( 
.A(n_1494),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1540),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_49),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1205),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1382),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_38),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_442),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1476),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_545),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1623),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_964),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_613),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1651),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1632),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1099),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_963),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1391),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_193),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_655),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_690),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1007),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1452),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1536),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1542),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_816),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_668),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_105),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_695),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1291),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1134),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_11),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_66),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1234),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1672),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1627),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_95),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1225),
.Y(n_1897)
);

CKINVDCx16_ASAP7_75t_R g1898 ( 
.A(n_1444),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1353),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1571),
.Y(n_1900)
);

BUFx2_ASAP7_75t_SL g1901 ( 
.A(n_1674),
.Y(n_1901)
);

CKINVDCx16_ASAP7_75t_R g1902 ( 
.A(n_1523),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1437),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_467),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1136),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_99),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_839),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_902),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_710),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1495),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1574),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_949),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_467),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_282),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1579),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_513),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_663),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1021),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1303),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_289),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_987),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1143),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1479),
.Y(n_1923)
);

BUFx8_ASAP7_75t_SL g1924 ( 
.A(n_1237),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_204),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_792),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1498),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_100),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1102),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_165),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1555),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_843),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_760),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_14),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_821),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1567),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_443),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1238),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1368),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_479),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1549),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_728),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1323),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_592),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_154),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1563),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_385),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1301),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_605),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_431),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_572),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_140),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1386),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_781),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1516),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1364),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1421),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1357),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_233),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1120),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1480),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_11),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1051),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_725),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_841),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1341),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_858),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1475),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_73),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1330),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1447),
.Y(n_1971)
);

INVx4_ASAP7_75t_R g1972 ( 
.A(n_1520),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_769),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_944),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1521),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1198),
.Y(n_1976)
);

BUFx2_ASAP7_75t_L g1977 ( 
.A(n_1680),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1624),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1199),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1137),
.Y(n_1980)
);

CKINVDCx16_ASAP7_75t_R g1981 ( 
.A(n_720),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_929),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_914),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_779),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1029),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1339),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_997),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_573),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_337),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1426),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1525),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_569),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_989),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_856),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1423),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1505),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_657),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_596),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1259),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_925),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1581),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_333),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1256),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1547),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_970),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1464),
.Y(n_2006)
);

CKINVDCx16_ASAP7_75t_R g2007 ( 
.A(n_966),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1509),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_577),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_213),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1528),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1415),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1219),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_31),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_173),
.Y(n_2015)
);

CKINVDCx16_ASAP7_75t_R g2016 ( 
.A(n_261),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1226),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_757),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1435),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_811),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_753),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1286),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_95),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_953),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1440),
.Y(n_2025)
);

CKINVDCx11_ASAP7_75t_R g2026 ( 
.A(n_1200),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1262),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1066),
.Y(n_2028)
);

INVx2_ASAP7_75t_SL g2029 ( 
.A(n_1324),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_555),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1429),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_28),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_210),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_908),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_32),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_152),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1607),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1473),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_78),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_600),
.Y(n_2040)
);

INVx1_ASAP7_75t_SL g2041 ( 
.A(n_1505),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_849),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_79),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_473),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_822),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1401),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1636),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1566),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_363),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1465),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1299),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1495),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_956),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1576),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_901),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_892),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_348),
.Y(n_2057)
);

CKINVDCx20_ASAP7_75t_R g2058 ( 
.A(n_1141),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1211),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_402),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_715),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1487),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1072),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_726),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_885),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1467),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_240),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1461),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_747),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_837),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_231),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_785),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1472),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1459),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1160),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_995),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1373),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_568),
.Y(n_2078)
);

CKINVDCx20_ASAP7_75t_R g2079 ( 
.A(n_780),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_33),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1485),
.Y(n_2081)
);

CKINVDCx16_ASAP7_75t_R g2082 ( 
.A(n_1053),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_696),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_398),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_962),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1513),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_1289),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1302),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1508),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_701),
.Y(n_2090)
);

BUFx10_ASAP7_75t_L g2091 ( 
.A(n_1629),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_380),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1225),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1561),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_257),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1600),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1092),
.Y(n_2097)
);

INVxp33_ASAP7_75t_R g2098 ( 
.A(n_704),
.Y(n_2098)
);

BUFx2_ASAP7_75t_L g2099 ( 
.A(n_223),
.Y(n_2099)
);

BUFx2_ASAP7_75t_L g2100 ( 
.A(n_1541),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_819),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1478),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_550),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_203),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1427),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_580),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1288),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_998),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1543),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1679),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_1545),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_1072),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_758),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_1558),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1377),
.Y(n_2115)
);

CKINVDCx20_ASAP7_75t_R g2116 ( 
.A(n_1129),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_1345),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1531),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1565),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_465),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_588),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_1333),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_298),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_204),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_746),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_1532),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1044),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_1607),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_820),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1273),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_351),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1288),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1481),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_360),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1229),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1591),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_647),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_470),
.Y(n_2138)
);

CKINVDCx20_ASAP7_75t_R g2139 ( 
.A(n_478),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1192),
.Y(n_2140)
);

INVx1_ASAP7_75t_SL g2141 ( 
.A(n_834),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_476),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1590),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1218),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_481),
.Y(n_2145)
);

CKINVDCx20_ASAP7_75t_R g2146 ( 
.A(n_1493),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_638),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1482),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_941),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_890),
.Y(n_2150)
);

CKINVDCx20_ASAP7_75t_R g2151 ( 
.A(n_1021),
.Y(n_2151)
);

BUFx10_ASAP7_75t_L g2152 ( 
.A(n_1430),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_468),
.Y(n_2153)
);

BUFx10_ASAP7_75t_L g2154 ( 
.A(n_1025),
.Y(n_2154)
);

BUFx8_ASAP7_75t_SL g2155 ( 
.A(n_408),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_60),
.Y(n_2156)
);

BUFx2_ASAP7_75t_L g2157 ( 
.A(n_1216),
.Y(n_2157)
);

CKINVDCx20_ASAP7_75t_R g2158 ( 
.A(n_1083),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1506),
.Y(n_2159)
);

BUFx2_ASAP7_75t_L g2160 ( 
.A(n_481),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_633),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_272),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1060),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1564),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1532),
.Y(n_2165)
);

CKINVDCx16_ASAP7_75t_R g2166 ( 
.A(n_1153),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1439),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_166),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1447),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_709),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1559),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1209),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1210),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1380),
.Y(n_2174)
);

INVxp67_ASAP7_75t_L g2175 ( 
.A(n_1543),
.Y(n_2175)
);

CKINVDCx16_ASAP7_75t_R g2176 ( 
.A(n_1197),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_364),
.Y(n_2177)
);

INVx1_ASAP7_75t_SL g2178 ( 
.A(n_637),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1537),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1489),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_940),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1114),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1012),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_551),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_749),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_366),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_290),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_614),
.Y(n_2188)
);

INVx1_ASAP7_75t_SL g2189 ( 
.A(n_1040),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_330),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_962),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_721),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_181),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1531),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_896),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1094),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_147),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1348),
.Y(n_2198)
);

CKINVDCx16_ASAP7_75t_R g2199 ( 
.A(n_1560),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_153),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_1672),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1436),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1466),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_1599),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_939),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_335),
.Y(n_2206)
);

CKINVDCx16_ASAP7_75t_R g2207 ( 
.A(n_472),
.Y(n_2207)
);

CKINVDCx20_ASAP7_75t_R g2208 ( 
.A(n_545),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1065),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1484),
.Y(n_2210)
);

BUFx10_ASAP7_75t_L g2211 ( 
.A(n_1669),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_866),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1645),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_700),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_204),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1561),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_138),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1553),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_451),
.Y(n_2219)
);

BUFx6f_ASAP7_75t_L g2220 ( 
.A(n_1325),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1217),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1067),
.Y(n_2222)
);

CKINVDCx20_ASAP7_75t_R g2223 ( 
.A(n_826),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1165),
.Y(n_2224)
);

CKINVDCx20_ASAP7_75t_R g2225 ( 
.A(n_897),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_1492),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_971),
.Y(n_2227)
);

CKINVDCx20_ASAP7_75t_R g2228 ( 
.A(n_1555),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_592),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1454),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_1041),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_783),
.Y(n_2232)
);

BUFx5_ASAP7_75t_L g2233 ( 
.A(n_532),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1303),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_161),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1127),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1424),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1631),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_265),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_271),
.Y(n_2240)
);

BUFx10_ASAP7_75t_L g2241 ( 
.A(n_933),
.Y(n_2241)
);

BUFx2_ASAP7_75t_SL g2242 ( 
.A(n_1471),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_862),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1552),
.Y(n_2244)
);

CKINVDCx20_ASAP7_75t_R g2245 ( 
.A(n_228),
.Y(n_2245)
);

CKINVDCx16_ASAP7_75t_R g2246 ( 
.A(n_1441),
.Y(n_2246)
);

HB1xp67_ASAP7_75t_L g2247 ( 
.A(n_173),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_823),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_356),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1460),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1567),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_526),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1630),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1242),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1434),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1343),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_1487),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1422),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_1016),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1100),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1246),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_69),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1181),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1071),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1094),
.Y(n_2265)
);

BUFx10_ASAP7_75t_L g2266 ( 
.A(n_73),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_241),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_1499),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_609),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1254),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_896),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_620),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_745),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_136),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_489),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1457),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_166),
.Y(n_2277)
);

BUFx3_ASAP7_75t_L g2278 ( 
.A(n_1084),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_501),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1538),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_1350),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_293),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_378),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1362),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1649),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_1275),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_342),
.Y(n_2287)
);

BUFx5_ASAP7_75t_L g2288 ( 
.A(n_1533),
.Y(n_2288)
);

BUFx2_ASAP7_75t_L g2289 ( 
.A(n_886),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1160),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1454),
.Y(n_2291)
);

INVx2_ASAP7_75t_SL g2292 ( 
.A(n_933),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_452),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_252),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1381),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_106),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_210),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1415),
.Y(n_2298)
);

CKINVDCx16_ASAP7_75t_R g2299 ( 
.A(n_299),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_121),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_633),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_596),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1163),
.Y(n_2303)
);

BUFx5_ASAP7_75t_L g2304 ( 
.A(n_1562),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1521),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_1425),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1220),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_274),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1015),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_343),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_74),
.Y(n_2311)
);

CKINVDCx20_ASAP7_75t_R g2312 ( 
.A(n_1417),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_98),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_726),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_704),
.Y(n_2315)
);

INVx2_ASAP7_75t_SL g2316 ( 
.A(n_318),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_700),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_258),
.Y(n_2318)
);

INVxp67_ASAP7_75t_L g2319 ( 
.A(n_815),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_336),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_953),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_405),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_1530),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1011),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1291),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_268),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1245),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_880),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_1629),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_733),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_80),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_1510),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1033),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_1262),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_1069),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1574),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_797),
.Y(n_2337)
);

CKINVDCx16_ASAP7_75t_R g2338 ( 
.A(n_1577),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1581),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_503),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_1462),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1079),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1501),
.Y(n_2343)
);

INVxp67_ASAP7_75t_L g2344 ( 
.A(n_1644),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_1588),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_5),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1084),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_1321),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1511),
.Y(n_2349)
);

BUFx8_ASAP7_75t_SL g2350 ( 
.A(n_1575),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_802),
.Y(n_2351)
);

CKINVDCx20_ASAP7_75t_R g2352 ( 
.A(n_479),
.Y(n_2352)
);

INVx2_ASAP7_75t_SL g2353 ( 
.A(n_1207),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1556),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_4),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_932),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_885),
.Y(n_2357)
);

BUFx8_ASAP7_75t_SL g2358 ( 
.A(n_99),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_667),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1260),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1512),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_512),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1041),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_1643),
.Y(n_2364)
);

BUFx6f_ASAP7_75t_L g2365 ( 
.A(n_1469),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_443),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_77),
.Y(n_2367)
);

CKINVDCx20_ASAP7_75t_R g2368 ( 
.A(n_296),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_631),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_340),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_215),
.Y(n_2371)
);

BUFx2_ASAP7_75t_L g2372 ( 
.A(n_1428),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1476),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1190),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_427),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_198),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_688),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_624),
.Y(n_2378)
);

BUFx2_ASAP7_75t_SL g2379 ( 
.A(n_539),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_317),
.Y(n_2380)
);

INVxp67_ASAP7_75t_L g2381 ( 
.A(n_1593),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_1134),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1088),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_1625),
.Y(n_2384)
);

BUFx3_ASAP7_75t_L g2385 ( 
.A(n_411),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1540),
.Y(n_2386)
);

INVx1_ASAP7_75t_SL g2387 ( 
.A(n_1297),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_749),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_298),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_631),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_994),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_1572),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_42),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_1490),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_1100),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_192),
.Y(n_2396)
);

BUFx10_ASAP7_75t_L g2397 ( 
.A(n_961),
.Y(n_2397)
);

CKINVDCx16_ASAP7_75t_R g2398 ( 
.A(n_1662),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_1334),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_961),
.Y(n_2400)
);

CKINVDCx16_ASAP7_75t_R g2401 ( 
.A(n_1241),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_1582),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_1587),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_137),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_181),
.Y(n_2405)
);

INVxp33_ASAP7_75t_R g2406 ( 
.A(n_787),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1539),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1449),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_515),
.Y(n_2409)
);

CKINVDCx20_ASAP7_75t_R g2410 ( 
.A(n_1445),
.Y(n_2410)
);

INVx1_ASAP7_75t_SL g2411 ( 
.A(n_64),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_1488),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_1477),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_499),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_932),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1064),
.Y(n_2416)
);

CKINVDCx5p33_ASAP7_75t_R g2417 ( 
.A(n_1008),
.Y(n_2417)
);

BUFx6f_ASAP7_75t_L g2418 ( 
.A(n_1003),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_748),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_250),
.Y(n_2420)
);

BUFx2_ASAP7_75t_L g2421 ( 
.A(n_1307),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_140),
.Y(n_2422)
);

CKINVDCx20_ASAP7_75t_R g2423 ( 
.A(n_712),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_82),
.Y(n_2424)
);

CKINVDCx16_ASAP7_75t_R g2425 ( 
.A(n_187),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1500),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_383),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_1141),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_563),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1085),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_533),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_549),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_1548),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_1542),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_1079),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_1144),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_1081),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_211),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_824),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_519),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_871),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_447),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_721),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_1458),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_956),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_L g2446 ( 
.A(n_736),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_1619),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_1252),
.Y(n_2448)
);

BUFx6f_ASAP7_75t_L g2449 ( 
.A(n_512),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_126),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_242),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_919),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1066),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_1124),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_861),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_1186),
.Y(n_2456)
);

INVx1_ASAP7_75t_SL g2457 ( 
.A(n_1231),
.Y(n_2457)
);

BUFx3_ASAP7_75t_L g2458 ( 
.A(n_495),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_55),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_1082),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_74),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_922),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_252),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_1433),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_1649),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_1444),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_729),
.Y(n_2467)
);

BUFx6f_ASAP7_75t_L g2468 ( 
.A(n_919),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1659),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_1566),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_1240),
.Y(n_2471)
);

CKINVDCx20_ASAP7_75t_R g2472 ( 
.A(n_1580),
.Y(n_2472)
);

CKINVDCx16_ASAP7_75t_R g2473 ( 
.A(n_1497),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_1573),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_1409),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_954),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_35),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_1076),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_1280),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_125),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_743),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_829),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_59),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_1277),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_573),
.Y(n_2485)
);

CKINVDCx20_ASAP7_75t_R g2486 ( 
.A(n_1522),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_163),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_263),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1000),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_1423),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_551),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_1107),
.Y(n_2492)
);

CKINVDCx20_ASAP7_75t_R g2493 ( 
.A(n_762),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_1615),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_1210),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_806),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_616),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_1630),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_1435),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_1551),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_167),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_1057),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_1027),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_1535),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_414),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_610),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_1524),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_1293),
.Y(n_2508)
);

CKINVDCx16_ASAP7_75t_R g2509 ( 
.A(n_37),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_1514),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_375),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_50),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_1302),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_1316),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_582),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_1074),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_1518),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_1496),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_1224),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_799),
.Y(n_2520)
);

BUFx6f_ASAP7_75t_L g2521 ( 
.A(n_1405),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_1017),
.Y(n_2522)
);

INVx1_ASAP7_75t_SL g2523 ( 
.A(n_946),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_1390),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_189),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_911),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_1045),
.Y(n_2527)
);

CKINVDCx20_ASAP7_75t_R g2528 ( 
.A(n_1534),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1568),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_537),
.Y(n_2530)
);

HB1xp67_ASAP7_75t_L g2531 ( 
.A(n_1169),
.Y(n_2531)
);

BUFx5_ASAP7_75t_L g2532 ( 
.A(n_1235),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_1556),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_397),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_1486),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_1161),
.Y(n_2536)
);

BUFx5_ASAP7_75t_L g2537 ( 
.A(n_72),
.Y(n_2537)
);

CKINVDCx20_ASAP7_75t_R g2538 ( 
.A(n_173),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_1242),
.Y(n_2539)
);

CKINVDCx20_ASAP7_75t_R g2540 ( 
.A(n_1529),
.Y(n_2540)
);

INVx1_ASAP7_75t_SL g2541 ( 
.A(n_25),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_229),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_1032),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_1712),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1712),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_1712),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_1712),
.Y(n_2547)
);

CKINVDCx20_ASAP7_75t_R g2548 ( 
.A(n_1824),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_1712),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2537),
.Y(n_2550)
);

INVx3_ASAP7_75t_L g2551 ( 
.A(n_1704),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2537),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2537),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2537),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_1725),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_1725),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_2358),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2016),
.Y(n_2558)
);

CKINVDCx20_ASAP7_75t_R g2559 ( 
.A(n_1699),
.Y(n_2559)
);

INVxp33_ASAP7_75t_SL g2560 ( 
.A(n_2039),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_1725),
.Y(n_2561)
);

INVxp67_ASAP7_75t_L g2562 ( 
.A(n_2071),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_1725),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_1725),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2099),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_1842),
.Y(n_2566)
);

BUFx3_ASAP7_75t_L g2567 ( 
.A(n_1723),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_1842),
.Y(n_2568)
);

INVxp67_ASAP7_75t_L g2569 ( 
.A(n_2123),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_1842),
.Y(n_2570)
);

INVxp67_ASAP7_75t_L g2571 ( 
.A(n_2247),
.Y(n_2571)
);

INVxp67_ASAP7_75t_SL g2572 ( 
.A(n_2355),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1845),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_1920),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1845),
.Y(n_2575)
);

INVxp67_ASAP7_75t_L g2576 ( 
.A(n_1760),
.Y(n_2576)
);

INVxp33_ASAP7_75t_L g2577 ( 
.A(n_1688),
.Y(n_2577)
);

CKINVDCx20_ASAP7_75t_R g2578 ( 
.A(n_1766),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_1845),
.Y(n_2579)
);

INVxp67_ASAP7_75t_SL g2580 ( 
.A(n_1905),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1845),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2233),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2233),
.Y(n_2583)
);

INVxp33_ASAP7_75t_SL g2584 ( 
.A(n_1865),
.Y(n_2584)
);

INVxp67_ASAP7_75t_L g2585 ( 
.A(n_1812),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_2026),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2233),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2233),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2288),
.Y(n_2589)
);

INVxp67_ASAP7_75t_SL g2590 ( 
.A(n_1905),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2288),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2288),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2288),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2288),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2304),
.Y(n_2595)
);

INVxp33_ASAP7_75t_SL g2596 ( 
.A(n_2065),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2304),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2304),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2304),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2304),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_1924),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2532),
.Y(n_2602)
);

CKINVDCx20_ASAP7_75t_R g2603 ( 
.A(n_1898),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2532),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2532),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2266),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_2155),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2532),
.Y(n_2608)
);

CKINVDCx20_ASAP7_75t_R g2609 ( 
.A(n_1902),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2532),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2542),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1702),
.Y(n_2612)
);

CKINVDCx20_ASAP7_75t_R g2613 ( 
.A(n_1981),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_1718),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2350),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2299),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_1719),
.Y(n_2617)
);

CKINVDCx20_ASAP7_75t_R g2618 ( 
.A(n_2007),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2425),
.Y(n_2619)
);

BUFx3_ASAP7_75t_L g2620 ( 
.A(n_1930),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_1887),
.Y(n_2621)
);

CKINVDCx20_ASAP7_75t_R g2622 ( 
.A(n_2082),
.Y(n_2622)
);

INVxp67_ASAP7_75t_SL g2623 ( 
.A(n_2128),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_1891),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1892),
.Y(n_2625)
);

CKINVDCx20_ASAP7_75t_R g2626 ( 
.A(n_2166),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_1906),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_1914),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_1928),
.Y(n_2629)
);

INVxp67_ASAP7_75t_SL g2630 ( 
.A(n_2128),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_1945),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2509),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2176),
.Y(n_2633)
);

CKINVDCx20_ASAP7_75t_R g2634 ( 
.A(n_2199),
.Y(n_2634)
);

INVxp67_ASAP7_75t_SL g2635 ( 
.A(n_2499),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_1959),
.Y(n_2636)
);

CKINVDCx14_ASAP7_75t_R g2637 ( 
.A(n_1888),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_1969),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2207),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2010),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_2246),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2015),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2033),
.Y(n_2643)
);

INVx1_ASAP7_75t_SL g2644 ( 
.A(n_1947),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_2338),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2036),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2398),
.Y(n_2647)
);

INVxp67_ASAP7_75t_SL g2648 ( 
.A(n_2499),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2067),
.Y(n_2649)
);

CKINVDCx20_ASAP7_75t_R g2650 ( 
.A(n_2401),
.Y(n_2650)
);

INVxp33_ASAP7_75t_SL g2651 ( 
.A(n_2226),
.Y(n_2651)
);

INVx2_ASAP7_75t_SL g2652 ( 
.A(n_2266),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2080),
.Y(n_2653)
);

INVx4_ASAP7_75t_R g2654 ( 
.A(n_1684),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2095),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2104),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2124),
.Y(n_2657)
);

CKINVDCx16_ASAP7_75t_R g2658 ( 
.A(n_2473),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2131),
.Y(n_2659)
);

INVxp33_ASAP7_75t_L g2660 ( 
.A(n_2248),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2162),
.Y(n_2661)
);

BUFx3_ASAP7_75t_L g2662 ( 
.A(n_2326),
.Y(n_2662)
);

BUFx2_ASAP7_75t_SL g2663 ( 
.A(n_1727),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2200),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2206),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2235),
.Y(n_2666)
);

INVxp67_ASAP7_75t_L g2667 ( 
.A(n_1974),
.Y(n_2667)
);

INVxp67_ASAP7_75t_SL g2668 ( 
.A(n_2524),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2249),
.Y(n_2669)
);

INVx1_ASAP7_75t_SL g2670 ( 
.A(n_1977),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_1706),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2262),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2282),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2294),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2300),
.Y(n_2675)
);

CKINVDCx14_ASAP7_75t_R g2676 ( 
.A(n_2004),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2308),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2313),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2320),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2331),
.Y(n_2680)
);

INVx1_ASAP7_75t_SL g2681 ( 
.A(n_2100),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2405),
.Y(n_2682)
);

CKINVDCx20_ASAP7_75t_R g2683 ( 
.A(n_1746),
.Y(n_2683)
);

INVx1_ASAP7_75t_SL g2684 ( 
.A(n_2112),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_2157),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2346),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_1709),
.Y(n_2687)
);

CKINVDCx14_ASAP7_75t_R g2688 ( 
.A(n_2160),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2370),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2371),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2393),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2450),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2459),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2463),
.Y(n_2694)
);

INVxp67_ASAP7_75t_SL g2695 ( 
.A(n_1920),
.Y(n_2695)
);

CKINVDCx16_ASAP7_75t_R g2696 ( 
.A(n_1749),
.Y(n_2696)
);

INVxp67_ASAP7_75t_L g2697 ( 
.A(n_2289),
.Y(n_2697)
);

INVxp67_ASAP7_75t_L g2698 ( 
.A(n_2372),
.Y(n_2698)
);

CKINVDCx16_ASAP7_75t_R g2699 ( 
.A(n_1749),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2480),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_1717),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2366),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_1920),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_1721),
.Y(n_2704)
);

CKINVDCx5p33_ASAP7_75t_R g2705 ( 
.A(n_1751),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_1820),
.Y(n_2706)
);

INVxp67_ASAP7_75t_L g2707 ( 
.A(n_2421),
.Y(n_2707)
);

INVxp67_ASAP7_75t_SL g2708 ( 
.A(n_2531),
.Y(n_2708)
);

INVxp67_ASAP7_75t_SL g2709 ( 
.A(n_1704),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_1852),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_1755),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_1878),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_1764),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2190),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2501),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_1761),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_1765),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_1704),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_1708),
.Y(n_2719)
);

CKINVDCx20_ASAP7_75t_R g2720 ( 
.A(n_1769),
.Y(n_2720)
);

INVxp33_ASAP7_75t_SL g2721 ( 
.A(n_1777),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_1781),
.Y(n_2722)
);

INVxp67_ASAP7_75t_SL g2723 ( 
.A(n_1708),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_1785),
.Y(n_2724)
);

CKINVDCx20_ASAP7_75t_R g2725 ( 
.A(n_1771),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_1708),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_1809),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_1809),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_1788),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_1789),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_1818),
.Y(n_2731)
);

CKINVDCx20_ASAP7_75t_R g2732 ( 
.A(n_1782),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_1818),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_1797),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_1822),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_1822),
.Y(n_2736)
);

CKINVDCx16_ASAP7_75t_R g2737 ( 
.A(n_1763),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_1870),
.Y(n_2738)
);

CKINVDCx20_ASAP7_75t_R g2739 ( 
.A(n_1790),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_1870),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_1838),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_1893),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_1853),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_1855),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_1863),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_1893),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1893),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_1907),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_1866),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_1907),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_1896),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_1925),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_1826),
.B(n_0),
.Y(n_2753)
);

INVxp67_ASAP7_75t_SL g2754 ( 
.A(n_1941),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_1934),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_1997),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_1997),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2049),
.Y(n_2758)
);

INVxp67_ASAP7_75t_SL g2759 ( 
.A(n_2049),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2059),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2059),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2709),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2708),
.B(n_1731),
.Y(n_2763)
);

INVx4_ASAP7_75t_L g2764 ( 
.A(n_2671),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2658),
.B(n_2696),
.Y(n_2765)
);

BUFx3_ASAP7_75t_L g2766 ( 
.A(n_2567),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2723),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2738),
.Y(n_2768)
);

BUFx2_ASAP7_75t_L g2769 ( 
.A(n_2559),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2572),
.B(n_1802),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2580),
.B(n_2126),
.Y(n_2771)
);

OAI22x1_ASAP7_75t_L g2772 ( 
.A1(n_2644),
.A2(n_1962),
.B1(n_1989),
.B2(n_1952),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2633),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2558),
.Y(n_2774)
);

AND2x2_ASAP7_75t_SL g2775 ( 
.A(n_2753),
.B(n_2126),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2590),
.B(n_1881),
.Y(n_2776)
);

OA21x2_ASAP7_75t_L g2777 ( 
.A1(n_2544),
.A2(n_1693),
.B(n_1686),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2574),
.Y(n_2778)
);

BUFx12f_ASAP7_75t_L g2779 ( 
.A(n_2601),
.Y(n_2779)
);

CKINVDCx20_ASAP7_75t_R g2780 ( 
.A(n_2683),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2574),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2623),
.B(n_2126),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2630),
.B(n_2635),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2546),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2584),
.A2(n_2002),
.B1(n_2023),
.B2(n_2014),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2703),
.Y(n_2786)
);

BUFx3_ASAP7_75t_L g2787 ( 
.A(n_2620),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_2687),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2754),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2759),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2695),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2639),
.Y(n_2792)
);

BUFx3_ASAP7_75t_L g2793 ( 
.A(n_2662),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2648),
.B(n_1908),
.Y(n_2794)
);

INVx6_ASAP7_75t_L g2795 ( 
.A(n_2682),
.Y(n_2795)
);

BUFx12f_ASAP7_75t_L g2796 ( 
.A(n_2607),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2562),
.B(n_1910),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2545),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2596),
.A2(n_2035),
.B1(n_2057),
.B2(n_2043),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2547),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2551),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2578),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2565),
.B(n_1916),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2668),
.B(n_1943),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2549),
.Y(n_2805)
);

AND2x6_ASAP7_75t_L g2806 ( 
.A(n_2670),
.B(n_1703),
.Y(n_2806)
);

OAI22x1_ASAP7_75t_SL g2807 ( 
.A1(n_2713),
.A2(n_1710),
.B1(n_1854),
.B2(n_1783),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2672),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2550),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2689),
.Y(n_2810)
);

CKINVDCx6p67_ASAP7_75t_R g2811 ( 
.A(n_2548),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2663),
.B(n_2205),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_2710),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_SL g2814 ( 
.A(n_2681),
.B(n_1763),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_2615),
.Y(n_2815)
);

BUFx2_ASAP7_75t_L g2816 ( 
.A(n_2603),
.Y(n_2816)
);

AND2x4_ASAP7_75t_L g2817 ( 
.A(n_2569),
.B(n_1982),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2552),
.Y(n_2818)
);

HB1xp67_ASAP7_75t_L g2819 ( 
.A(n_2641),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2553),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2554),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2718),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2719),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2726),
.Y(n_2824)
);

AND2x2_ASAP7_75t_SL g2825 ( 
.A(n_2699),
.B(n_2205),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2727),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2701),
.Y(n_2827)
);

BUFx8_ASAP7_75t_L g2828 ( 
.A(n_2606),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2728),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2576),
.B(n_1986),
.Y(n_2830)
);

BUFx12f_ASAP7_75t_L g2831 ( 
.A(n_2586),
.Y(n_2831)
);

INVx3_ASAP7_75t_L g2832 ( 
.A(n_2731),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2704),
.B(n_2220),
.Y(n_2833)
);

INVx5_ASAP7_75t_L g2834 ( 
.A(n_2652),
.Y(n_2834)
);

BUFx6f_ASAP7_75t_L g2835 ( 
.A(n_2733),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2735),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2736),
.Y(n_2837)
);

OA21x2_ASAP7_75t_L g2838 ( 
.A1(n_2555),
.A2(n_1738),
.B(n_1730),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2705),
.Y(n_2839)
);

OAI22xp33_ASAP7_75t_R g2840 ( 
.A1(n_2684),
.A2(n_1707),
.B1(n_2032),
.B2(n_1791),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2740),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2742),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2746),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2747),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2711),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2748),
.Y(n_2846)
);

AND2x4_ASAP7_75t_L g2847 ( 
.A(n_2585),
.B(n_2278),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2750),
.Y(n_2848)
);

AND2x2_ASAP7_75t_SL g2849 ( 
.A(n_2737),
.B(n_2220),
.Y(n_2849)
);

NAND2x1p5_ASAP7_75t_L g2850 ( 
.A(n_2611),
.B(n_2220),
.Y(n_2850)
);

CKINVDCx5p33_ASAP7_75t_R g2851 ( 
.A(n_2716),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_2717),
.Y(n_2852)
);

INVx5_ASAP7_75t_L g2853 ( 
.A(n_2556),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2651),
.A2(n_2156),
.B1(n_2187),
.B2(n_2168),
.Y(n_2854)
);

OA21x2_ASAP7_75t_L g2855 ( 
.A1(n_2561),
.A2(n_1807),
.B(n_1762),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2756),
.Y(n_2856)
);

INVx3_ASAP7_75t_L g2857 ( 
.A(n_2757),
.Y(n_2857)
);

INVx3_ASAP7_75t_L g2858 ( 
.A(n_2758),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2721),
.B(n_2277),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2560),
.A2(n_2193),
.B1(n_2215),
.B2(n_2197),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2760),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2637),
.B(n_2676),
.Y(n_2862)
);

AND2x4_ASAP7_75t_L g2863 ( 
.A(n_2667),
.B(n_2332),
.Y(n_2863)
);

BUFx6f_ASAP7_75t_L g2864 ( 
.A(n_2761),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2755),
.B(n_2227),
.Y(n_2865)
);

BUFx3_ASAP7_75t_L g2866 ( 
.A(n_2563),
.Y(n_2866)
);

AND2x6_ASAP7_75t_L g2867 ( 
.A(n_2612),
.B(n_2411),
.Y(n_2867)
);

INVxp33_ASAP7_75t_SL g2868 ( 
.A(n_2645),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2566),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2647),
.Y(n_2870)
);

INVx5_ASAP7_75t_L g2871 ( 
.A(n_2564),
.Y(n_2871)
);

OAI21x1_ASAP7_75t_L g2872 ( 
.A1(n_2568),
.A2(n_1819),
.B(n_1813),
.Y(n_2872)
);

BUFx6f_ASAP7_75t_L g2873 ( 
.A(n_2614),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2600),
.Y(n_2874)
);

XNOR2x2_ASAP7_75t_L g2875 ( 
.A(n_2617),
.B(n_2541),
.Y(n_2875)
);

CKINVDCx6p67_ASAP7_75t_R g2876 ( 
.A(n_2609),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2621),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2616),
.A2(n_2217),
.B1(n_2240),
.B2(n_2239),
.Y(n_2878)
);

BUFx8_ASAP7_75t_L g2879 ( 
.A(n_2624),
.Y(n_2879)
);

NOR2x1_ASAP7_75t_L g2880 ( 
.A(n_2570),
.B(n_2385),
.Y(n_2880)
);

BUFx6f_ASAP7_75t_L g2881 ( 
.A(n_2625),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2573),
.Y(n_2882)
);

OAI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2575),
.A2(n_1879),
.B(n_1874),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2619),
.B(n_2227),
.Y(n_2884)
);

AOI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2688),
.A2(n_2267),
.B1(n_2287),
.B2(n_2274),
.Y(n_2885)
);

OA21x2_ASAP7_75t_L g2886 ( 
.A1(n_2579),
.A2(n_1938),
.B(n_1913),
.Y(n_2886)
);

BUFx6f_ASAP7_75t_L g2887 ( 
.A(n_2627),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2581),
.Y(n_2888)
);

NOR2xp33_ASAP7_75t_L g2889 ( 
.A(n_2722),
.B(n_2316),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2628),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2582),
.Y(n_2891)
);

INVx2_ASAP7_75t_SL g2892 ( 
.A(n_2724),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_2729),
.Y(n_2893)
);

OAI21x1_ASAP7_75t_L g2894 ( 
.A1(n_2583),
.A2(n_1967),
.B(n_1963),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2752),
.B(n_2227),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2730),
.B(n_2365),
.Y(n_2896)
);

BUFx12f_ASAP7_75t_L g2897 ( 
.A(n_2734),
.Y(n_2897)
);

BUFx2_ASAP7_75t_L g2898 ( 
.A(n_2613),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2741),
.B(n_2365),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2751),
.B(n_2365),
.Y(n_2900)
);

CKINVDCx16_ASAP7_75t_R g2901 ( 
.A(n_2618),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2743),
.B(n_2744),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_L g2903 ( 
.A(n_2629),
.Y(n_2903)
);

OA21x2_ASAP7_75t_L g2904 ( 
.A1(n_2587),
.A2(n_2069),
.B(n_2056),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2745),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2588),
.Y(n_2906)
);

INVx3_ASAP7_75t_L g2907 ( 
.A(n_2631),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_2636),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2685),
.A2(n_2297),
.B1(n_2310),
.B2(n_2296),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2589),
.Y(n_2910)
);

BUFx6f_ASAP7_75t_L g2911 ( 
.A(n_2638),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2591),
.Y(n_2912)
);

AOI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2697),
.A2(n_2311),
.B1(n_2367),
.B2(n_2318),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2749),
.B(n_2592),
.Y(n_2914)
);

BUFx2_ASAP7_75t_L g2915 ( 
.A(n_2622),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2698),
.A2(n_2376),
.B1(n_2389),
.B2(n_2380),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2577),
.B(n_2402),
.Y(n_2917)
);

HB1xp67_ASAP7_75t_L g2918 ( 
.A(n_2632),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2593),
.B(n_2594),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2707),
.A2(n_2396),
.B1(n_2420),
.B2(n_2404),
.Y(n_2920)
);

OAI22xp5_ASAP7_75t_SL g2921 ( 
.A1(n_2626),
.A2(n_2368),
.B1(n_2538),
.B2(n_2245),
.Y(n_2921)
);

AND2x2_ASAP7_75t_L g2922 ( 
.A(n_2660),
.B(n_2458),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2595),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2597),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2598),
.Y(n_2925)
);

AND2x4_ASAP7_75t_L g2926 ( 
.A(n_2571),
.B(n_2479),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2599),
.Y(n_2927)
);

INVx3_ASAP7_75t_L g2928 ( 
.A(n_2640),
.Y(n_2928)
);

INVx3_ASAP7_75t_L g2929 ( 
.A(n_2642),
.Y(n_2929)
);

BUFx6f_ASAP7_75t_L g2930 ( 
.A(n_2643),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2646),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2602),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2604),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2605),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2702),
.B(n_1923),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2873),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_2827),
.Y(n_2937)
);

BUFx2_ASAP7_75t_L g2938 ( 
.A(n_2806),
.Y(n_2938)
);

CKINVDCx5p33_ASAP7_75t_R g2939 ( 
.A(n_2839),
.Y(n_2939)
);

NOR2xp67_ASAP7_75t_L g2940 ( 
.A(n_2764),
.B(n_2557),
.Y(n_2940)
);

CKINVDCx5p33_ASAP7_75t_R g2941 ( 
.A(n_2845),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2881),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_2851),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2887),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_2852),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2778),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2914),
.B(n_2608),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2783),
.B(n_2610),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2903),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_2893),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2866),
.Y(n_2951)
);

INVxp67_ASAP7_75t_L g2952 ( 
.A(n_2814),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_R g2953 ( 
.A(n_2815),
.B(n_2720),
.Y(n_2953)
);

CKINVDCx20_ASAP7_75t_R g2954 ( 
.A(n_2780),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2775),
.A2(n_2175),
.B1(n_2319),
.B2(n_1918),
.Y(n_2955)
);

CKINVDCx5p33_ASAP7_75t_R g2956 ( 
.A(n_2905),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2911),
.Y(n_2957)
);

CKINVDCx5p33_ASAP7_75t_R g2958 ( 
.A(n_2897),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_R g2959 ( 
.A(n_2901),
.B(n_2779),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_R g2960 ( 
.A(n_2796),
.B(n_2725),
.Y(n_2960)
);

CKINVDCx20_ASAP7_75t_R g2961 ( 
.A(n_2876),
.Y(n_2961)
);

CKINVDCx20_ASAP7_75t_R g2962 ( 
.A(n_2811),
.Y(n_2962)
);

CKINVDCx5p33_ASAP7_75t_R g2963 ( 
.A(n_2868),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2833),
.B(n_2649),
.Y(n_2964)
);

CKINVDCx5p33_ASAP7_75t_R g2965 ( 
.A(n_2831),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2930),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2931),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2768),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2862),
.B(n_2653),
.Y(n_2969)
);

CKINVDCx5p33_ASAP7_75t_R g2970 ( 
.A(n_2788),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_2892),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2798),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_2769),
.Y(n_2973)
);

CKINVDCx16_ASAP7_75t_R g2974 ( 
.A(n_2802),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2784),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2874),
.Y(n_2976)
);

CKINVDCx5p33_ASAP7_75t_R g2977 ( 
.A(n_2816),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_R g2978 ( 
.A(n_2898),
.B(n_2732),
.Y(n_2978)
);

CKINVDCx5p33_ASAP7_75t_R g2979 ( 
.A(n_2915),
.Y(n_2979)
);

BUFx3_ASAP7_75t_L g2980 ( 
.A(n_2766),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2902),
.Y(n_2981)
);

CKINVDCx5p33_ASAP7_75t_R g2982 ( 
.A(n_2828),
.Y(n_2982)
);

CKINVDCx20_ASAP7_75t_R g2983 ( 
.A(n_2773),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_2792),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2808),
.Y(n_2985)
);

CKINVDCx5p33_ASAP7_75t_R g2986 ( 
.A(n_2819),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2800),
.Y(n_2987)
);

OAI22xp33_ASAP7_75t_SL g2988 ( 
.A1(n_2865),
.A2(n_2424),
.B1(n_2438),
.B2(n_2422),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_2870),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_2787),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2793),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_2825),
.Y(n_2992)
);

BUFx10_ASAP7_75t_L g2993 ( 
.A(n_2889),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2805),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2895),
.B(n_2634),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2810),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_2917),
.Y(n_2997)
);

HB1xp67_ASAP7_75t_L g2998 ( 
.A(n_2922),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2849),
.Y(n_2999)
);

CKINVDCx5p33_ASAP7_75t_R g3000 ( 
.A(n_2795),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_2896),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2809),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2899),
.B(n_2650),
.Y(n_3003)
);

CKINVDCx20_ASAP7_75t_R g3004 ( 
.A(n_2765),
.Y(n_3004)
);

CKINVDCx20_ASAP7_75t_R g3005 ( 
.A(n_2918),
.Y(n_3005)
);

BUFx2_ASAP7_75t_L g3006 ( 
.A(n_2806),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2786),
.Y(n_3007)
);

CKINVDCx5p33_ASAP7_75t_R g3008 ( 
.A(n_2900),
.Y(n_3008)
);

INVxp67_ASAP7_75t_L g3009 ( 
.A(n_2859),
.Y(n_3009)
);

NOR2xp67_ASAP7_75t_L g3010 ( 
.A(n_2834),
.B(n_2655),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2762),
.B(n_2451),
.Y(n_3011)
);

CKINVDCx20_ASAP7_75t_R g3012 ( 
.A(n_2921),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2885),
.Y(n_3013)
);

CKINVDCx5p33_ASAP7_75t_R g3014 ( 
.A(n_2807),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2776),
.B(n_2656),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2818),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2878),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_R g3018 ( 
.A(n_2791),
.B(n_2739),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2767),
.B(n_2461),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2821),
.Y(n_3020)
);

CKINVDCx20_ASAP7_75t_R g3021 ( 
.A(n_2774),
.Y(n_3021)
);

NOR2xp67_ASAP7_75t_L g3022 ( 
.A(n_2853),
.B(n_2657),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2869),
.Y(n_3023)
);

CKINVDCx20_ASAP7_75t_R g3024 ( 
.A(n_2770),
.Y(n_3024)
);

CKINVDCx5p33_ASAP7_75t_R g3025 ( 
.A(n_2854),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2882),
.Y(n_3026)
);

CKINVDCx20_ASAP7_75t_R g3027 ( 
.A(n_2794),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2888),
.Y(n_3028)
);

NOR2xp67_ASAP7_75t_L g3029 ( 
.A(n_2853),
.B(n_2659),
.Y(n_3029)
);

HB1xp67_ASAP7_75t_L g3030 ( 
.A(n_2812),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_SL g3031 ( 
.A(n_2763),
.B(n_2375),
.Y(n_3031)
);

INVx3_ASAP7_75t_L g3032 ( 
.A(n_2820),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_2804),
.Y(n_3033)
);

CKINVDCx5p33_ASAP7_75t_R g3034 ( 
.A(n_2785),
.Y(n_3034)
);

CKINVDCx5p33_ASAP7_75t_R g3035 ( 
.A(n_2799),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2836),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_2909),
.Y(n_3037)
);

CKINVDCx5p33_ASAP7_75t_R g3038 ( 
.A(n_2860),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2842),
.Y(n_3039)
);

NAND2xp33_ASAP7_75t_R g3040 ( 
.A(n_2935),
.B(n_2797),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2891),
.Y(n_3041)
);

CKINVDCx5p33_ASAP7_75t_R g3042 ( 
.A(n_2875),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2910),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_2913),
.Y(n_3044)
);

NOR2xp67_ASAP7_75t_L g3045 ( 
.A(n_2871),
.B(n_2661),
.Y(n_3045)
);

CKINVDCx5p33_ASAP7_75t_R g3046 ( 
.A(n_2916),
.Y(n_3046)
);

CKINVDCx5p33_ASAP7_75t_R g3047 ( 
.A(n_2920),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2932),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2934),
.Y(n_3049)
);

CKINVDCx20_ASAP7_75t_R g3050 ( 
.A(n_2884),
.Y(n_3050)
);

CKINVDCx5p33_ASAP7_75t_R g3051 ( 
.A(n_2772),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2830),
.B(n_2375),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2789),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_2790),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2843),
.Y(n_3055)
);

CKINVDCx5p33_ASAP7_75t_R g3056 ( 
.A(n_2847),
.Y(n_3056)
);

CKINVDCx5p33_ASAP7_75t_R g3057 ( 
.A(n_2863),
.Y(n_3057)
);

CKINVDCx20_ASAP7_75t_R g3058 ( 
.A(n_2879),
.Y(n_3058)
);

CKINVDCx5p33_ASAP7_75t_R g3059 ( 
.A(n_2803),
.Y(n_3059)
);

BUFx2_ASAP7_75t_L g3060 ( 
.A(n_2867),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_R g3061 ( 
.A(n_2771),
.B(n_1805),
.Y(n_3061)
);

BUFx2_ASAP7_75t_L g3062 ( 
.A(n_2867),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2906),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2912),
.Y(n_3064)
);

CKINVDCx20_ASAP7_75t_R g3065 ( 
.A(n_2782),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2923),
.Y(n_3066)
);

OAI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_2817),
.A2(n_2381),
.B1(n_2344),
.B2(n_2477),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_2926),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2823),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_R g3070 ( 
.A(n_2877),
.B(n_1831),
.Y(n_3070)
);

CKINVDCx20_ASAP7_75t_R g3071 ( 
.A(n_2919),
.Y(n_3071)
);

CKINVDCx5p33_ASAP7_75t_R g3072 ( 
.A(n_2835),
.Y(n_3072)
);

CKINVDCx5p33_ASAP7_75t_R g3073 ( 
.A(n_2844),
.Y(n_3073)
);

AOI21x1_ASAP7_75t_L g3074 ( 
.A1(n_2924),
.A2(n_2665),
.B(n_2664),
.Y(n_3074)
);

BUFx3_ASAP7_75t_L g3075 ( 
.A(n_2777),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_R g3076 ( 
.A(n_2890),
.B(n_1861),
.Y(n_3076)
);

CKINVDCx5p33_ASAP7_75t_R g3077 ( 
.A(n_2864),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2925),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2927),
.Y(n_3079)
);

INVx5_ASAP7_75t_L g3080 ( 
.A(n_2781),
.Y(n_3080)
);

CKINVDCx20_ASAP7_75t_R g3081 ( 
.A(n_2838),
.Y(n_3081)
);

CKINVDCx5p33_ASAP7_75t_R g3082 ( 
.A(n_2907),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2933),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2871),
.B(n_2666),
.Y(n_3084)
);

CKINVDCx5p33_ASAP7_75t_R g3085 ( 
.A(n_2929),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_2908),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2855),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2822),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2886),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2824),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_2928),
.Y(n_3091)
);

CKINVDCx5p33_ASAP7_75t_R g3092 ( 
.A(n_2813),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2880),
.B(n_2418),
.Y(n_3093)
);

AOI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2872),
.A2(n_2673),
.B(n_2669),
.Y(n_3094)
);

CKINVDCx5p33_ASAP7_75t_R g3095 ( 
.A(n_2801),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2829),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2904),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_R g3098 ( 
.A(n_2826),
.B(n_1885),
.Y(n_3098)
);

CKINVDCx6p67_ASAP7_75t_R g3099 ( 
.A(n_2840),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_2837),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2883),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2832),
.B(n_2674),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2841),
.B(n_2675),
.Y(n_3103)
);

CKINVDCx5p33_ASAP7_75t_R g3104 ( 
.A(n_2846),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_2848),
.Y(n_3105)
);

CKINVDCx5p33_ASAP7_75t_R g3106 ( 
.A(n_2856),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_2861),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2894),
.Y(n_3108)
);

BUFx10_ASAP7_75t_L g3109 ( 
.A(n_2850),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2857),
.B(n_2483),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2858),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_2862),
.B(n_2677),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2873),
.Y(n_3113)
);

INVx3_ASAP7_75t_L g3114 ( 
.A(n_2866),
.Y(n_3114)
);

CKINVDCx20_ASAP7_75t_R g3115 ( 
.A(n_2780),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2778),
.Y(n_3116)
);

CKINVDCx5p33_ASAP7_75t_R g3117 ( 
.A(n_2827),
.Y(n_3117)
);

CKINVDCx5p33_ASAP7_75t_R g3118 ( 
.A(n_2827),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_2827),
.Y(n_3119)
);

CKINVDCx20_ASAP7_75t_R g3120 ( 
.A(n_2780),
.Y(n_3120)
);

BUFx6f_ASAP7_75t_L g3121 ( 
.A(n_2781),
.Y(n_3121)
);

INVxp67_ASAP7_75t_SL g3122 ( 
.A(n_3075),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3094),
.Y(n_3123)
);

INVx3_ASAP7_75t_L g3124 ( 
.A(n_3121),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2975),
.Y(n_3125)
);

AND2x4_ASAP7_75t_L g3126 ( 
.A(n_2980),
.B(n_2985),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2976),
.Y(n_3127)
);

BUFx6f_ASAP7_75t_L g3128 ( 
.A(n_3121),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2968),
.Y(n_3129)
);

BUFx6f_ASAP7_75t_L g3130 ( 
.A(n_3121),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2996),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_3033),
.B(n_2418),
.Y(n_3132)
);

NAND2x1p5_ASAP7_75t_L g3133 ( 
.A(n_2997),
.B(n_2678),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_3009),
.B(n_2098),
.Y(n_3134)
);

AND2x6_ASAP7_75t_L g3135 ( 
.A(n_2969),
.B(n_2418),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_3080),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_3032),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2972),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2987),
.Y(n_3139)
);

INVx4_ASAP7_75t_L g3140 ( 
.A(n_3000),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2998),
.B(n_2679),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_3032),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_2981),
.B(n_3001),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2994),
.Y(n_3144)
);

NAND2x1p5_ASAP7_75t_L g3145 ( 
.A(n_2951),
.B(n_2680),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_3064),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3002),
.Y(n_3147)
);

AND2x6_ASAP7_75t_L g3148 ( 
.A(n_3112),
.B(n_2443),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_3008),
.B(n_2443),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_3015),
.B(n_2686),
.Y(n_3150)
);

AND2x4_ASAP7_75t_L g3151 ( 
.A(n_2936),
.B(n_2942),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3016),
.Y(n_3152)
);

OR2x2_ASAP7_75t_L g3153 ( 
.A(n_3030),
.B(n_2955),
.Y(n_3153)
);

INVxp33_ASAP7_75t_SL g3154 ( 
.A(n_2953),
.Y(n_3154)
);

AND2x2_ASAP7_75t_SL g3155 ( 
.A(n_2938),
.B(n_2406),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_3007),
.Y(n_3156)
);

BUFx3_ASAP7_75t_L g3157 ( 
.A(n_3069),
.Y(n_3157)
);

INVx2_ASAP7_75t_SL g3158 ( 
.A(n_3092),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3020),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3023),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3026),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3028),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2947),
.B(n_2446),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3041),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_3043),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_3053),
.B(n_1803),
.Y(n_3166)
);

NAND3xp33_ASAP7_75t_L g3167 ( 
.A(n_3054),
.B(n_2488),
.C(n_2487),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_3080),
.Y(n_3168)
);

OR2x6_ASAP7_75t_L g3169 ( 
.A(n_3060),
.B(n_1901),
.Y(n_3169)
);

BUFx8_ASAP7_75t_SL g3170 ( 
.A(n_3120),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2948),
.B(n_2446),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_3080),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_3071),
.B(n_1833),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_3048),
.Y(n_3174)
);

NAND2xp33_ASAP7_75t_L g3175 ( 
.A(n_3081),
.B(n_2449),
.Y(n_3175)
);

OAI22xp33_ASAP7_75t_SL g3176 ( 
.A1(n_3042),
.A2(n_2525),
.B1(n_2512),
.B2(n_1886),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3049),
.B(n_2449),
.Y(n_3177)
);

NAND3xp33_ASAP7_75t_L g3178 ( 
.A(n_3011),
.B(n_1682),
.C(n_1681),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3102),
.Y(n_3179)
);

OR2x6_ASAP7_75t_L g3180 ( 
.A(n_3062),
.B(n_2242),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_SL g3181 ( 
.A(n_3082),
.B(n_2449),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3036),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_3085),
.B(n_2468),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3039),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3055),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2964),
.B(n_2951),
.Y(n_3186)
);

NOR2xp33_ASAP7_75t_L g3187 ( 
.A(n_3065),
.B(n_1873),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_2937),
.Y(n_3188)
);

AND2x4_ASAP7_75t_L g3189 ( 
.A(n_2944),
.B(n_2690),
.Y(n_3189)
);

BUFx6f_ASAP7_75t_L g3190 ( 
.A(n_3074),
.Y(n_3190)
);

INVx4_ASAP7_75t_L g3191 ( 
.A(n_3072),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3114),
.B(n_2468),
.Y(n_3192)
);

CKINVDCx5p33_ASAP7_75t_R g3193 ( 
.A(n_2939),
.Y(n_3193)
);

INVx4_ASAP7_75t_L g3194 ( 
.A(n_3073),
.Y(n_3194)
);

OAI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_3034),
.A2(n_2055),
.B1(n_2078),
.B2(n_2041),
.Y(n_3195)
);

AND2x6_ASAP7_75t_L g3196 ( 
.A(n_2995),
.B(n_2468),
.Y(n_3196)
);

CKINVDCx5p33_ASAP7_75t_R g3197 ( 
.A(n_2941),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3086),
.B(n_2691),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_2943),
.Y(n_3199)
);

AND2x4_ASAP7_75t_L g3200 ( 
.A(n_2949),
.B(n_2692),
.Y(n_3200)
);

INVx5_ASAP7_75t_L g3201 ( 
.A(n_3006),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3088),
.Y(n_3202)
);

INVx2_ASAP7_75t_SL g3203 ( 
.A(n_3091),
.Y(n_3203)
);

INVx1_ASAP7_75t_SL g3204 ( 
.A(n_3076),
.Y(n_3204)
);

BUFx3_ASAP7_75t_L g3205 ( 
.A(n_3077),
.Y(n_3205)
);

NAND3xp33_ASAP7_75t_L g3206 ( 
.A(n_3019),
.B(n_1685),
.C(n_1683),
.Y(n_3206)
);

NAND2xp33_ASAP7_75t_L g3207 ( 
.A(n_3017),
.B(n_2521),
.Y(n_3207)
);

AND2x2_ASAP7_75t_SL g3208 ( 
.A(n_2974),
.B(n_2521),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3090),
.Y(n_3209)
);

BUFx6f_ASAP7_75t_L g3210 ( 
.A(n_3109),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2993),
.B(n_2113),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3096),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3114),
.B(n_2521),
.Y(n_3213)
);

AND2x4_ASAP7_75t_L g3214 ( 
.A(n_2957),
.B(n_2693),
.Y(n_3214)
);

INVx3_ASAP7_75t_L g3215 ( 
.A(n_2946),
.Y(n_3215)
);

NAND3xp33_ASAP7_75t_L g3216 ( 
.A(n_3003),
.B(n_1691),
.C(n_1687),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3087),
.B(n_1733),
.Y(n_3217)
);

BUFx3_ASAP7_75t_L g3218 ( 
.A(n_2954),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2993),
.B(n_2141),
.Y(n_3219)
);

CKINVDCx5p33_ASAP7_75t_R g3220 ( 
.A(n_2945),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_3116),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3089),
.B(n_1835),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3097),
.B(n_1851),
.Y(n_3223)
);

NOR2x1p5_ASAP7_75t_L g3224 ( 
.A(n_2982),
.B(n_1694),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3111),
.Y(n_3225)
);

NOR2xp33_ASAP7_75t_L g3226 ( 
.A(n_2952),
.B(n_2178),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_2970),
.B(n_2971),
.Y(n_3227)
);

OR2x2_ASAP7_75t_L g3228 ( 
.A(n_3067),
.B(n_2189),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3061),
.B(n_2694),
.Y(n_3229)
);

AND2x4_ASAP7_75t_L g3230 ( 
.A(n_2966),
.B(n_2700),
.Y(n_3230)
);

INVx4_ASAP7_75t_L g3231 ( 
.A(n_2990),
.Y(n_3231)
);

NAND2x1p5_ASAP7_75t_L g3232 ( 
.A(n_2967),
.B(n_2706),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_3113),
.B(n_2712),
.Y(n_3233)
);

CKINVDCx5p33_ASAP7_75t_R g3234 ( 
.A(n_2950),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3063),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3066),
.B(n_1946),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_3115),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3103),
.Y(n_3238)
);

BUFx2_ASAP7_75t_L g3239 ( 
.A(n_3005),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3078),
.Y(n_3240)
);

AND2x6_ASAP7_75t_L g3241 ( 
.A(n_3101),
.B(n_1689),
.Y(n_3241)
);

INVx2_ASAP7_75t_SL g3242 ( 
.A(n_3100),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3079),
.Y(n_3243)
);

INVx1_ASAP7_75t_SL g3244 ( 
.A(n_3098),
.Y(n_3244)
);

OR2x2_ASAP7_75t_L g3245 ( 
.A(n_3031),
.B(n_2387),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3083),
.Y(n_3246)
);

BUFx6f_ASAP7_75t_L g3247 ( 
.A(n_3109),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3110),
.B(n_2011),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_3104),
.B(n_2455),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3108),
.B(n_2029),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3105),
.Y(n_3251)
);

OR2x2_ASAP7_75t_L g3252 ( 
.A(n_2992),
.B(n_2457),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3106),
.B(n_3107),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3084),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2988),
.B(n_1696),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3024),
.B(n_1767),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3095),
.B(n_2940),
.Y(n_3257)
);

INVx3_ASAP7_75t_L g3258 ( 
.A(n_3068),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3035),
.A2(n_2379),
.B1(n_2089),
.B2(n_2094),
.Y(n_3259)
);

INVx4_ASAP7_75t_L g3260 ( 
.A(n_2991),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_3037),
.A2(n_2523),
.B1(n_2494),
.B2(n_1698),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3093),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3052),
.Y(n_3263)
);

BUFx6f_ASAP7_75t_L g3264 ( 
.A(n_3056),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_3044),
.B(n_1697),
.Y(n_3265)
);

INVx4_ASAP7_75t_L g3266 ( 
.A(n_2958),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_3057),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3027),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3059),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_SL g3270 ( 
.A(n_3046),
.B(n_3047),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_2999),
.B(n_1701),
.Y(n_3271)
);

INVx3_ASAP7_75t_L g3272 ( 
.A(n_2977),
.Y(n_3272)
);

BUFx10_ASAP7_75t_L g3273 ( 
.A(n_2965),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3099),
.B(n_2034),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3022),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_3038),
.B(n_1705),
.Y(n_3276)
);

AND2x6_ASAP7_75t_L g3277 ( 
.A(n_3040),
.B(n_1690),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_3025),
.B(n_2272),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3013),
.B(n_2292),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3010),
.B(n_2353),
.Y(n_3280)
);

AND2x4_ASAP7_75t_L g3281 ( 
.A(n_2973),
.B(n_2714),
.Y(n_3281)
);

INVx4_ASAP7_75t_L g3282 ( 
.A(n_2956),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_SL g3283 ( 
.A(n_3018),
.B(n_1711),
.Y(n_3283)
);

INVx4_ASAP7_75t_L g3284 ( 
.A(n_3117),
.Y(n_3284)
);

INVxp67_ASAP7_75t_L g3285 ( 
.A(n_2984),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3029),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_2986),
.B(n_1810),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3045),
.Y(n_3288)
);

AND2x6_ASAP7_75t_L g3289 ( 
.A(n_2959),
.B(n_1692),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3051),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3050),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_SL g3292 ( 
.A(n_3118),
.B(n_1714),
.Y(n_3292)
);

BUFx6f_ASAP7_75t_L g3293 ( 
.A(n_2979),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_3119),
.B(n_1715),
.Y(n_3294)
);

CKINVDCx5p33_ASAP7_75t_R g3295 ( 
.A(n_2960),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2989),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3021),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_2978),
.B(n_1810),
.Y(n_3298)
);

AND2x6_ASAP7_75t_L g3299 ( 
.A(n_3004),
.B(n_1695),
.Y(n_3299)
);

INVx4_ASAP7_75t_L g3300 ( 
.A(n_3014),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_2983),
.B(n_1720),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3012),
.Y(n_3302)
);

OR2x2_ASAP7_75t_L g3303 ( 
.A(n_2961),
.B(n_2456),
.Y(n_3303)
);

NOR2xp33_ASAP7_75t_L g3304 ( 
.A(n_2962),
.B(n_1722),
.Y(n_3304)
);

BUFx6f_ASAP7_75t_L g3305 ( 
.A(n_3058),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2947),
.B(n_1729),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_2980),
.B(n_2715),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_3081),
.A2(n_2084),
.B1(n_2119),
.B2(n_2072),
.Y(n_3308)
);

AND2x4_ASAP7_75t_L g3309 ( 
.A(n_2980),
.B(n_1700),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3094),
.Y(n_3310)
);

INVx6_ASAP7_75t_L g3311 ( 
.A(n_3080),
.Y(n_3311)
);

NAND2x1p5_ASAP7_75t_L g3312 ( 
.A(n_2997),
.B(n_1713),
.Y(n_3312)
);

BUFx6f_ASAP7_75t_L g3313 ( 
.A(n_3121),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3094),
.Y(n_3314)
);

OAI22xp5_ASAP7_75t_L g3315 ( 
.A1(n_3081),
.A2(n_1735),
.B1(n_1736),
.B2(n_1734),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3094),
.Y(n_3316)
);

NAND3xp33_ASAP7_75t_L g3317 ( 
.A(n_3033),
.B(n_1739),
.C(n_1737),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3094),
.Y(n_3318)
);

INVx3_ASAP7_75t_L g3319 ( 
.A(n_3121),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3094),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_3121),
.Y(n_3321)
);

BUFx6f_ASAP7_75t_L g3322 ( 
.A(n_3121),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3094),
.Y(n_3323)
);

AOI22xp33_ASAP7_75t_L g3324 ( 
.A1(n_3081),
.A2(n_2169),
.B1(n_2202),
.B2(n_2133),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3094),
.Y(n_3325)
);

BUFx3_ASAP7_75t_L g3326 ( 
.A(n_2980),
.Y(n_3326)
);

OAI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3081),
.A2(n_1741),
.B1(n_1743),
.B2(n_1740),
.Y(n_3327)
);

CKINVDCx20_ASAP7_75t_R g3328 ( 
.A(n_2954),
.Y(n_3328)
);

BUFx3_ASAP7_75t_L g3329 ( 
.A(n_2980),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3009),
.B(n_1744),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3094),
.Y(n_3331)
);

BUFx6f_ASAP7_75t_L g3332 ( 
.A(n_3121),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2947),
.B(n_1747),
.Y(n_3333)
);

AND2x4_ASAP7_75t_L g3334 ( 
.A(n_2980),
.B(n_1716),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_SL g3335 ( 
.A(n_2963),
.B(n_1890),
.Y(n_3335)
);

NOR2xp33_ASAP7_75t_L g3336 ( 
.A(n_3009),
.B(n_1750),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3094),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3094),
.Y(n_3338)
);

CKINVDCx5p33_ASAP7_75t_R g3339 ( 
.A(n_2937),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2947),
.B(n_1753),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3094),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3094),
.Y(n_3342)
);

BUFx10_ASAP7_75t_L g3343 ( 
.A(n_2963),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_SL g3344 ( 
.A(n_3033),
.B(n_1756),
.Y(n_3344)
);

NAND3x1_ASAP7_75t_L g3345 ( 
.A(n_2995),
.B(n_1726),
.C(n_1724),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3081),
.A2(n_1758),
.B1(n_1759),
.B2(n_1757),
.Y(n_3346)
);

HB1xp67_ASAP7_75t_L g3347 ( 
.A(n_2998),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3094),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_L g3349 ( 
.A(n_3009),
.B(n_1768),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3094),
.Y(n_3350)
);

INVx3_ASAP7_75t_L g3351 ( 
.A(n_3121),
.Y(n_3351)
);

AND2x4_ASAP7_75t_L g3352 ( 
.A(n_2980),
.B(n_1728),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_2975),
.Y(n_3353)
);

AND2x6_ASAP7_75t_L g3354 ( 
.A(n_2969),
.B(n_1732),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_3033),
.B(n_1770),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3094),
.Y(n_3356)
);

INVx1_ASAP7_75t_SL g3357 ( 
.A(n_3070),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_3009),
.B(n_1773),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_3081),
.A2(n_2258),
.B1(n_2283),
.B2(n_2222),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_R g3360 ( 
.A(n_3188),
.B(n_1894),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3238),
.B(n_1775),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3186),
.B(n_1776),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3122),
.B(n_1778),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3306),
.B(n_1779),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3138),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3125),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3127),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3143),
.B(n_1990),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3139),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3129),
.Y(n_3370)
);

AND2x4_ASAP7_75t_L g3371 ( 
.A(n_3157),
.B(n_1742),
.Y(n_3371)
);

AOI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3175),
.A2(n_1996),
.B1(n_2020),
.B2(n_1991),
.Y(n_3372)
);

A2O1A1Ixp33_ASAP7_75t_L g3373 ( 
.A1(n_3226),
.A2(n_1748),
.B(n_1752),
.C(n_1745),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3333),
.B(n_3340),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3241),
.A2(n_2030),
.B1(n_2058),
.B2(n_2021),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3308),
.A2(n_2079),
.B1(n_2083),
.B2(n_2075),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3144),
.Y(n_3377)
);

AND2x6_ASAP7_75t_SL g3378 ( 
.A(n_3304),
.B(n_1754),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3147),
.Y(n_3379)
);

NOR3xp33_ASAP7_75t_L g3380 ( 
.A(n_3134),
.B(n_3265),
.C(n_3173),
.Y(n_3380)
);

NOR2xp67_ASAP7_75t_L g3381 ( 
.A(n_3282),
.B(n_1784),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_3249),
.B(n_2087),
.Y(n_3382)
);

NAND2x1_ASAP7_75t_L g3383 ( 
.A(n_3190),
.B(n_2654),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3152),
.Y(n_3384)
);

HB1xp67_ASAP7_75t_L g3385 ( 
.A(n_3281),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3159),
.Y(n_3386)
);

OAI221xp5_ASAP7_75t_L g3387 ( 
.A1(n_3259),
.A2(n_1780),
.B1(n_1786),
.B2(n_1774),
.C(n_1772),
.Y(n_3387)
);

OAI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_3153),
.A2(n_2139),
.B1(n_2146),
.B2(n_2116),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_3211),
.B(n_2151),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_3219),
.B(n_2158),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3241),
.A2(n_2208),
.B1(n_2223),
.B2(n_2204),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3160),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3179),
.B(n_1792),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3150),
.B(n_1793),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3161),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3330),
.B(n_1794),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3198),
.B(n_2091),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3162),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3164),
.Y(n_3399)
);

INVx8_ASAP7_75t_L g3400 ( 
.A(n_3170),
.Y(n_3400)
);

NAND2xp33_ASAP7_75t_L g3401 ( 
.A(n_3277),
.B(n_3210),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3336),
.B(n_1795),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3349),
.B(n_1798),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3358),
.B(n_1799),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_SL g3405 ( 
.A(n_3242),
.B(n_2225),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3229),
.B(n_3248),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_3128),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3165),
.B(n_1800),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3353),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3174),
.B(n_1801),
.Y(n_3410)
);

INVx2_ASAP7_75t_SL g3411 ( 
.A(n_3307),
.Y(n_3411)
);

AOI22xp33_ASAP7_75t_L g3412 ( 
.A1(n_3324),
.A2(n_2257),
.B1(n_2312),
.B2(n_2228),
.Y(n_3412)
);

A2O1A1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_3359),
.A2(n_1796),
.B(n_1804),
.C(n_1787),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3204),
.B(n_2352),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3163),
.B(n_1806),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3156),
.Y(n_3416)
);

OR2x2_ASAP7_75t_L g3417 ( 
.A(n_3252),
.B(n_1808),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_3251),
.B(n_3244),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3254),
.B(n_1814),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3171),
.B(n_1815),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3278),
.A2(n_2410),
.B1(n_2423),
.B2(n_2394),
.Y(n_3421)
);

BUFx3_ASAP7_75t_L g3422 ( 
.A(n_3205),
.Y(n_3422)
);

A2O1A1Ixp33_ASAP7_75t_L g3423 ( 
.A1(n_3216),
.A2(n_1816),
.B(n_1829),
.C(n_1811),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3240),
.Y(n_3424)
);

BUFx3_ASAP7_75t_L g3425 ( 
.A(n_3326),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3217),
.B(n_1817),
.Y(n_3426)
);

BUFx8_ASAP7_75t_L g3427 ( 
.A(n_3305),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3243),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3246),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3222),
.B(n_1821),
.Y(n_3430)
);

AOI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_3279),
.A2(n_2472),
.B1(n_2486),
.B2(n_2465),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3223),
.B(n_1823),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_3128),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_3357),
.B(n_2493),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3141),
.B(n_1825),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3227),
.B(n_2500),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3250),
.B(n_1827),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_3187),
.B(n_2502),
.Y(n_3438)
);

AOI22x1_ASAP7_75t_L g3439 ( 
.A1(n_3262),
.A2(n_1830),
.B1(n_1834),
.B2(n_1828),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3182),
.B(n_3184),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3133),
.B(n_2091),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3185),
.B(n_1836),
.Y(n_3442)
);

INVx3_ASAP7_75t_L g3443 ( 
.A(n_3130),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3202),
.B(n_1837),
.Y(n_3444)
);

BUFx2_ASAP7_75t_L g3445 ( 
.A(n_3239),
.Y(n_3445)
);

INVx3_ASAP7_75t_L g3446 ( 
.A(n_3130),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_L g3447 ( 
.A(n_3154),
.B(n_2528),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_SL g3448 ( 
.A(n_3203),
.B(n_2534),
.Y(n_3448)
);

AO221x1_ASAP7_75t_L g3449 ( 
.A1(n_3195),
.A2(n_1849),
.B1(n_1858),
.B2(n_1841),
.C(n_1832),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3208),
.B(n_2540),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3209),
.Y(n_3451)
);

BUFx3_ASAP7_75t_L g3452 ( 
.A(n_3329),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3212),
.Y(n_3453)
);

OAI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3335),
.A2(n_1840),
.B1(n_1843),
.B2(n_1839),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3287),
.B(n_2152),
.Y(n_3455)
);

INVx2_ASAP7_75t_SL g3456 ( 
.A(n_3309),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3196),
.B(n_1844),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3235),
.Y(n_3458)
);

INVx2_ASAP7_75t_SL g3459 ( 
.A(n_3334),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3196),
.B(n_1846),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3225),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3137),
.Y(n_3462)
);

OR2x6_ASAP7_75t_L g3463 ( 
.A(n_3191),
.B(n_3194),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3142),
.B(n_1848),
.Y(n_3464)
);

AND2x6_ASAP7_75t_SL g3465 ( 
.A(n_3302),
.B(n_1868),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3146),
.B(n_1850),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_3294),
.B(n_3347),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3257),
.B(n_1856),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3276),
.B(n_1857),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3233),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3192),
.B(n_1859),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3215),
.Y(n_3472)
);

OAI22xp5_ASAP7_75t_L g3473 ( 
.A1(n_3310),
.A2(n_1860),
.B1(n_1864),
.B2(n_1862),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3213),
.B(n_1867),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3221),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3177),
.Y(n_3476)
);

BUFx3_ASAP7_75t_L g3477 ( 
.A(n_3247),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3189),
.Y(n_3478)
);

NOR2xp33_ASAP7_75t_L g3479 ( 
.A(n_3270),
.B(n_1875),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3298),
.B(n_2152),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3201),
.B(n_1876),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_SL g3482 ( 
.A(n_3201),
.B(n_1877),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3228),
.A2(n_2539),
.B1(n_2323),
.B2(n_1869),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3354),
.A2(n_3255),
.B1(n_3206),
.B2(n_3178),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3314),
.A2(n_1871),
.B1(n_1880),
.B2(n_1872),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_3285),
.B(n_1883),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3316),
.B(n_1884),
.Y(n_3487)
);

NOR2xp33_ASAP7_75t_L g3488 ( 
.A(n_3291),
.B(n_3271),
.Y(n_3488)
);

NAND2x1_ASAP7_75t_L g3489 ( 
.A(n_3318),
.B(n_1847),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_L g3490 ( 
.A1(n_3320),
.A2(n_1904),
.B1(n_1909),
.B2(n_1882),
.Y(n_3490)
);

AOI22xp5_ASAP7_75t_L g3491 ( 
.A1(n_3317),
.A2(n_1895),
.B1(n_1897),
.B2(n_1889),
.Y(n_3491)
);

NAND2xp33_ASAP7_75t_L g3492 ( 
.A(n_3247),
.B(n_3193),
.Y(n_3492)
);

OAI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_3323),
.A2(n_1900),
.B1(n_1903),
.B2(n_1899),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3325),
.B(n_1911),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3312),
.B(n_2154),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3331),
.B(n_1912),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3236),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3200),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_3158),
.B(n_1917),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3214),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3337),
.B(n_1921),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3344),
.B(n_1922),
.Y(n_3502)
);

OAI221xp5_ASAP7_75t_L g3503 ( 
.A1(n_3261),
.A2(n_1926),
.B1(n_1932),
.B2(n_1919),
.C(n_1915),
.Y(n_3503)
);

AND2x4_ASAP7_75t_SL g3504 ( 
.A(n_3140),
.B(n_3343),
.Y(n_3504)
);

AND2x4_ASAP7_75t_L g3505 ( 
.A(n_3126),
.B(n_1933),
.Y(n_3505)
);

BUFx3_ASAP7_75t_L g3506 ( 
.A(n_3328),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3231),
.B(n_1927),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3338),
.B(n_1929),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_SL g3509 ( 
.A1(n_3155),
.A2(n_1935),
.B1(n_1936),
.B2(n_1931),
.Y(n_3509)
);

NOR3xp33_ASAP7_75t_L g3510 ( 
.A(n_3301),
.B(n_1940),
.C(n_1939),
.Y(n_3510)
);

NOR2xp33_ASAP7_75t_L g3511 ( 
.A(n_3355),
.B(n_1942),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3272),
.B(n_2154),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_3313),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3341),
.B(n_1944),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3296),
.B(n_3315),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3327),
.B(n_1948),
.Y(n_3516)
);

INVx3_ASAP7_75t_L g3517 ( 
.A(n_3313),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_3346),
.B(n_1950),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3342),
.B(n_1953),
.Y(n_3519)
);

BUFx6f_ASAP7_75t_L g3520 ( 
.A(n_3321),
.Y(n_3520)
);

NOR2x1p5_ASAP7_75t_L g3521 ( 
.A(n_3266),
.B(n_1956),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3230),
.Y(n_3522)
);

OR2x2_ASAP7_75t_L g3523 ( 
.A(n_3297),
.B(n_3268),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_3292),
.B(n_1958),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3260),
.B(n_1960),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3256),
.B(n_2211),
.Y(n_3526)
);

NAND2xp33_ASAP7_75t_L g3527 ( 
.A(n_3197),
.B(n_1961),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3348),
.B(n_1964),
.Y(n_3528)
);

INVx2_ASAP7_75t_SL g3529 ( 
.A(n_3352),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3131),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3145),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3350),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3151),
.Y(n_3533)
);

AOI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_3167),
.A2(n_1966),
.B1(n_1968),
.B2(n_1965),
.Y(n_3534)
);

NAND3xp33_ASAP7_75t_L g3535 ( 
.A(n_3207),
.B(n_1971),
.C(n_1970),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3263),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3356),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3149),
.B(n_1973),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3135),
.B(n_1975),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3135),
.B(n_1976),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3124),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3319),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3351),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3293),
.B(n_3284),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3232),
.Y(n_3545)
);

AOI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3132),
.A2(n_1980),
.B1(n_1983),
.B2(n_1978),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3321),
.Y(n_3547)
);

OR2x6_ASAP7_75t_L g3548 ( 
.A(n_3264),
.B(n_1937),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_SL g3549 ( 
.A(n_3199),
.B(n_3220),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3280),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3148),
.B(n_3245),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3322),
.Y(n_3552)
);

INVxp67_ASAP7_75t_L g3553 ( 
.A(n_3303),
.Y(n_3553)
);

NOR2x1p5_ASAP7_75t_L g3554 ( 
.A(n_3295),
.B(n_3258),
.Y(n_3554)
);

INVx2_ASAP7_75t_SL g3555 ( 
.A(n_3311),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3148),
.B(n_1988),
.Y(n_3556)
);

HB1xp67_ASAP7_75t_L g3557 ( 
.A(n_3322),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_3234),
.B(n_3339),
.Y(n_3558)
);

INVx8_ASAP7_75t_L g3559 ( 
.A(n_3169),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3275),
.B(n_1992),
.Y(n_3560)
);

NOR2xp33_ASAP7_75t_L g3561 ( 
.A(n_3283),
.B(n_1993),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3286),
.B(n_1994),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3288),
.B(n_1995),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3332),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3181),
.B(n_1998),
.Y(n_3565)
);

O2A1O1Ixp33_ASAP7_75t_L g3566 ( 
.A1(n_3176),
.A2(n_1951),
.B(n_1954),
.C(n_1949),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_3290),
.B(n_2000),
.Y(n_3567)
);

AND2x6_ASAP7_75t_SL g3568 ( 
.A(n_3269),
.B(n_1955),
.Y(n_3568)
);

BUFx12f_ASAP7_75t_L g3569 ( 
.A(n_3273),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3183),
.B(n_2003),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3345),
.B(n_2008),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3267),
.B(n_2012),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_3274),
.B(n_2013),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3218),
.B(n_2018),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3237),
.B(n_2019),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3264),
.B(n_2022),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3136),
.B(n_1957),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3180),
.B(n_2024),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3136),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3168),
.B(n_2025),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3168),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3172),
.B(n_2027),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3299),
.B(n_2028),
.Y(n_3583)
);

BUFx6f_ASAP7_75t_L g3584 ( 
.A(n_3305),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3224),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3289),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3300),
.B(n_2037),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3138),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3125),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3125),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3238),
.B(n_2040),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3125),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_3125),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3238),
.B(n_2042),
.Y(n_3594)
);

BUFx5_ASAP7_75t_L g3595 ( 
.A(n_3123),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3238),
.B(n_2044),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3122),
.A2(n_1984),
.B(n_1979),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3125),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3238),
.B(n_2045),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_3253),
.B(n_2052),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3125),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3238),
.B(n_2054),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3238),
.B(n_2060),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3122),
.A2(n_1987),
.B(n_1985),
.Y(n_3604)
);

HB1xp67_ASAP7_75t_L g3605 ( 
.A(n_3281),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3138),
.Y(n_3606)
);

INVxp67_ASAP7_75t_SL g3607 ( 
.A(n_3122),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_SL g3608 ( 
.A(n_3253),
.B(n_2070),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3125),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3238),
.B(n_2076),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3125),
.Y(n_3611)
);

NOR3xp33_ASAP7_75t_L g3612 ( 
.A(n_3143),
.B(n_2085),
.C(n_2081),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3138),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_SL g3614 ( 
.A(n_3253),
.B(n_2088),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_SL g3615 ( 
.A(n_3253),
.B(n_2090),
.Y(n_3615)
);

NAND2xp33_ASAP7_75t_L g3616 ( 
.A(n_3241),
.B(n_2092),
.Y(n_3616)
);

INVx2_ASAP7_75t_SL g3617 ( 
.A(n_3281),
.Y(n_3617)
);

BUFx3_ASAP7_75t_L g3618 ( 
.A(n_3157),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3238),
.B(n_2093),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3238),
.B(n_2096),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3238),
.B(n_2097),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3238),
.B(n_2101),
.Y(n_3622)
);

OAI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3253),
.A2(n_2103),
.B1(n_2105),
.B2(n_2102),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3238),
.B(n_2106),
.Y(n_3624)
);

BUFx3_ASAP7_75t_L g3625 ( 
.A(n_3157),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3138),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3166),
.B(n_2241),
.Y(n_3627)
);

NOR3xp33_ASAP7_75t_L g3628 ( 
.A(n_3143),
.B(n_2110),
.C(n_2109),
.Y(n_3628)
);

OR2x2_ASAP7_75t_L g3629 ( 
.A(n_3252),
.B(n_2111),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3374),
.B(n_2114),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3406),
.B(n_2117),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3607),
.A2(n_2001),
.B(n_1999),
.Y(n_3632)
);

AO21x1_ASAP7_75t_L g3633 ( 
.A1(n_3396),
.A2(n_2006),
.B(n_2005),
.Y(n_3633)
);

AO21x1_ASAP7_75t_L g3634 ( 
.A1(n_3402),
.A2(n_2017),
.B(n_2009),
.Y(n_3634)
);

OAI21xp33_ASAP7_75t_L g3635 ( 
.A1(n_3382),
.A2(n_3390),
.B(n_3389),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3532),
.Y(n_3636)
);

BUFx12f_ASAP7_75t_L g3637 ( 
.A(n_3427),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3537),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3476),
.A2(n_2038),
.B(n_2031),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3515),
.B(n_2121),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3366),
.Y(n_3641)
);

AOI21xp33_ASAP7_75t_L g3642 ( 
.A1(n_3438),
.A2(n_2129),
.B(n_2122),
.Y(n_3642)
);

A2O1A1Ixp33_ASAP7_75t_L g3643 ( 
.A1(n_3516),
.A2(n_2046),
.B(n_2048),
.C(n_2047),
.Y(n_3643)
);

INVxp67_ASAP7_75t_L g3644 ( 
.A(n_3523),
.Y(n_3644)
);

O2A1O1Ixp5_ASAP7_75t_L g3645 ( 
.A1(n_3489),
.A2(n_2050),
.B(n_2053),
.C(n_2051),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3362),
.B(n_2130),
.Y(n_3646)
);

AO22x1_ASAP7_75t_L g3647 ( 
.A1(n_3436),
.A2(n_2136),
.B1(n_2137),
.B2(n_2134),
.Y(n_3647)
);

AOI21xp33_ASAP7_75t_L g3648 ( 
.A1(n_3518),
.A2(n_2140),
.B(n_2138),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3367),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3497),
.A2(n_2062),
.B(n_2061),
.Y(n_3650)
);

AOI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_3550),
.A2(n_2064),
.B(n_2063),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3403),
.B(n_2144),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3365),
.Y(n_3653)
);

OAI21xp33_ASAP7_75t_L g3654 ( 
.A1(n_3412),
.A2(n_2147),
.B(n_2145),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3404),
.B(n_2149),
.Y(n_3655)
);

AOI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_3440),
.A2(n_2068),
.B(n_2066),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3364),
.B(n_2150),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_L g3658 ( 
.A(n_3414),
.B(n_2163),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3370),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3369),
.Y(n_3660)
);

AO21x1_ASAP7_75t_L g3661 ( 
.A1(n_3561),
.A2(n_2074),
.B(n_2073),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3363),
.A2(n_3430),
.B(n_3426),
.Y(n_3662)
);

O2A1O1Ixp33_ASAP7_75t_L g3663 ( 
.A1(n_3503),
.A2(n_2077),
.B(n_2107),
.C(n_2086),
.Y(n_3663)
);

AOI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_3432),
.A2(n_2115),
.B(n_2108),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3377),
.Y(n_3665)
);

OAI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3487),
.A2(n_3496),
.B(n_3494),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3379),
.Y(n_3667)
);

OAI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3501),
.A2(n_2120),
.B(n_2118),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3384),
.B(n_2174),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3467),
.B(n_2177),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3386),
.B(n_2180),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3380),
.B(n_3488),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3392),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3468),
.A2(n_2127),
.B(n_2125),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3395),
.B(n_2183),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3398),
.B(n_2184),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3399),
.B(n_2185),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_3437),
.A2(n_2135),
.B(n_2132),
.Y(n_3678)
);

A2O1A1Ixp33_ASAP7_75t_L g3679 ( 
.A1(n_3469),
.A2(n_2142),
.B(n_2148),
.C(n_2143),
.Y(n_3679)
);

OAI22xp5_ASAP7_75t_L g3680 ( 
.A1(n_3588),
.A2(n_2188),
.B1(n_2191),
.B2(n_2186),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3420),
.A2(n_2159),
.B(n_2153),
.Y(n_3681)
);

A2O1A1Ixp33_ASAP7_75t_L g3682 ( 
.A1(n_3502),
.A2(n_3511),
.B(n_3524),
.C(n_3479),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3606),
.B(n_2192),
.Y(n_3683)
);

OAI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3508),
.A2(n_2164),
.B(n_2161),
.Y(n_3684)
);

OAI22xp5_ASAP7_75t_L g3685 ( 
.A1(n_3613),
.A2(n_2196),
.B1(n_2201),
.B2(n_2194),
.Y(n_3685)
);

NOR2xp33_ASAP7_75t_L g3686 ( 
.A(n_3368),
.B(n_3388),
.Y(n_3686)
);

O2A1O1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3373),
.A2(n_2165),
.B(n_2170),
.C(n_2167),
.Y(n_3687)
);

HB1xp67_ASAP7_75t_L g3688 ( 
.A(n_3385),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3471),
.A2(n_2172),
.B(n_2171),
.Y(n_3689)
);

INVx4_ASAP7_75t_L g3690 ( 
.A(n_3584),
.Y(n_3690)
);

AOI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_3474),
.A2(n_2179),
.B(n_2173),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3383),
.A2(n_2182),
.B(n_2181),
.Y(n_3692)
);

O2A1O1Ixp33_ASAP7_75t_L g3693 ( 
.A1(n_3423),
.A2(n_2195),
.B(n_2203),
.C(n_2198),
.Y(n_3693)
);

INVx3_ASAP7_75t_L g3694 ( 
.A(n_3477),
.Y(n_3694)
);

OAI21xp33_ASAP7_75t_SL g3695 ( 
.A1(n_3626),
.A2(n_3536),
.B(n_3428),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_3415),
.A2(n_2210),
.B(n_2209),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_3400),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3372),
.B(n_2213),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3514),
.A2(n_2216),
.B(n_2212),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_L g3700 ( 
.A(n_3447),
.B(n_2214),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3627),
.B(n_2218),
.Y(n_3701)
);

O2A1O1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_3623),
.A2(n_2219),
.B(n_2224),
.C(n_2221),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3361),
.B(n_3591),
.Y(n_3703)
);

AOI21x1_ASAP7_75t_L g3704 ( 
.A1(n_3519),
.A2(n_2230),
.B(n_2229),
.Y(n_3704)
);

BUFx6f_ASAP7_75t_L g3705 ( 
.A(n_3433),
.Y(n_3705)
);

AOI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3528),
.A2(n_2236),
.B(n_2234),
.Y(n_3706)
);

INVx2_ASAP7_75t_SL g3707 ( 
.A(n_3605),
.Y(n_3707)
);

HB1xp67_ASAP7_75t_L g3708 ( 
.A(n_3445),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3594),
.B(n_2231),
.Y(n_3709)
);

INVx4_ASAP7_75t_L g3710 ( 
.A(n_3584),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3596),
.B(n_2232),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3599),
.A2(n_2250),
.B(n_2243),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3602),
.A2(n_2253),
.B(n_2252),
.Y(n_3713)
);

INVx4_ASAP7_75t_L g3714 ( 
.A(n_3422),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3424),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3603),
.B(n_2237),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3610),
.A2(n_2260),
.B(n_2256),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3619),
.B(n_2238),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3429),
.A2(n_2244),
.B1(n_2254),
.B2(n_2251),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3620),
.A2(n_2269),
.B(n_2263),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3621),
.A2(n_2271),
.B(n_2270),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3622),
.B(n_2255),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3624),
.B(n_2259),
.Y(n_3723)
);

OAI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_3419),
.A2(n_2276),
.B(n_2273),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_L g3725 ( 
.A(n_3421),
.B(n_2261),
.Y(n_3725)
);

OAI21x1_ASAP7_75t_L g3726 ( 
.A1(n_3462),
.A2(n_2285),
.B(n_2279),
.Y(n_3726)
);

A2O1A1Ixp33_ASAP7_75t_L g3727 ( 
.A1(n_3567),
.A2(n_2295),
.B(n_2298),
.C(n_2293),
.Y(n_3727)
);

AOI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3394),
.A2(n_2303),
.B(n_2302),
.Y(n_3728)
);

O2A1O1Ixp33_ASAP7_75t_SL g3729 ( 
.A1(n_3413),
.A2(n_2307),
.B(n_2317),
.C(n_2309),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3464),
.A2(n_2324),
.B(n_2321),
.Y(n_3730)
);

AOI21x1_ASAP7_75t_L g3731 ( 
.A1(n_3458),
.A2(n_2327),
.B(n_2325),
.Y(n_3731)
);

OR2x6_ASAP7_75t_L g3732 ( 
.A(n_3400),
.B(n_2333),
.Y(n_3732)
);

O2A1O1Ixp33_ASAP7_75t_L g3733 ( 
.A1(n_3435),
.A2(n_2336),
.B(n_2342),
.C(n_2339),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3397),
.B(n_3480),
.Y(n_3734)
);

INVx3_ASAP7_75t_L g3735 ( 
.A(n_3618),
.Y(n_3735)
);

AND2x4_ASAP7_75t_L g3736 ( 
.A(n_3625),
.B(n_2343),
.Y(n_3736)
);

AND2x4_ASAP7_75t_L g3737 ( 
.A(n_3425),
.B(n_2347),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3451),
.B(n_2264),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_SL g3739 ( 
.A(n_3484),
.B(n_2265),
.Y(n_3739)
);

A2O1A1Ixp33_ASAP7_75t_L g3740 ( 
.A1(n_3573),
.A2(n_2356),
.B(n_2360),
.C(n_2349),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3453),
.B(n_2268),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_SL g3742 ( 
.A(n_3544),
.B(n_2275),
.Y(n_3742)
);

AOI22xp5_ASAP7_75t_L g3743 ( 
.A1(n_3612),
.A2(n_2280),
.B1(n_2284),
.B2(n_2281),
.Y(n_3743)
);

OAI321xp33_ASAP7_75t_L g3744 ( 
.A1(n_3376),
.A2(n_2378),
.A3(n_2373),
.B1(n_2386),
.B2(n_2383),
.C(n_2374),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_3472),
.B(n_3475),
.Y(n_3745)
);

AOI33xp33_ASAP7_75t_L g3746 ( 
.A1(n_3483),
.A2(n_2408),
.A3(n_2409),
.B1(n_2426),
.B2(n_2416),
.B3(n_2407),
.Y(n_3746)
);

INVx3_ASAP7_75t_L g3747 ( 
.A(n_3452),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3466),
.A2(n_2430),
.B(n_2429),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3461),
.Y(n_3749)
);

BUFx8_ASAP7_75t_L g3750 ( 
.A(n_3569),
.Y(n_3750)
);

OAI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3485),
.A2(n_2286),
.B1(n_2291),
.B2(n_2290),
.Y(n_3751)
);

O2A1O1Ixp33_ASAP7_75t_L g3752 ( 
.A1(n_3566),
.A2(n_3571),
.B(n_3393),
.C(n_3410),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_3450),
.B(n_2301),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3409),
.Y(n_3754)
);

NOR2x2_ASAP7_75t_L g3755 ( 
.A(n_3548),
.B(n_1972),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3416),
.A2(n_2439),
.B(n_2431),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3455),
.B(n_2397),
.Y(n_3757)
);

O2A1O1Ixp33_ASAP7_75t_L g3758 ( 
.A1(n_3408),
.A2(n_2442),
.B(n_2453),
.C(n_2452),
.Y(n_3758)
);

NOR2xp33_ASAP7_75t_SL g3759 ( 
.A(n_3504),
.B(n_2397),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3589),
.B(n_2305),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3590),
.A2(n_2474),
.B(n_2469),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_SL g3762 ( 
.A(n_3512),
.B(n_2306),
.Y(n_3762)
);

NOR2xp67_ASAP7_75t_SL g3763 ( 
.A(n_3549),
.B(n_2489),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3431),
.B(n_2314),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_SL g3765 ( 
.A(n_3531),
.B(n_2315),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3592),
.B(n_3593),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3598),
.B(n_2322),
.Y(n_3767)
);

AO21x1_ASAP7_75t_L g3768 ( 
.A1(n_3628),
.A2(n_2498),
.B(n_2496),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3601),
.B(n_2328),
.Y(n_3769)
);

AOI21xp33_ASAP7_75t_L g3770 ( 
.A1(n_3417),
.A2(n_2330),
.B(n_2329),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3609),
.A2(n_2506),
.B(n_2504),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3611),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_3434),
.B(n_2334),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3490),
.B(n_2335),
.Y(n_3774)
);

NOR2x1p5_ASAP7_75t_SL g3775 ( 
.A(n_3595),
.B(n_2510),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_L g3776 ( 
.A(n_3405),
.B(n_2337),
.Y(n_3776)
);

BUFx6f_ASAP7_75t_L g3777 ( 
.A(n_3513),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3595),
.B(n_2340),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_SL g3779 ( 
.A(n_3486),
.B(n_2341),
.Y(n_3779)
);

NOR2xp33_ASAP7_75t_L g3780 ( 
.A(n_3448),
.B(n_2345),
.Y(n_3780)
);

BUFx12f_ASAP7_75t_L g3781 ( 
.A(n_3463),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3572),
.A2(n_2543),
.B(n_2529),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3597),
.B(n_2348),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3604),
.B(n_2351),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3551),
.A2(n_2357),
.B(n_2354),
.Y(n_3785)
);

INVx3_ASAP7_75t_L g3786 ( 
.A(n_3520),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3530),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_L g3788 ( 
.A1(n_3444),
.A2(n_2361),
.B(n_2359),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3542),
.Y(n_3789)
);

AOI21xp5_ASAP7_75t_L g3790 ( 
.A1(n_3442),
.A2(n_2363),
.B(n_2362),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3526),
.B(n_2364),
.Y(n_3791)
);

BUFx6f_ASAP7_75t_L g3792 ( 
.A(n_3520),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3560),
.A2(n_2377),
.B(n_2369),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3629),
.B(n_2382),
.Y(n_3794)
);

NOR2xp67_ASAP7_75t_L g3795 ( 
.A(n_3535),
.B(n_2384),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3441),
.B(n_2388),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_3553),
.B(n_2390),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3541),
.Y(n_3798)
);

AOI21x1_ASAP7_75t_L g3799 ( 
.A1(n_3600),
.A2(n_361),
.B(n_360),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3543),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3547),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3552),
.Y(n_3802)
);

AOI22xp5_ASAP7_75t_L g3803 ( 
.A1(n_3608),
.A2(n_2392),
.B1(n_2395),
.B2(n_2391),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3564),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_L g3805 ( 
.A(n_3418),
.B(n_2399),
.Y(n_3805)
);

AO21x1_ASAP7_75t_L g3806 ( 
.A1(n_3614),
.A2(n_362),
.B(n_361),
.Y(n_3806)
);

CKINVDCx5p33_ASAP7_75t_R g3807 ( 
.A(n_3506),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3562),
.A2(n_2403),
.B(n_2400),
.Y(n_3808)
);

AOI21x1_ASAP7_75t_L g3809 ( 
.A1(n_3615),
.A2(n_363),
.B(n_362),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3495),
.B(n_2412),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3473),
.B(n_2413),
.Y(n_3811)
);

A2O1A1Ixp33_ASAP7_75t_L g3812 ( 
.A1(n_3538),
.A2(n_2415),
.B(n_2417),
.C(n_2414),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3360),
.B(n_3478),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3493),
.B(n_3381),
.Y(n_3814)
);

INVx4_ASAP7_75t_L g3815 ( 
.A(n_3463),
.Y(n_3815)
);

HB1xp67_ASAP7_75t_L g3816 ( 
.A(n_3617),
.Y(n_3816)
);

OAI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3563),
.A2(n_2427),
.B(n_2419),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_SL g3818 ( 
.A(n_3498),
.B(n_2428),
.Y(n_3818)
);

BUFx6f_ASAP7_75t_L g3819 ( 
.A(n_3407),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3505),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3533),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3411),
.A2(n_2433),
.B(n_2432),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3574),
.B(n_2434),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3579),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_3500),
.A2(n_2436),
.B(n_2435),
.Y(n_3825)
);

O2A1O1Ixp33_ASAP7_75t_L g3826 ( 
.A1(n_3387),
.A2(n_2440),
.B(n_2441),
.C(n_2437),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_SL g3827 ( 
.A(n_3522),
.B(n_2444),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_3575),
.B(n_2445),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3580),
.A2(n_2448),
.B(n_2447),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3510),
.B(n_2454),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3557),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3443),
.B(n_2460),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3446),
.B(n_2462),
.Y(n_3833)
);

BUFx6f_ASAP7_75t_L g3834 ( 
.A(n_3517),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_3558),
.B(n_2464),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3454),
.B(n_2466),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_SL g3837 ( 
.A(n_3456),
.B(n_2467),
.Y(n_3837)
);

AND2x2_ASAP7_75t_SL g3838 ( 
.A(n_3492),
.B(n_365),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3459),
.B(n_2470),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3470),
.Y(n_3840)
);

OAI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_3565),
.A2(n_2475),
.B(n_2471),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3581),
.Y(n_3842)
);

NOR3xp33_ASAP7_75t_L g3843 ( 
.A(n_3509),
.B(n_2478),
.C(n_2476),
.Y(n_3843)
);

NOR2xp67_ASAP7_75t_L g3844 ( 
.A(n_3587),
.B(n_2481),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3375),
.B(n_2482),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3449),
.B(n_2484),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3439),
.A2(n_2490),
.B1(n_2491),
.B2(n_2485),
.Y(n_3847)
);

AOI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_3582),
.A2(n_2495),
.B(n_2492),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3499),
.A2(n_2503),
.B(n_2497),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3391),
.B(n_2505),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3576),
.A2(n_2508),
.B(n_2507),
.Y(n_3851)
);

A2O1A1Ixp33_ASAP7_75t_L g3852 ( 
.A1(n_3570),
.A2(n_2513),
.B(n_2514),
.C(n_2511),
.Y(n_3852)
);

BUFx2_ASAP7_75t_SL g3853 ( 
.A(n_3555),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3401),
.A2(n_3529),
.B(n_3525),
.Y(n_3854)
);

A2O1A1Ixp33_ASAP7_75t_L g3855 ( 
.A1(n_3586),
.A2(n_2516),
.B(n_2517),
.C(n_2515),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3577),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3682),
.A2(n_3616),
.B(n_3507),
.Y(n_3857)
);

A2O1A1Ixp33_ASAP7_75t_L g3858 ( 
.A1(n_3635),
.A2(n_3583),
.B(n_3460),
.C(n_3457),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_R g3859 ( 
.A(n_3697),
.B(n_3527),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3703),
.B(n_3491),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3734),
.B(n_3371),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3662),
.A2(n_3545),
.B(n_3482),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3666),
.A2(n_3481),
.B(n_3585),
.Y(n_3863)
);

INVx3_ASAP7_75t_SL g3864 ( 
.A(n_3807),
.Y(n_3864)
);

BUFx12f_ASAP7_75t_L g3865 ( 
.A(n_3637),
.Y(n_3865)
);

O2A1O1Ixp33_ASAP7_75t_SL g3866 ( 
.A1(n_3855),
.A2(n_3540),
.B(n_3556),
.C(n_3539),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3653),
.Y(n_3867)
);

NOR2xp33_ASAP7_75t_R g3868 ( 
.A(n_3735),
.B(n_3559),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3660),
.Y(n_3869)
);

INVx5_ASAP7_75t_L g3870 ( 
.A(n_3705),
.Y(n_3870)
);

OAI22xp5_ASAP7_75t_L g3871 ( 
.A1(n_3686),
.A2(n_3554),
.B1(n_3578),
.B2(n_3534),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3665),
.Y(n_3872)
);

OR2x6_ASAP7_75t_L g3873 ( 
.A(n_3690),
.B(n_3521),
.Y(n_3873)
);

OAI22xp5_ASAP7_75t_SL g3874 ( 
.A1(n_3838),
.A2(n_3378),
.B1(n_3546),
.B2(n_3465),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_SL g3875 ( 
.A1(n_3828),
.A2(n_3568),
.B1(n_2519),
.B2(n_2520),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3752),
.A2(n_2522),
.B(n_2518),
.Y(n_3876)
);

INVx1_ASAP7_75t_SL g3877 ( 
.A(n_3831),
.Y(n_3877)
);

AOI21x1_ASAP7_75t_L g3878 ( 
.A1(n_3814),
.A2(n_366),
.B(n_365),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_SL g3879 ( 
.A(n_3644),
.B(n_2526),
.Y(n_3879)
);

NOR3xp33_ASAP7_75t_L g3880 ( 
.A(n_3658),
.B(n_2530),
.C(n_2527),
.Y(n_3880)
);

A2O1A1Ixp33_ASAP7_75t_L g3881 ( 
.A1(n_3724),
.A2(n_2535),
.B(n_2536),
.C(n_2533),
.Y(n_3881)
);

INVxp67_ASAP7_75t_L g3882 ( 
.A(n_3688),
.Y(n_3882)
);

BUFx6f_ASAP7_75t_L g3883 ( 
.A(n_3705),
.Y(n_3883)
);

NOR3xp33_ASAP7_75t_SL g3884 ( 
.A(n_3725),
.B(n_3813),
.C(n_3764),
.Y(n_3884)
);

O2A1O1Ixp5_ASAP7_75t_L g3885 ( 
.A1(n_3668),
.A2(n_3684),
.B(n_3661),
.C(n_3640),
.Y(n_3885)
);

AO32x1_ASAP7_75t_L g3886 ( 
.A1(n_3680),
.A2(n_2),
.A3(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_3886)
);

O2A1O1Ixp33_ASAP7_75t_L g3887 ( 
.A1(n_3648),
.A2(n_368),
.B(n_369),
.C(n_367),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3630),
.B(n_3631),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3667),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3700),
.A2(n_369),
.B1(n_370),
.B2(n_367),
.Y(n_3890)
);

NOR2xp33_ASAP7_75t_L g3891 ( 
.A(n_3823),
.B(n_370),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3705),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3707),
.B(n_3835),
.Y(n_3893)
);

HAxp5_ASAP7_75t_L g3894 ( 
.A(n_3755),
.B(n_3698),
.CON(n_3894),
.SN(n_3894)
);

NAND3xp33_ASAP7_75t_L g3895 ( 
.A(n_3642),
.B(n_3),
.C(n_4),
.Y(n_3895)
);

O2A1O1Ixp33_ASAP7_75t_L g3896 ( 
.A1(n_3643),
.A2(n_372),
.B(n_374),
.C(n_371),
.Y(n_3896)
);

CKINVDCx6p67_ASAP7_75t_R g3897 ( 
.A(n_3781),
.Y(n_3897)
);

A2O1A1Ixp33_ASAP7_75t_SL g3898 ( 
.A1(n_3763),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_3898)
);

OR2x4_ASAP7_75t_L g3899 ( 
.A(n_3753),
.B(n_3773),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3759),
.B(n_374),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3652),
.A2(n_376),
.B(n_375),
.Y(n_3901)
);

O2A1O1Ixp33_ASAP7_75t_L g3902 ( 
.A1(n_3770),
.A2(n_377),
.B(n_378),
.C(n_376),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_SL g3903 ( 
.A(n_3856),
.B(n_377),
.Y(n_3903)
);

AND2x4_ASAP7_75t_L g3904 ( 
.A(n_3747),
.B(n_379),
.Y(n_3904)
);

BUFx5_ASAP7_75t_L g3905 ( 
.A(n_3673),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3715),
.Y(n_3906)
);

A2O1A1Ixp33_ASAP7_75t_L g3907 ( 
.A1(n_3826),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_3907)
);

BUFx6f_ASAP7_75t_L g3908 ( 
.A(n_3777),
.Y(n_3908)
);

INVx2_ASAP7_75t_SL g3909 ( 
.A(n_3710),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3749),
.A2(n_380),
.B1(n_381),
.B2(n_379),
.Y(n_3910)
);

BUFx4f_ASAP7_75t_L g3911 ( 
.A(n_3777),
.Y(n_3911)
);

BUFx3_ASAP7_75t_L g3912 ( 
.A(n_3777),
.Y(n_3912)
);

NOR2xp33_ASAP7_75t_R g3913 ( 
.A(n_3694),
.B(n_381),
.Y(n_3913)
);

OAI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_3695),
.A2(n_8),
.B(n_9),
.Y(n_3914)
);

INVx2_ASAP7_75t_SL g3915 ( 
.A(n_3792),
.Y(n_3915)
);

BUFx12f_ASAP7_75t_L g3916 ( 
.A(n_3750),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3636),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3655),
.B(n_8),
.Y(n_3918)
);

NAND2x1p5_ASAP7_75t_L g3919 ( 
.A(n_3792),
.B(n_382),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3638),
.Y(n_3920)
);

AOI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3646),
.A2(n_385),
.B(n_384),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3657),
.B(n_9),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_L g3923 ( 
.A(n_3670),
.B(n_384),
.Y(n_3923)
);

BUFx2_ASAP7_75t_L g3924 ( 
.A(n_3792),
.Y(n_3924)
);

NOR2xp33_ASAP7_75t_L g3925 ( 
.A(n_3709),
.B(n_3711),
.Y(n_3925)
);

BUFx6f_ASAP7_75t_L g3926 ( 
.A(n_3819),
.Y(n_3926)
);

OAI22xp5_ASAP7_75t_L g3927 ( 
.A1(n_3778),
.A2(n_387),
.B1(n_388),
.B2(n_386),
.Y(n_3927)
);

A2O1A1Ixp33_ASAP7_75t_L g3928 ( 
.A1(n_3776),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_3928)
);

OAI21xp33_ASAP7_75t_L g3929 ( 
.A1(n_3845),
.A2(n_10),
.B(n_12),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3810),
.B(n_387),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3722),
.A2(n_390),
.B(n_389),
.Y(n_3931)
);

OAI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3716),
.A2(n_391),
.B1(n_392),
.B2(n_390),
.Y(n_3932)
);

AO21x1_ASAP7_75t_L g3933 ( 
.A1(n_3739),
.A2(n_3702),
.B(n_3846),
.Y(n_3933)
);

BUFx2_ASAP7_75t_L g3934 ( 
.A(n_3786),
.Y(n_3934)
);

O2A1O1Ixp33_ASAP7_75t_SL g3935 ( 
.A1(n_3836),
.A2(n_13),
.B(n_10),
.C(n_12),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3718),
.A2(n_392),
.B(n_391),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_SL g3937 ( 
.A(n_3796),
.B(n_393),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3723),
.A2(n_394),
.B(n_393),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3805),
.B(n_394),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3641),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3701),
.B(n_13),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3766),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3649),
.Y(n_3943)
);

INVx5_ASAP7_75t_L g3944 ( 
.A(n_3819),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3791),
.B(n_395),
.Y(n_3945)
);

HB1xp67_ASAP7_75t_L g3946 ( 
.A(n_3816),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3744),
.B(n_395),
.Y(n_3947)
);

CKINVDCx5p33_ASAP7_75t_R g3948 ( 
.A(n_3732),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3659),
.Y(n_3949)
);

AOI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3854),
.A2(n_397),
.B(n_396),
.Y(n_3950)
);

OAI22xp5_ASAP7_75t_L g3951 ( 
.A1(n_3772),
.A2(n_398),
.B1(n_399),
.B2(n_396),
.Y(n_3951)
);

HB1xp67_ASAP7_75t_L g3952 ( 
.A(n_3820),
.Y(n_3952)
);

O2A1O1Ixp33_ASAP7_75t_L g3953 ( 
.A1(n_3811),
.A2(n_401),
.B(n_402),
.C(n_399),
.Y(n_3953)
);

NAND2x1p5_ASAP7_75t_L g3954 ( 
.A(n_3815),
.B(n_401),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3762),
.A2(n_404),
.B(n_403),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_SL g3956 ( 
.A(n_3780),
.B(n_403),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3850),
.B(n_15),
.Y(n_3957)
);

OAI22x1_ASAP7_75t_L g3958 ( 
.A1(n_3765),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_3958)
);

NOR2xp33_ASAP7_75t_L g3959 ( 
.A(n_3779),
.B(n_405),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3757),
.B(n_406),
.Y(n_3960)
);

CKINVDCx5p33_ASAP7_75t_R g3961 ( 
.A(n_3819),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3840),
.B(n_406),
.Y(n_3962)
);

OAI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3787),
.A2(n_408),
.B1(n_409),
.B2(n_407),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3754),
.Y(n_3964)
);

O2A1O1Ixp33_ASAP7_75t_L g3965 ( 
.A1(n_3679),
.A2(n_409),
.B(n_410),
.C(n_407),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3844),
.B(n_15),
.Y(n_3966)
);

O2A1O1Ixp5_ASAP7_75t_L g3967 ( 
.A1(n_3633),
.A2(n_411),
.B(n_412),
.C(n_410),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3821),
.Y(n_3968)
);

CKINVDCx5p33_ASAP7_75t_R g3969 ( 
.A(n_3834),
.Y(n_3969)
);

OAI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3798),
.A2(n_3800),
.B1(n_3789),
.B2(n_3801),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3804),
.Y(n_3971)
);

AO21x1_ASAP7_75t_L g3972 ( 
.A1(n_3731),
.A2(n_415),
.B(n_413),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_SL g3973 ( 
.A(n_3797),
.B(n_3843),
.Y(n_3973)
);

BUFx2_ASAP7_75t_L g3974 ( 
.A(n_3834),
.Y(n_3974)
);

AO32x1_ASAP7_75t_L g3975 ( 
.A1(n_3685),
.A2(n_18),
.A3(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_3975)
);

O2A1O1Ixp5_ASAP7_75t_L g3976 ( 
.A1(n_3634),
.A2(n_416),
.B(n_417),
.C(n_415),
.Y(n_3976)
);

BUFx12f_ASAP7_75t_L g3977 ( 
.A(n_3834),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_SL g3978 ( 
.A(n_3736),
.B(n_16),
.Y(n_3978)
);

BUFx6f_ASAP7_75t_L g3979 ( 
.A(n_3737),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3746),
.B(n_17),
.Y(n_3980)
);

NAND3xp33_ASAP7_75t_L g3981 ( 
.A(n_3647),
.B(n_19),
.C(n_20),
.Y(n_3981)
);

BUFx6f_ASAP7_75t_L g3982 ( 
.A(n_3824),
.Y(n_3982)
);

NAND3xp33_ASAP7_75t_SL g3983 ( 
.A(n_3768),
.B(n_20),
.C(n_21),
.Y(n_3983)
);

OAI21x1_ASAP7_75t_L g3984 ( 
.A1(n_3726),
.A2(n_21),
.B(n_22),
.Y(n_3984)
);

OAI22xp5_ASAP7_75t_L g3985 ( 
.A1(n_3802),
.A2(n_419),
.B1(n_420),
.B2(n_418),
.Y(n_3985)
);

AOI21x1_ASAP7_75t_L g3986 ( 
.A1(n_3704),
.A2(n_420),
.B(n_419),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_3760),
.A2(n_422),
.B(n_421),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3767),
.A2(n_423),
.B(n_421),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3669),
.B(n_21),
.Y(n_3989)
);

BUFx2_ASAP7_75t_L g3990 ( 
.A(n_3842),
.Y(n_3990)
);

A2O1A1Ixp33_ASAP7_75t_L g3991 ( 
.A1(n_3733),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_L g3992 ( 
.A(n_3794),
.B(n_423),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3830),
.B(n_424),
.Y(n_3993)
);

OAI22xp5_ASAP7_75t_L g3994 ( 
.A1(n_3671),
.A2(n_426),
.B1(n_427),
.B2(n_425),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3675),
.B(n_22),
.Y(n_3995)
);

CKINVDCx20_ASAP7_75t_R g3996 ( 
.A(n_3742),
.Y(n_3996)
);

AOI21x1_ASAP7_75t_L g3997 ( 
.A1(n_3799),
.A2(n_426),
.B(n_425),
.Y(n_3997)
);

BUFx6f_ASAP7_75t_L g3998 ( 
.A(n_3809),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3745),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3743),
.B(n_428),
.Y(n_4000)
);

AOI21xp5_ASAP7_75t_L g4001 ( 
.A1(n_3769),
.A2(n_429),
.B(n_428),
.Y(n_4001)
);

O2A1O1Ixp33_ASAP7_75t_L g4002 ( 
.A1(n_3740),
.A2(n_430),
.B(n_432),
.C(n_429),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_L g4003 ( 
.A(n_3654),
.B(n_430),
.Y(n_4003)
);

O2A1O1Ixp33_ASAP7_75t_L g4004 ( 
.A1(n_3727),
.A2(n_3852),
.B(n_3812),
.C(n_3758),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3818),
.A2(n_433),
.B(n_432),
.Y(n_4005)
);

NOR2xp67_ASAP7_75t_L g4006 ( 
.A(n_3832),
.B(n_23),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3632),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_L g4008 ( 
.A(n_3676),
.B(n_23),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3827),
.A2(n_434),
.B(n_433),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3677),
.B(n_24),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_SL g4011 ( 
.A(n_3683),
.B(n_435),
.Y(n_4011)
);

AND2x2_ASAP7_75t_SL g4012 ( 
.A(n_3774),
.B(n_435),
.Y(n_4012)
);

BUFx3_ASAP7_75t_L g4013 ( 
.A(n_3833),
.Y(n_4013)
);

OAI22xp5_ASAP7_75t_L g4014 ( 
.A1(n_3738),
.A2(n_438),
.B1(n_439),
.B2(n_437),
.Y(n_4014)
);

A2O1A1Ixp33_ASAP7_75t_L g4015 ( 
.A1(n_3775),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_4015)
);

AND2x4_ASAP7_75t_L g4016 ( 
.A(n_3837),
.B(n_440),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_L g4017 ( 
.A(n_3741),
.B(n_440),
.Y(n_4017)
);

AND2x4_ASAP7_75t_L g4018 ( 
.A(n_3839),
.B(n_441),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_3825),
.A2(n_444),
.B(n_441),
.Y(n_4019)
);

OAI22xp5_ASAP7_75t_L g4020 ( 
.A1(n_3783),
.A2(n_445),
.B1(n_446),
.B2(n_444),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3645),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3784),
.A2(n_448),
.B(n_447),
.Y(n_4022)
);

NOR2x1_ASAP7_75t_L g4023 ( 
.A(n_3795),
.B(n_448),
.Y(n_4023)
);

INVx4_ASAP7_75t_L g4024 ( 
.A(n_3806),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3817),
.B(n_449),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_3674),
.A2(n_450),
.B(n_449),
.Y(n_4026)
);

INVx1_ASAP7_75t_SL g4027 ( 
.A(n_3692),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_3728),
.A2(n_452),
.B(n_450),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3719),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_R g4030 ( 
.A(n_3847),
.B(n_453),
.Y(n_4030)
);

NOR2x1_ASAP7_75t_L g4031 ( 
.A(n_3822),
.B(n_453),
.Y(n_4031)
);

O2A1O1Ixp33_ASAP7_75t_L g4032 ( 
.A1(n_3663),
.A2(n_455),
.B(n_456),
.C(n_454),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3639),
.Y(n_4033)
);

CKINVDCx8_ASAP7_75t_R g4034 ( 
.A(n_3785),
.Y(n_4034)
);

NOR2xp33_ASAP7_75t_L g4035 ( 
.A(n_3803),
.B(n_454),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3751),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3756),
.A2(n_3771),
.B(n_3761),
.Y(n_4037)
);

O2A1O1Ixp5_ASAP7_75t_SL g4038 ( 
.A1(n_3841),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_4038)
);

OAI22xp5_ASAP7_75t_L g4039 ( 
.A1(n_3788),
.A2(n_456),
.B1(n_457),
.B2(n_455),
.Y(n_4039)
);

A2O1A1Ixp33_ASAP7_75t_L g4040 ( 
.A1(n_3790),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_4040)
);

AOI21x1_ASAP7_75t_L g4041 ( 
.A1(n_3699),
.A2(n_459),
.B(n_458),
.Y(n_4041)
);

INVxp67_ASAP7_75t_SL g4042 ( 
.A(n_3650),
.Y(n_4042)
);

BUFx8_ASAP7_75t_L g4043 ( 
.A(n_3782),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3656),
.Y(n_4044)
);

INVx3_ASAP7_75t_L g4045 ( 
.A(n_3651),
.Y(n_4045)
);

A2O1A1Ixp33_ASAP7_75t_L g4046 ( 
.A1(n_3793),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_4046)
);

O2A1O1Ixp33_ASAP7_75t_L g4047 ( 
.A1(n_3706),
.A2(n_461),
.B(n_462),
.C(n_460),
.Y(n_4047)
);

INVx3_ASAP7_75t_SL g4048 ( 
.A(n_3712),
.Y(n_4048)
);

NAND2x2_ASAP7_75t_L g4049 ( 
.A(n_3851),
.B(n_29),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3713),
.B(n_29),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3717),
.A2(n_464),
.B(n_463),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3720),
.B(n_3721),
.Y(n_4052)
);

BUFx8_ASAP7_75t_L g4053 ( 
.A(n_3730),
.Y(n_4053)
);

OAI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3808),
.A2(n_3848),
.B(n_3829),
.Y(n_4054)
);

INVxp67_ASAP7_75t_SL g4055 ( 
.A(n_3687),
.Y(n_4055)
);

OAI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3748),
.A2(n_30),
.B(n_31),
.Y(n_4056)
);

BUFx6f_ASAP7_75t_L g4057 ( 
.A(n_3729),
.Y(n_4057)
);

AOI21xp5_ASAP7_75t_L g4058 ( 
.A1(n_3664),
.A2(n_464),
.B(n_463),
.Y(n_4058)
);

NOR3xp33_ASAP7_75t_SL g4059 ( 
.A(n_3849),
.B(n_32),
.C(n_33),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3681),
.B(n_3696),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_SL g4061 ( 
.A(n_3678),
.B(n_465),
.Y(n_4061)
);

NOR2xp33_ASAP7_75t_L g4062 ( 
.A(n_3689),
.B(n_3691),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3693),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3653),
.Y(n_4064)
);

OAI22xp5_ASAP7_75t_L g4065 ( 
.A1(n_3682),
.A2(n_469),
.B1(n_470),
.B2(n_466),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3635),
.B(n_32),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3635),
.B(n_33),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3653),
.Y(n_4068)
);

OR2x2_ASAP7_75t_L g4069 ( 
.A(n_3644),
.B(n_34),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3734),
.B(n_469),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3682),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_4071)
);

NOR2xp33_ASAP7_75t_SL g4072 ( 
.A(n_3714),
.B(n_34),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3635),
.B(n_35),
.Y(n_4073)
);

NOR2xp33_ASAP7_75t_L g4074 ( 
.A(n_3635),
.B(n_474),
.Y(n_4074)
);

INVx6_ASAP7_75t_L g4075 ( 
.A(n_3690),
.Y(n_4075)
);

CKINVDCx8_ASAP7_75t_R g4076 ( 
.A(n_3853),
.Y(n_4076)
);

HB1xp67_ASAP7_75t_L g4077 ( 
.A(n_3708),
.Y(n_4077)
);

O2A1O1Ixp5_ASAP7_75t_SL g4078 ( 
.A1(n_3672),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_4078)
);

AOI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_3682),
.A2(n_475),
.B(n_474),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_3637),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3653),
.Y(n_4081)
);

OAI21x1_ASAP7_75t_L g4082 ( 
.A1(n_3862),
.A2(n_36),
.B(n_37),
.Y(n_4082)
);

AO31x2_ASAP7_75t_L g4083 ( 
.A1(n_3933),
.A2(n_39),
.A3(n_36),
.B(n_38),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3925),
.B(n_39),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3872),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3889),
.Y(n_4086)
);

AO31x2_ASAP7_75t_L g4087 ( 
.A1(n_3972),
.A2(n_41),
.A3(n_39),
.B(n_40),
.Y(n_4087)
);

OA21x2_ASAP7_75t_L g4088 ( 
.A1(n_3914),
.A2(n_40),
.B(n_41),
.Y(n_4088)
);

INVx5_ASAP7_75t_L g4089 ( 
.A(n_3977),
.Y(n_4089)
);

A2O1A1Ixp33_ASAP7_75t_L g4090 ( 
.A1(n_3885),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4064),
.Y(n_4091)
);

OAI21x1_ASAP7_75t_L g4092 ( 
.A1(n_3984),
.A2(n_3857),
.B(n_4054),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_4077),
.B(n_477),
.Y(n_4093)
);

INVx3_ASAP7_75t_L g4094 ( 
.A(n_4076),
.Y(n_4094)
);

AO21x1_ASAP7_75t_L g4095 ( 
.A1(n_4025),
.A2(n_482),
.B(n_480),
.Y(n_4095)
);

CKINVDCx14_ASAP7_75t_R g4096 ( 
.A(n_3916),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3888),
.B(n_44),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3860),
.B(n_45),
.Y(n_4098)
);

INVx3_ASAP7_75t_L g4099 ( 
.A(n_4075),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_L g4100 ( 
.A(n_3899),
.B(n_483),
.Y(n_4100)
);

NOR2xp67_ASAP7_75t_L g4101 ( 
.A(n_3882),
.B(n_45),
.Y(n_4101)
);

A2O1A1Ixp33_ASAP7_75t_L g4102 ( 
.A1(n_3891),
.A2(n_4004),
.B(n_4062),
.C(n_3884),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3942),
.B(n_46),
.Y(n_4103)
);

OAI21x1_ASAP7_75t_SL g4104 ( 
.A1(n_4079),
.A2(n_47),
.B(n_48),
.Y(n_4104)
);

NOR2x1_ASAP7_75t_SL g4105 ( 
.A(n_3998),
.B(n_483),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_4060),
.A2(n_485),
.B(n_484),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_4070),
.B(n_48),
.Y(n_4107)
);

INVx3_ASAP7_75t_L g4108 ( 
.A(n_4075),
.Y(n_4108)
);

OA21x2_ASAP7_75t_L g4109 ( 
.A1(n_3950),
.A2(n_49),
.B(n_50),
.Y(n_4109)
);

INVx2_ASAP7_75t_SL g4110 ( 
.A(n_3944),
.Y(n_4110)
);

BUFx5_ASAP7_75t_L g4111 ( 
.A(n_3999),
.Y(n_4111)
);

BUFx6f_ASAP7_75t_L g4112 ( 
.A(n_3911),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3867),
.Y(n_4113)
);

OAI22x1_ASAP7_75t_L g4114 ( 
.A1(n_4074),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_4114)
);

AO31x2_ASAP7_75t_L g4115 ( 
.A1(n_4024),
.A2(n_53),
.A3(n_51),
.B(n_52),
.Y(n_4115)
);

AND2x6_ASAP7_75t_L g4116 ( 
.A(n_4033),
.B(n_4057),
.Y(n_4116)
);

BUFx6f_ASAP7_75t_L g4117 ( 
.A(n_3870),
.Y(n_4117)
);

A2O1A1Ixp33_ASAP7_75t_L g4118 ( 
.A1(n_3992),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_4118)
);

AOI22xp33_ASAP7_75t_L g4119 ( 
.A1(n_4035),
.A2(n_4003),
.B1(n_4000),
.B2(n_4030),
.Y(n_4119)
);

OA21x2_ASAP7_75t_L g4120 ( 
.A1(n_3863),
.A2(n_56),
.B(n_57),
.Y(n_4120)
);

BUFx10_ASAP7_75t_L g4121 ( 
.A(n_4080),
.Y(n_4121)
);

BUFx2_ASAP7_75t_L g4122 ( 
.A(n_3861),
.Y(n_4122)
);

CKINVDCx5p33_ASAP7_75t_R g4123 ( 
.A(n_3865),
.Y(n_4123)
);

OAI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3973),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_4124)
);

OAI21x1_ASAP7_75t_L g4125 ( 
.A1(n_4037),
.A2(n_60),
.B(n_61),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_4029),
.B(n_61),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_4052),
.A2(n_487),
.B(n_486),
.Y(n_4127)
);

NOR3xp33_ASAP7_75t_L g4128 ( 
.A(n_3874),
.B(n_61),
.C(n_62),
.Y(n_4128)
);

CKINVDCx12_ASAP7_75t_R g4129 ( 
.A(n_3873),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_3877),
.Y(n_4130)
);

AOI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_4042),
.A2(n_488),
.B(n_487),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3894),
.B(n_62),
.Y(n_4132)
);

OAI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_3893),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_4133)
);

OAI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_3858),
.A2(n_63),
.B(n_65),
.Y(n_4134)
);

AOI21xp5_ASAP7_75t_L g4135 ( 
.A1(n_3866),
.A2(n_491),
.B(n_490),
.Y(n_4135)
);

AO31x2_ASAP7_75t_L g4136 ( 
.A1(n_4021),
.A2(n_67),
.A3(n_65),
.B(n_66),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3869),
.Y(n_4137)
);

NAND3xp33_ASAP7_75t_SL g4138 ( 
.A(n_3880),
.B(n_66),
.C(n_67),
.Y(n_4138)
);

AO21x2_ASAP7_75t_L g4139 ( 
.A1(n_3876),
.A2(n_67),
.B(n_68),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_4017),
.B(n_68),
.Y(n_4140)
);

AOI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_4045),
.A2(n_491),
.B(n_490),
.Y(n_4141)
);

INVx5_ASAP7_75t_L g4142 ( 
.A(n_3883),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_4044),
.A2(n_493),
.B(n_492),
.Y(n_4143)
);

INVxp67_ASAP7_75t_L g4144 ( 
.A(n_3946),
.Y(n_4144)
);

BUFx2_ASAP7_75t_L g4145 ( 
.A(n_3924),
.Y(n_4145)
);

OAI22x1_ASAP7_75t_L g4146 ( 
.A1(n_3890),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_4146)
);

AOI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3959),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_L g4148 ( 
.A1(n_4007),
.A2(n_3871),
.B(n_4027),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_3917),
.Y(n_4149)
);

AO31x2_ASAP7_75t_L g4150 ( 
.A1(n_4065),
.A2(n_72),
.A3(n_70),
.B(n_71),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_4055),
.A2(n_494),
.B(n_493),
.Y(n_4151)
);

AO31x2_ASAP7_75t_L g4152 ( 
.A1(n_4071),
.A2(n_73),
.A3(n_71),
.B(n_72),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3918),
.B(n_74),
.Y(n_4153)
);

OAI21x1_ASAP7_75t_L g4154 ( 
.A1(n_3997),
.A2(n_4056),
.B(n_4041),
.Y(n_4154)
);

BUFx6f_ASAP7_75t_L g4155 ( 
.A(n_3870),
.Y(n_4155)
);

INVx6_ASAP7_75t_L g4156 ( 
.A(n_3944),
.Y(n_4156)
);

AOI21xp5_ASAP7_75t_L g4157 ( 
.A1(n_4063),
.A2(n_497),
.B(n_496),
.Y(n_4157)
);

AO31x2_ASAP7_75t_L g4158 ( 
.A1(n_4015),
.A2(n_77),
.A3(n_75),
.B(n_76),
.Y(n_4158)
);

AO31x2_ASAP7_75t_L g4159 ( 
.A1(n_3907),
.A2(n_78),
.A3(n_76),
.B(n_77),
.Y(n_4159)
);

OAI21x1_ASAP7_75t_SL g4160 ( 
.A1(n_3878),
.A2(n_78),
.B(n_79),
.Y(n_4160)
);

AOI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_4036),
.A2(n_497),
.B(n_496),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3922),
.A2(n_499),
.B(n_498),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_3945),
.B(n_79),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_4012),
.B(n_80),
.Y(n_4164)
);

AOI21x1_ASAP7_75t_SL g4165 ( 
.A1(n_3957),
.A2(n_80),
.B(n_81),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3906),
.Y(n_4166)
);

OAI21x1_ASAP7_75t_L g4167 ( 
.A1(n_3986),
.A2(n_81),
.B(n_82),
.Y(n_4167)
);

OAI21x1_ASAP7_75t_L g4168 ( 
.A1(n_3970),
.A2(n_83),
.B(n_84),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3940),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3990),
.B(n_83),
.Y(n_4170)
);

AOI221xp5_ASAP7_75t_L g4171 ( 
.A1(n_3929),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.C(n_87),
.Y(n_4171)
);

AOI22xp5_ASAP7_75t_L g4172 ( 
.A1(n_3923),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4068),
.Y(n_4173)
);

AOI31xp67_ASAP7_75t_L g4174 ( 
.A1(n_4061),
.A2(n_501),
.A3(n_502),
.B(n_500),
.Y(n_4174)
);

AOI21xp5_ASAP7_75t_SL g4175 ( 
.A1(n_4013),
.A2(n_503),
.B(n_502),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3989),
.B(n_88),
.Y(n_4176)
);

INVx5_ASAP7_75t_L g4177 ( 
.A(n_3883),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3995),
.B(n_89),
.Y(n_4178)
);

HB1xp67_ASAP7_75t_L g4179 ( 
.A(n_3952),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4008),
.B(n_90),
.Y(n_4180)
);

NOR2x1_ASAP7_75t_L g4181 ( 
.A(n_3895),
.B(n_504),
.Y(n_4181)
);

OAI22xp5_ASAP7_75t_L g4182 ( 
.A1(n_3996),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_4182)
);

O2A1O1Ixp33_ASAP7_75t_SL g4183 ( 
.A1(n_4040),
.A2(n_507),
.B(n_508),
.C(n_506),
.Y(n_4183)
);

AND2x6_ASAP7_75t_L g4184 ( 
.A(n_4057),
.B(n_508),
.Y(n_4184)
);

OAI21x1_ASAP7_75t_L g4185 ( 
.A1(n_4019),
.A2(n_92),
.B(n_93),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_4010),
.B(n_93),
.Y(n_4186)
);

OAI21x1_ASAP7_75t_L g4187 ( 
.A1(n_4038),
.A2(n_94),
.B(n_95),
.Y(n_4187)
);

OAI21x1_ASAP7_75t_L g4188 ( 
.A1(n_4078),
.A2(n_94),
.B(n_96),
.Y(n_4188)
);

AOI211x1_ASAP7_75t_L g4189 ( 
.A1(n_3939),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3943),
.Y(n_4190)
);

INVx2_ASAP7_75t_SL g4191 ( 
.A(n_3926),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3949),
.Y(n_4192)
);

INVx4_ASAP7_75t_L g4193 ( 
.A(n_3961),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_3947),
.A2(n_510),
.B(n_509),
.Y(n_4194)
);

NOR2x1_ASAP7_75t_L g4195 ( 
.A(n_3981),
.B(n_511),
.Y(n_4195)
);

INVx4_ASAP7_75t_L g4196 ( 
.A(n_3969),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_4066),
.B(n_100),
.Y(n_4197)
);

NAND2x1p5_ASAP7_75t_L g4198 ( 
.A(n_3974),
.B(n_3892),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_4067),
.B(n_102),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4073),
.B(n_103),
.Y(n_4200)
);

NAND3xp33_ASAP7_75t_SL g4201 ( 
.A(n_3875),
.B(n_103),
.C(n_104),
.Y(n_4201)
);

O2A1O1Ixp5_ASAP7_75t_L g4202 ( 
.A1(n_3956),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_4202)
);

OA21x2_ASAP7_75t_L g4203 ( 
.A1(n_3967),
.A2(n_105),
.B(n_106),
.Y(n_4203)
);

AND2x4_ASAP7_75t_L g4204 ( 
.A(n_3912),
.B(n_3934),
.Y(n_4204)
);

OAI21x1_ASAP7_75t_L g4205 ( 
.A1(n_3987),
.A2(n_4001),
.B(n_3988),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_3892),
.Y(n_4206)
);

AOI21x1_ASAP7_75t_SL g4207 ( 
.A1(n_3966),
.A2(n_3980),
.B(n_4050),
.Y(n_4207)
);

AO31x2_ASAP7_75t_L g4208 ( 
.A1(n_4046),
.A2(n_3928),
.A3(n_3991),
.B(n_4039),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3941),
.B(n_108),
.Y(n_4209)
);

AOI221x1_ASAP7_75t_L g4210 ( 
.A1(n_3983),
.A2(n_517),
.B1(n_518),
.B2(n_516),
.C(n_514),
.Y(n_4210)
);

OR2x6_ASAP7_75t_L g4211 ( 
.A(n_3873),
.B(n_517),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3920),
.B(n_109),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4081),
.Y(n_4213)
);

BUFx6f_ASAP7_75t_L g4214 ( 
.A(n_3908),
.Y(n_4214)
);

OAI21x1_ASAP7_75t_L g4215 ( 
.A1(n_3901),
.A2(n_109),
.B(n_110),
.Y(n_4215)
);

OAI21x1_ASAP7_75t_L g4216 ( 
.A1(n_3936),
.A2(n_111),
.B(n_112),
.Y(n_4216)
);

OAI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_3881),
.A2(n_111),
.B(n_112),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_SL g4218 ( 
.A(n_3905),
.B(n_518),
.Y(n_4218)
);

OA21x2_ASAP7_75t_L g4219 ( 
.A1(n_3976),
.A2(n_113),
.B(n_114),
.Y(n_4219)
);

AO31x2_ASAP7_75t_L g4220 ( 
.A1(n_3927),
.A2(n_4020),
.A3(n_3932),
.B(n_3958),
.Y(n_4220)
);

INVx1_ASAP7_75t_SL g4221 ( 
.A(n_3864),
.Y(n_4221)
);

OAI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4048),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_3909),
.B(n_521),
.Y(n_4223)
);

INVxp67_ASAP7_75t_SL g4224 ( 
.A(n_3968),
.Y(n_4224)
);

OA21x2_ASAP7_75t_L g4225 ( 
.A1(n_3931),
.A2(n_115),
.B(n_116),
.Y(n_4225)
);

OA21x2_ASAP7_75t_L g4226 ( 
.A1(n_3938),
.A2(n_117),
.B(n_118),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3971),
.Y(n_4227)
);

OAI21x1_ASAP7_75t_L g4228 ( 
.A1(n_3921),
.A2(n_4031),
.B(n_4022),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3964),
.Y(n_4229)
);

AOI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_4028),
.A2(n_523),
.B(n_522),
.Y(n_4230)
);

CKINVDCx14_ASAP7_75t_R g4231 ( 
.A(n_3859),
.Y(n_4231)
);

AOI21xp5_ASAP7_75t_L g4232 ( 
.A1(n_4026),
.A2(n_524),
.B(n_523),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3905),
.Y(n_4233)
);

INVx3_ASAP7_75t_SL g4234 ( 
.A(n_3897),
.Y(n_4234)
);

OA21x2_ASAP7_75t_L g4235 ( 
.A1(n_4005),
.A2(n_118),
.B(n_119),
.Y(n_4235)
);

BUFx6f_ASAP7_75t_L g4236 ( 
.A(n_3979),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3930),
.B(n_119),
.Y(n_4237)
);

OAI21x1_ASAP7_75t_L g4238 ( 
.A1(n_4058),
.A2(n_121),
.B(n_122),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_SL g4239 ( 
.A(n_3905),
.B(n_524),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4059),
.B(n_121),
.Y(n_4240)
);

AOI21xp5_ASAP7_75t_SL g4241 ( 
.A1(n_3896),
.A2(n_527),
.B(n_525),
.Y(n_4241)
);

BUFx6f_ASAP7_75t_L g4242 ( 
.A(n_3979),
.Y(n_4242)
);

INVxp67_ASAP7_75t_SL g4243 ( 
.A(n_3982),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3905),
.B(n_4072),
.Y(n_4244)
);

OAI21x1_ASAP7_75t_L g4245 ( 
.A1(n_4051),
.A2(n_122),
.B(n_123),
.Y(n_4245)
);

AOI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_3887),
.A2(n_527),
.B(n_525),
.Y(n_4246)
);

BUFx10_ASAP7_75t_L g4247 ( 
.A(n_3904),
.Y(n_4247)
);

OAI21x1_ASAP7_75t_L g4248 ( 
.A1(n_4009),
.A2(n_123),
.B(n_124),
.Y(n_4248)
);

OA21x2_ASAP7_75t_L g4249 ( 
.A1(n_3955),
.A2(n_124),
.B(n_125),
.Y(n_4249)
);

OA21x2_ASAP7_75t_L g4250 ( 
.A1(n_4011),
.A2(n_124),
.B(n_125),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3982),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4224),
.Y(n_4252)
);

OAI21x1_ASAP7_75t_L g4253 ( 
.A1(n_4092),
.A2(n_3965),
.B(n_3902),
.Y(n_4253)
);

OAI21x1_ASAP7_75t_L g4254 ( 
.A1(n_4154),
.A2(n_4002),
.B(n_3953),
.Y(n_4254)
);

OAI22xp33_ASAP7_75t_L g4255 ( 
.A1(n_4147),
.A2(n_4172),
.B1(n_4201),
.B2(n_4140),
.Y(n_4255)
);

INVx5_ASAP7_75t_SL g4256 ( 
.A(n_4112),
.Y(n_4256)
);

BUFx3_ASAP7_75t_L g4257 ( 
.A(n_4206),
.Y(n_4257)
);

BUFx3_ASAP7_75t_L g4258 ( 
.A(n_4099),
.Y(n_4258)
);

OAI21x1_ASAP7_75t_L g4259 ( 
.A1(n_4125),
.A2(n_4047),
.B(n_4032),
.Y(n_4259)
);

AOI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_4119),
.A2(n_4049),
.B1(n_3993),
.B2(n_4023),
.Y(n_4260)
);

BUFx3_ASAP7_75t_L g4261 ( 
.A(n_4108),
.Y(n_4261)
);

OAI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_4102),
.A2(n_3900),
.B1(n_3937),
.B2(n_4006),
.Y(n_4262)
);

INVx1_ASAP7_75t_SL g4263 ( 
.A(n_4122),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4098),
.B(n_3962),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4113),
.Y(n_4265)
);

OA21x2_ASAP7_75t_L g4266 ( 
.A1(n_4135),
.A2(n_3903),
.B(n_3960),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4130),
.B(n_4016),
.Y(n_4267)
);

OAI21x1_ASAP7_75t_L g4268 ( 
.A1(n_4082),
.A2(n_3985),
.B(n_3994),
.Y(n_4268)
);

OAI22xp5_ASAP7_75t_L g4269 ( 
.A1(n_4084),
.A2(n_4034),
.B1(n_3954),
.B2(n_4018),
.Y(n_4269)
);

OAI211xp5_ASAP7_75t_SL g4270 ( 
.A1(n_4128),
.A2(n_3879),
.B(n_4069),
.C(n_4014),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4137),
.Y(n_4271)
);

AO32x2_ASAP7_75t_L g4272 ( 
.A1(n_4222),
.A2(n_3910),
.A3(n_3963),
.B1(n_3951),
.B2(n_3886),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4166),
.Y(n_4273)
);

OAI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_4134),
.A2(n_4148),
.B(n_4217),
.Y(n_4274)
);

OAI21x1_ASAP7_75t_L g4275 ( 
.A1(n_4205),
.A2(n_3919),
.B(n_3886),
.Y(n_4275)
);

OA21x2_ASAP7_75t_L g4276 ( 
.A1(n_4228),
.A2(n_3898),
.B(n_3975),
.Y(n_4276)
);

NOR2xp33_ASAP7_75t_L g4277 ( 
.A(n_4221),
.B(n_3978),
.Y(n_4277)
);

OAI21x1_ASAP7_75t_L g4278 ( 
.A1(n_4167),
.A2(n_3975),
.B(n_3935),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4173),
.Y(n_4279)
);

OAI21x1_ASAP7_75t_L g4280 ( 
.A1(n_4185),
.A2(n_4207),
.B(n_4238),
.Y(n_4280)
);

OA21x2_ASAP7_75t_L g4281 ( 
.A1(n_4090),
.A2(n_3915),
.B(n_3948),
.Y(n_4281)
);

NAND2x1p5_ASAP7_75t_L g4282 ( 
.A(n_4089),
.B(n_4142),
.Y(n_4282)
);

OA21x2_ASAP7_75t_L g4283 ( 
.A1(n_4168),
.A2(n_4043),
.B(n_4053),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4132),
.B(n_3913),
.Y(n_4284)
);

OAI21x1_ASAP7_75t_L g4285 ( 
.A1(n_4245),
.A2(n_3868),
.B(n_126),
.Y(n_4285)
);

BUFx2_ASAP7_75t_L g4286 ( 
.A(n_4145),
.Y(n_4286)
);

BUFx6f_ASAP7_75t_L g4287 ( 
.A(n_4112),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4149),
.Y(n_4288)
);

BUFx2_ASAP7_75t_L g4289 ( 
.A(n_4204),
.Y(n_4289)
);

AOI22xp33_ASAP7_75t_L g4290 ( 
.A1(n_4138),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_4179),
.B(n_528),
.Y(n_4291)
);

AO21x2_ASAP7_75t_L g4292 ( 
.A1(n_4160),
.A2(n_128),
.B(n_130),
.Y(n_4292)
);

BUFx2_ASAP7_75t_L g4293 ( 
.A(n_4198),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4213),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_4231),
.Y(n_4295)
);

BUFx2_ASAP7_75t_L g4296 ( 
.A(n_4243),
.Y(n_4296)
);

OAI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_4246),
.A2(n_130),
.B(n_131),
.Y(n_4297)
);

CKINVDCx5p33_ASAP7_75t_R g4298 ( 
.A(n_4096),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4227),
.Y(n_4299)
);

NOR2xp67_ASAP7_75t_L g4300 ( 
.A(n_4094),
.B(n_4144),
.Y(n_4300)
);

OAI21x1_ASAP7_75t_L g4301 ( 
.A1(n_4233),
.A2(n_130),
.B(n_131),
.Y(n_4301)
);

INVx2_ASAP7_75t_SL g4302 ( 
.A(n_4156),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_4117),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4169),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4240),
.B(n_529),
.Y(n_4305)
);

AOI22xp33_ASAP7_75t_L g4306 ( 
.A1(n_4171),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_4306)
);

BUFx3_ASAP7_75t_L g4307 ( 
.A(n_4155),
.Y(n_4307)
);

BUFx6f_ASAP7_75t_L g4308 ( 
.A(n_4155),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4229),
.Y(n_4309)
);

OR2x2_ASAP7_75t_L g4310 ( 
.A(n_4085),
.B(n_530),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4097),
.B(n_530),
.Y(n_4311)
);

AOI21xp5_ASAP7_75t_L g4312 ( 
.A1(n_4244),
.A2(n_533),
.B(n_531),
.Y(n_4312)
);

OAI21xp5_ASAP7_75t_L g4313 ( 
.A1(n_4106),
.A2(n_135),
.B(n_136),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4181),
.B(n_531),
.Y(n_4314)
);

OAI22xp33_ASAP7_75t_L g4315 ( 
.A1(n_4211),
.A2(n_4210),
.B1(n_4146),
.B2(n_4182),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4107),
.B(n_534),
.Y(n_4316)
);

INVxp67_ASAP7_75t_L g4317 ( 
.A(n_4251),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4086),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4164),
.B(n_534),
.Y(n_4319)
);

OAI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4127),
.A2(n_139),
.B(n_140),
.Y(n_4320)
);

OAI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_4230),
.A2(n_141),
.B(n_142),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4190),
.Y(n_4322)
);

AO31x2_ASAP7_75t_L g4323 ( 
.A1(n_4095),
.A2(n_4232),
.A3(n_4143),
.B(n_4141),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4091),
.Y(n_4324)
);

OAI21x1_ASAP7_75t_L g4325 ( 
.A1(n_4215),
.A2(n_143),
.B(n_144),
.Y(n_4325)
);

INVx1_ASAP7_75t_SL g4326 ( 
.A(n_4247),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4194),
.A2(n_143),
.B(n_144),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4192),
.Y(n_4328)
);

AO21x2_ASAP7_75t_L g4329 ( 
.A1(n_4104),
.A2(n_145),
.B(n_146),
.Y(n_4329)
);

OAI21x1_ASAP7_75t_L g4330 ( 
.A1(n_4216),
.A2(n_145),
.B(n_146),
.Y(n_4330)
);

AOI21x1_ASAP7_75t_L g4331 ( 
.A1(n_4218),
.A2(n_147),
.B(n_148),
.Y(n_4331)
);

BUFx6f_ASAP7_75t_L g4332 ( 
.A(n_4214),
.Y(n_4332)
);

AO31x2_ASAP7_75t_L g4333 ( 
.A1(n_4105),
.A2(n_150),
.A3(n_148),
.B(n_149),
.Y(n_4333)
);

OAI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4211),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4334)
);

AOI22xp33_ASAP7_75t_L g4335 ( 
.A1(n_4195),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_4335)
);

OAI21x1_ASAP7_75t_L g4336 ( 
.A1(n_4248),
.A2(n_151),
.B(n_152),
.Y(n_4336)
);

OAI221xp5_ASAP7_75t_L g4337 ( 
.A1(n_4118),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_4337)
);

INVx4_ASAP7_75t_SL g4338 ( 
.A(n_4184),
.Y(n_4338)
);

INVx3_ASAP7_75t_L g4339 ( 
.A(n_4193),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4241),
.A2(n_536),
.B(n_535),
.Y(n_4340)
);

OAI21x1_ASAP7_75t_L g4341 ( 
.A1(n_4120),
.A2(n_155),
.B(n_156),
.Y(n_4341)
);

OAI21x1_ASAP7_75t_L g4342 ( 
.A1(n_4131),
.A2(n_155),
.B(n_156),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4126),
.B(n_535),
.Y(n_4343)
);

AO21x2_ASAP7_75t_L g4344 ( 
.A1(n_4239),
.A2(n_155),
.B(n_156),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4111),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_4197),
.B(n_536),
.Y(n_4346)
);

OR2x2_ASAP7_75t_L g4347 ( 
.A(n_4199),
.B(n_537),
.Y(n_4347)
);

OAI21xp5_ASAP7_75t_L g4348 ( 
.A1(n_4151),
.A2(n_157),
.B(n_158),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4136),
.Y(n_4349)
);

AND2x4_ASAP7_75t_L g4350 ( 
.A(n_4089),
.B(n_538),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4111),
.Y(n_4351)
);

OAI21x1_ASAP7_75t_L g4352 ( 
.A1(n_4165),
.A2(n_157),
.B(n_158),
.Y(n_4352)
);

NOR2xp67_ASAP7_75t_L g4353 ( 
.A(n_4196),
.B(n_159),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4163),
.B(n_4250),
.Y(n_4354)
);

INVx2_ASAP7_75t_SL g4355 ( 
.A(n_4142),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4136),
.Y(n_4356)
);

OA21x2_ASAP7_75t_L g4357 ( 
.A1(n_4187),
.A2(n_159),
.B(n_160),
.Y(n_4357)
);

AOI21xp33_ASAP7_75t_SL g4358 ( 
.A1(n_4100),
.A2(n_160),
.B(n_161),
.Y(n_4358)
);

OA21x2_ASAP7_75t_L g4359 ( 
.A1(n_4161),
.A2(n_160),
.B(n_162),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_4200),
.B(n_538),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4083),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4111),
.Y(n_4362)
);

CKINVDCx5p33_ASAP7_75t_R g4363 ( 
.A(n_4123),
.Y(n_4363)
);

A2O1A1Ixp33_ASAP7_75t_L g4364 ( 
.A1(n_4162),
.A2(n_540),
.B(n_541),
.C(n_539),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4235),
.Y(n_4365)
);

BUFx3_ASAP7_75t_L g4366 ( 
.A(n_4236),
.Y(n_4366)
);

OAI21x1_ASAP7_75t_L g4367 ( 
.A1(n_4109),
.A2(n_162),
.B(n_163),
.Y(n_4367)
);

OAI21xp5_ASAP7_75t_L g4368 ( 
.A1(n_4157),
.A2(n_164),
.B(n_165),
.Y(n_4368)
);

HB1xp67_ASAP7_75t_SL g4369 ( 
.A(n_4214),
.Y(n_4369)
);

AND2x4_ASAP7_75t_L g4370 ( 
.A(n_4177),
.B(n_541),
.Y(n_4370)
);

OAI21x1_ASAP7_75t_L g4371 ( 
.A1(n_4226),
.A2(n_168),
.B(n_169),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4083),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4225),
.Y(n_4373)
);

OAI21x1_ASAP7_75t_L g4374 ( 
.A1(n_4253),
.A2(n_4249),
.B(n_4219),
.Y(n_4374)
);

INVx5_ASAP7_75t_L g4375 ( 
.A(n_4303),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4265),
.Y(n_4376)
);

AO31x2_ASAP7_75t_L g4377 ( 
.A1(n_4361),
.A2(n_4114),
.A3(n_4124),
.B(n_4133),
.Y(n_4377)
);

AND2x4_ASAP7_75t_L g4378 ( 
.A(n_4286),
.B(n_4177),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4271),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4273),
.Y(n_4380)
);

INVx1_ASAP7_75t_SL g4381 ( 
.A(n_4289),
.Y(n_4381)
);

BUFx6f_ASAP7_75t_L g4382 ( 
.A(n_4287),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4279),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4318),
.Y(n_4384)
);

AOI21xp5_ASAP7_75t_L g4385 ( 
.A1(n_4274),
.A2(n_4088),
.B(n_4183),
.Y(n_4385)
);

OAI21x1_ASAP7_75t_L g4386 ( 
.A1(n_4280),
.A2(n_4203),
.B(n_4188),
.Y(n_4386)
);

AOI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_4313),
.A2(n_4139),
.B(n_4175),
.Y(n_4387)
);

BUFx12f_ASAP7_75t_L g4388 ( 
.A(n_4298),
.Y(n_4388)
);

OAI221xp5_ASAP7_75t_L g4389 ( 
.A1(n_4260),
.A2(n_4176),
.B1(n_4186),
.B2(n_4180),
.C(n_4178),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_4252),
.B(n_4153),
.Y(n_4390)
);

OA21x2_ASAP7_75t_L g4391 ( 
.A1(n_4341),
.A2(n_4202),
.B(n_4209),
.Y(n_4391)
);

OR2x2_ASAP7_75t_L g4392 ( 
.A(n_4294),
.B(n_4093),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4299),
.Y(n_4393)
);

OA21x2_ASAP7_75t_L g4394 ( 
.A1(n_4275),
.A2(n_4103),
.B(n_4212),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4309),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_4320),
.A2(n_4116),
.B(n_4237),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4349),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4356),
.Y(n_4398)
);

HB1xp67_ASAP7_75t_L g4399 ( 
.A(n_4296),
.Y(n_4399)
);

A2O1A1Ixp33_ASAP7_75t_L g4400 ( 
.A1(n_4340),
.A2(n_4101),
.B(n_4110),
.C(n_4170),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4324),
.Y(n_4401)
);

AND2x4_ASAP7_75t_SL g4402 ( 
.A(n_4339),
.B(n_4121),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4263),
.B(n_4223),
.Y(n_4403)
);

OAI21x1_ASAP7_75t_L g4404 ( 
.A1(n_4254),
.A2(n_4116),
.B(n_4174),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4372),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4288),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4304),
.Y(n_4407)
);

AO21x2_ASAP7_75t_L g4408 ( 
.A1(n_4321),
.A2(n_4087),
.B(n_4115),
.Y(n_4408)
);

OAI21x1_ASAP7_75t_L g4409 ( 
.A1(n_4259),
.A2(n_4115),
.B(n_4158),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_4322),
.Y(n_4410)
);

AOI21x1_ASAP7_75t_L g4411 ( 
.A1(n_4331),
.A2(n_4191),
.B(n_4158),
.Y(n_4411)
);

OAI21x1_ASAP7_75t_L g4412 ( 
.A1(n_4268),
.A2(n_4208),
.B(n_4159),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4354),
.B(n_4159),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_SL g4414 ( 
.A1(n_4297),
.A2(n_4184),
.B1(n_4220),
.B2(n_4150),
.Y(n_4414)
);

AO21x2_ASAP7_75t_L g4415 ( 
.A1(n_4348),
.A2(n_4152),
.B(n_4150),
.Y(n_4415)
);

HB1xp67_ASAP7_75t_L g4416 ( 
.A(n_4365),
.Y(n_4416)
);

NAND2x1p5_ASAP7_75t_L g4417 ( 
.A(n_4293),
.B(n_4242),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4305),
.B(n_4152),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4328),
.Y(n_4419)
);

AOI21xp5_ASAP7_75t_L g4420 ( 
.A1(n_4368),
.A2(n_4242),
.B(n_4129),
.Y(n_4420)
);

OR2x2_ASAP7_75t_L g4421 ( 
.A(n_4267),
.B(n_4234),
.Y(n_4421)
);

AO31x2_ASAP7_75t_L g4422 ( 
.A1(n_4373),
.A2(n_4189),
.A3(n_170),
.B(n_168),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_4264),
.B(n_542),
.Y(n_4423)
);

AO21x2_ASAP7_75t_L g4424 ( 
.A1(n_4327),
.A2(n_169),
.B(n_170),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_4345),
.Y(n_4425)
);

AOI21x1_ASAP7_75t_L g4426 ( 
.A1(n_4312),
.A2(n_170),
.B(n_171),
.Y(n_4426)
);

OA21x2_ASAP7_75t_L g4427 ( 
.A1(n_4367),
.A2(n_4371),
.B(n_4285),
.Y(n_4427)
);

AOI22xp33_ASAP7_75t_L g4428 ( 
.A1(n_4337),
.A2(n_174),
.B1(n_171),
.B2(n_172),
.Y(n_4428)
);

OAI22xp5_ASAP7_75t_L g4429 ( 
.A1(n_4315),
.A2(n_174),
.B1(n_171),
.B2(n_172),
.Y(n_4429)
);

OR2x2_ASAP7_75t_L g4430 ( 
.A(n_4310),
.B(n_543),
.Y(n_4430)
);

OAI21x1_ASAP7_75t_L g4431 ( 
.A1(n_4278),
.A2(n_172),
.B(n_174),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4351),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4317),
.B(n_544),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4362),
.Y(n_4434)
);

BUFx6f_ASAP7_75t_L g4435 ( 
.A(n_4332),
.Y(n_4435)
);

AO21x2_ASAP7_75t_L g4436 ( 
.A1(n_4342),
.A2(n_175),
.B(n_176),
.Y(n_4436)
);

HB1xp67_ASAP7_75t_L g4437 ( 
.A(n_4323),
.Y(n_4437)
);

HB1xp67_ASAP7_75t_L g4438 ( 
.A(n_4323),
.Y(n_4438)
);

OR2x2_ASAP7_75t_L g4439 ( 
.A(n_4347),
.B(n_544),
.Y(n_4439)
);

OAI21x1_ASAP7_75t_L g4440 ( 
.A1(n_4336),
.A2(n_176),
.B(n_177),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4301),
.Y(n_4441)
);

OAI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_4364),
.A2(n_177),
.B(n_178),
.Y(n_4442)
);

INVx3_ASAP7_75t_SL g4443 ( 
.A(n_4295),
.Y(n_4443)
);

AOI21xp5_ASAP7_75t_L g4444 ( 
.A1(n_4262),
.A2(n_178),
.B(n_179),
.Y(n_4444)
);

AOI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_4266),
.A2(n_179),
.B(n_180),
.Y(n_4445)
);

INVxp33_ASAP7_75t_L g4446 ( 
.A(n_4300),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4291),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4343),
.B(n_546),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4311),
.B(n_546),
.Y(n_4449)
);

BUFx2_ASAP7_75t_L g4450 ( 
.A(n_4282),
.Y(n_4450)
);

INVx3_ASAP7_75t_L g4451 ( 
.A(n_4332),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4325),
.Y(n_4452)
);

OAI21x1_ASAP7_75t_L g4453 ( 
.A1(n_4330),
.A2(n_182),
.B(n_183),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4333),
.Y(n_4454)
);

BUFx8_ASAP7_75t_L g4455 ( 
.A(n_4303),
.Y(n_4455)
);

OAI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4255),
.A2(n_4269),
.B(n_4290),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4333),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4346),
.B(n_547),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4319),
.B(n_547),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4357),
.Y(n_4460)
);

AOI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4270),
.A2(n_4306),
.B1(n_4277),
.B2(n_4353),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4359),
.Y(n_4462)
);

OA21x2_ASAP7_75t_L g4463 ( 
.A1(n_4352),
.A2(n_182),
.B(n_183),
.Y(n_4463)
);

HB1xp67_ASAP7_75t_L g4464 ( 
.A(n_4283),
.Y(n_4464)
);

AOI21x1_ASAP7_75t_L g4465 ( 
.A1(n_4281),
.A2(n_184),
.B(n_185),
.Y(n_4465)
);

OAI21x1_ASAP7_75t_L g4466 ( 
.A1(n_4276),
.A2(n_184),
.B(n_185),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4292),
.Y(n_4467)
);

CKINVDCx6p67_ASAP7_75t_R g4468 ( 
.A(n_4258),
.Y(n_4468)
);

A2O1A1Ixp33_ASAP7_75t_L g4469 ( 
.A1(n_4358),
.A2(n_550),
.B(n_552),
.C(n_548),
.Y(n_4469)
);

OA21x2_ASAP7_75t_L g4470 ( 
.A1(n_4314),
.A2(n_186),
.B(n_187),
.Y(n_4470)
);

OR2x2_ASAP7_75t_L g4471 ( 
.A(n_4360),
.B(n_548),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_4329),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4344),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_4335),
.A2(n_4334),
.B(n_4284),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4272),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4272),
.Y(n_4476)
);

OAI21x1_ASAP7_75t_L g4477 ( 
.A1(n_4316),
.A2(n_190),
.B(n_191),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4338),
.Y(n_4478)
);

BUFx3_ASAP7_75t_L g4479 ( 
.A(n_4257),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4338),
.Y(n_4480)
);

OAI21x1_ASAP7_75t_SL g4481 ( 
.A1(n_4355),
.A2(n_190),
.B(n_191),
.Y(n_4481)
);

AOI21xp33_ASAP7_75t_L g4482 ( 
.A1(n_4326),
.A2(n_4302),
.B(n_4261),
.Y(n_4482)
);

AOI21xp5_ASAP7_75t_L g4483 ( 
.A1(n_4370),
.A2(n_192),
.B(n_193),
.Y(n_4483)
);

INVx2_ASAP7_75t_L g4484 ( 
.A(n_4384),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4376),
.Y(n_4485)
);

OAI21x1_ASAP7_75t_L g4486 ( 
.A1(n_4374),
.A2(n_4369),
.B(n_4256),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4379),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4380),
.Y(n_4488)
);

HB1xp67_ASAP7_75t_L g4489 ( 
.A(n_4399),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4383),
.Y(n_4490)
);

AO21x1_ASAP7_75t_SL g4491 ( 
.A1(n_4464),
.A2(n_4256),
.B(n_4350),
.Y(n_4491)
);

OAI21x1_ASAP7_75t_L g4492 ( 
.A1(n_4404),
.A2(n_4366),
.B(n_4308),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4393),
.Y(n_4493)
);

OAI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4387),
.A2(n_4307),
.B(n_4363),
.Y(n_4494)
);

INVx1_ASAP7_75t_SL g4495 ( 
.A(n_4381),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4401),
.Y(n_4496)
);

NOR2xp33_ASAP7_75t_L g4497 ( 
.A(n_4446),
.B(n_4308),
.Y(n_4497)
);

OR2x6_ASAP7_75t_L g4498 ( 
.A(n_4420),
.B(n_553),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_4395),
.Y(n_4499)
);

AO31x2_ASAP7_75t_L g4500 ( 
.A1(n_4467),
.A2(n_194),
.A3(n_192),
.B(n_193),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4447),
.B(n_553),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4397),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4425),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4432),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4398),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4405),
.Y(n_4506)
);

AND2x4_ASAP7_75t_L g4507 ( 
.A(n_4450),
.B(n_555),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4416),
.Y(n_4508)
);

HB1xp67_ASAP7_75t_L g4509 ( 
.A(n_4413),
.Y(n_4509)
);

OAI21x1_ASAP7_75t_L g4510 ( 
.A1(n_4412),
.A2(n_195),
.B(n_196),
.Y(n_4510)
);

HB1xp67_ASAP7_75t_L g4511 ( 
.A(n_4392),
.Y(n_4511)
);

INVx3_ASAP7_75t_L g4512 ( 
.A(n_4479),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4421),
.B(n_556),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4457),
.Y(n_4514)
);

OAI21x1_ASAP7_75t_L g4515 ( 
.A1(n_4409),
.A2(n_195),
.B(n_196),
.Y(n_4515)
);

BUFx2_ASAP7_75t_L g4516 ( 
.A(n_4378),
.Y(n_4516)
);

INVx2_ASAP7_75t_L g4517 ( 
.A(n_4434),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4454),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4406),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4407),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4410),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_4419),
.Y(n_4522)
);

OAI21x1_ASAP7_75t_L g4523 ( 
.A1(n_4386),
.A2(n_196),
.B(n_197),
.Y(n_4523)
);

AO21x2_ASAP7_75t_L g4524 ( 
.A1(n_4460),
.A2(n_197),
.B(n_198),
.Y(n_4524)
);

INVx2_ASAP7_75t_SL g4525 ( 
.A(n_4402),
.Y(n_4525)
);

INVx3_ASAP7_75t_L g4526 ( 
.A(n_4435),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4441),
.Y(n_4527)
);

AOI21xp33_ASAP7_75t_L g4528 ( 
.A1(n_4429),
.A2(n_197),
.B(n_198),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4462),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4473),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4472),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4437),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4418),
.B(n_557),
.Y(n_4533)
);

OA21x2_ASAP7_75t_L g4534 ( 
.A1(n_4466),
.A2(n_4431),
.B(n_4475),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4438),
.Y(n_4535)
);

OR2x6_ASAP7_75t_L g4536 ( 
.A(n_4385),
.B(n_558),
.Y(n_4536)
);

INVxp67_ASAP7_75t_L g4537 ( 
.A(n_4390),
.Y(n_4537)
);

HB1xp67_ASAP7_75t_L g4538 ( 
.A(n_4452),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4476),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4411),
.Y(n_4540)
);

BUFx6f_ASAP7_75t_L g4541 ( 
.A(n_4382),
.Y(n_4541)
);

HB1xp67_ASAP7_75t_L g4542 ( 
.A(n_4394),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4470),
.Y(n_4543)
);

CKINVDCx5p33_ASAP7_75t_R g4544 ( 
.A(n_4388),
.Y(n_4544)
);

AOI21x1_ASAP7_75t_L g4545 ( 
.A1(n_4465),
.A2(n_199),
.B(n_200),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4408),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_4427),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4403),
.B(n_559),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4415),
.Y(n_4549)
);

OA21x2_ASAP7_75t_L g4550 ( 
.A1(n_4445),
.A2(n_560),
.B(n_559),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4417),
.B(n_4478),
.Y(n_4551)
);

INVx3_ASAP7_75t_L g4552 ( 
.A(n_4468),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4480),
.B(n_560),
.Y(n_4553)
);

HB1xp67_ASAP7_75t_L g4554 ( 
.A(n_4391),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4433),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4482),
.B(n_561),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4451),
.B(n_562),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4414),
.B(n_562),
.Y(n_4558)
);

BUFx2_ASAP7_75t_L g4559 ( 
.A(n_4455),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4463),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4436),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4440),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4430),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4459),
.B(n_564),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4453),
.Y(n_4565)
);

INVx2_ASAP7_75t_SL g4566 ( 
.A(n_4375),
.Y(n_4566)
);

AOI21xp5_ASAP7_75t_L g4567 ( 
.A1(n_4456),
.A2(n_199),
.B(n_200),
.Y(n_4567)
);

AND2x4_ASAP7_75t_L g4568 ( 
.A(n_4375),
.B(n_565),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4443),
.B(n_565),
.Y(n_4569)
);

INVx3_ASAP7_75t_L g4570 ( 
.A(n_4382),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4422),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4422),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4477),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4423),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4426),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4424),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4471),
.Y(n_4577)
);

OR2x2_ASAP7_75t_L g4578 ( 
.A(n_4439),
.B(n_566),
.Y(n_4578)
);

NOR2xp33_ASAP7_75t_L g4579 ( 
.A(n_4389),
.B(n_566),
.Y(n_4579)
);

INVx3_ASAP7_75t_L g4580 ( 
.A(n_4474),
.Y(n_4580)
);

AOI21x1_ASAP7_75t_L g4581 ( 
.A1(n_4396),
.A2(n_201),
.B(n_202),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4377),
.Y(n_4582)
);

HB1xp67_ASAP7_75t_L g4583 ( 
.A(n_4400),
.Y(n_4583)
);

INVx3_ASAP7_75t_L g4584 ( 
.A(n_4448),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4449),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4458),
.B(n_567),
.Y(n_4586)
);

AO21x2_ASAP7_75t_L g4587 ( 
.A1(n_4444),
.A2(n_201),
.B(n_202),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4481),
.Y(n_4588)
);

BUFx3_ASAP7_75t_L g4589 ( 
.A(n_4461),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4442),
.B(n_4483),
.Y(n_4590)
);

OAI21x1_ASAP7_75t_L g4591 ( 
.A1(n_4428),
.A2(n_203),
.B(n_205),
.Y(n_4591)
);

INVxp67_ASAP7_75t_L g4592 ( 
.A(n_4469),
.Y(n_4592)
);

BUFx3_ASAP7_75t_L g4593 ( 
.A(n_4455),
.Y(n_4593)
);

OAI21x1_ASAP7_75t_L g4594 ( 
.A1(n_4374),
.A2(n_203),
.B(n_205),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4399),
.B(n_570),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4376),
.Y(n_4596)
);

INVx3_ASAP7_75t_L g4597 ( 
.A(n_4479),
.Y(n_4597)
);

BUFx6f_ASAP7_75t_L g4598 ( 
.A(n_4382),
.Y(n_4598)
);

INVx3_ASAP7_75t_L g4599 ( 
.A(n_4479),
.Y(n_4599)
);

AOI21xp5_ASAP7_75t_L g4600 ( 
.A1(n_4385),
.A2(n_205),
.B(n_206),
.Y(n_4600)
);

OAI21x1_ASAP7_75t_L g4601 ( 
.A1(n_4492),
.A2(n_206),
.B(n_207),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4529),
.Y(n_4602)
);

AOI22xp33_ASAP7_75t_L g4603 ( 
.A1(n_4589),
.A2(n_572),
.B1(n_574),
.B2(n_571),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4509),
.B(n_206),
.Y(n_4604)
);

OR2x2_ASAP7_75t_L g4605 ( 
.A(n_4511),
.B(n_207),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4504),
.Y(n_4606)
);

HB1xp67_ASAP7_75t_L g4607 ( 
.A(n_4489),
.Y(n_4607)
);

OAI22xp5_ASAP7_75t_L g4608 ( 
.A1(n_4536),
.A2(n_4592),
.B1(n_4583),
.B2(n_4590),
.Y(n_4608)
);

AO21x2_ASAP7_75t_L g4609 ( 
.A1(n_4546),
.A2(n_208),
.B(n_209),
.Y(n_4609)
);

OAI22xp33_ASAP7_75t_L g4610 ( 
.A1(n_4536),
.A2(n_574),
.B1(n_575),
.B2(n_571),
.Y(n_4610)
);

OAI22xp5_ASAP7_75t_L g4611 ( 
.A1(n_4558),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.Y(n_4611)
);

BUFx4f_ASAP7_75t_SL g4612 ( 
.A(n_4593),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4530),
.Y(n_4613)
);

OAI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4498),
.A2(n_214),
.B1(n_211),
.B2(n_212),
.Y(n_4614)
);

AO21x2_ASAP7_75t_L g4615 ( 
.A1(n_4542),
.A2(n_212),
.B(n_214),
.Y(n_4615)
);

AOI22xp33_ASAP7_75t_SL g4616 ( 
.A1(n_4494),
.A2(n_579),
.B1(n_580),
.B2(n_578),
.Y(n_4616)
);

OAI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_4498),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_4517),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4499),
.Y(n_4619)
);

INVx3_ASAP7_75t_L g4620 ( 
.A(n_4512),
.Y(n_4620)
);

OAI21x1_ASAP7_75t_L g4621 ( 
.A1(n_4486),
.A2(n_216),
.B(n_217),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4514),
.Y(n_4622)
);

AOI21xp33_ASAP7_75t_L g4623 ( 
.A1(n_4579),
.A2(n_581),
.B(n_579),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4485),
.Y(n_4624)
);

OA21x2_ASAP7_75t_L g4625 ( 
.A1(n_4547),
.A2(n_218),
.B(n_219),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4487),
.Y(n_4626)
);

AOI22xp33_ASAP7_75t_L g4627 ( 
.A1(n_4580),
.A2(n_584),
.B1(n_585),
.B2(n_583),
.Y(n_4627)
);

AOI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4528),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_4628)
);

AOI22xp33_ASAP7_75t_L g4629 ( 
.A1(n_4587),
.A2(n_587),
.B1(n_588),
.B2(n_586),
.Y(n_4629)
);

BUFx2_ASAP7_75t_L g4630 ( 
.A(n_4516),
.Y(n_4630)
);

AOI322xp5_ASAP7_75t_L g4631 ( 
.A1(n_4576),
.A2(n_225),
.A3(n_224),
.B1(n_222),
.B2(n_220),
.C1(n_221),
.C2(n_223),
.Y(n_4631)
);

OAI22xp33_ASAP7_75t_L g4632 ( 
.A1(n_4600),
.A2(n_4581),
.B1(n_4550),
.B2(n_4543),
.Y(n_4632)
);

INVx3_ASAP7_75t_L g4633 ( 
.A(n_4597),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4488),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4490),
.Y(n_4635)
);

OAI22xp33_ASAP7_75t_L g4636 ( 
.A1(n_4574),
.A2(n_590),
.B1(n_591),
.B2(n_589),
.Y(n_4636)
);

AOI22xp33_ASAP7_75t_L g4637 ( 
.A1(n_4577),
.A2(n_594),
.B1(n_595),
.B2(n_593),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4493),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_SL g4639 ( 
.A(n_4537),
.B(n_593),
.Y(n_4639)
);

AOI22xp33_ASAP7_75t_L g4640 ( 
.A1(n_4584),
.A2(n_4563),
.B1(n_4573),
.B2(n_4585),
.Y(n_4640)
);

AOI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_4588),
.A2(n_598),
.B1(n_599),
.B2(n_597),
.Y(n_4641)
);

AOI22xp33_ASAP7_75t_L g4642 ( 
.A1(n_4555),
.A2(n_601),
.B1(n_602),
.B2(n_599),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4508),
.B(n_601),
.Y(n_4643)
);

OAI22xp5_ASAP7_75t_L g4644 ( 
.A1(n_4566),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_4644)
);

OAI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4561),
.A2(n_603),
.B1(n_604),
.B2(n_602),
.Y(n_4645)
);

OAI22xp5_ASAP7_75t_L g4646 ( 
.A1(n_4495),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4551),
.B(n_224),
.Y(n_4647)
);

AOI22xp33_ASAP7_75t_L g4648 ( 
.A1(n_4575),
.A2(n_607),
.B1(n_608),
.B2(n_606),
.Y(n_4648)
);

AOI22xp33_ASAP7_75t_L g4649 ( 
.A1(n_4524),
.A2(n_612),
.B1(n_613),
.B2(n_611),
.Y(n_4649)
);

AOI222xp33_ASAP7_75t_L g4650 ( 
.A1(n_4586),
.A2(n_227),
.B1(n_229),
.B2(n_225),
.C1(n_226),
.C2(n_228),
.Y(n_4650)
);

OAI332xp33_ASAP7_75t_L g4651 ( 
.A1(n_4549),
.A2(n_232),
.A3(n_231),
.B1(n_229),
.B2(n_233),
.B3(n_226),
.C1(n_227),
.C2(n_230),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4596),
.Y(n_4652)
);

AOI22xp33_ASAP7_75t_L g4653 ( 
.A1(n_4556),
.A2(n_612),
.B1(n_614),
.B2(n_611),
.Y(n_4653)
);

OR2x2_ASAP7_75t_L g4654 ( 
.A(n_4531),
.B(n_230),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_4544),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4599),
.B(n_232),
.Y(n_4656)
);

AND2x4_ASAP7_75t_L g4657 ( 
.A(n_4521),
.B(n_615),
.Y(n_4657)
);

BUFx3_ASAP7_75t_L g4658 ( 
.A(n_4559),
.Y(n_4658)
);

INVx2_ASAP7_75t_SL g4659 ( 
.A(n_4525),
.Y(n_4659)
);

AOI22xp33_ASAP7_75t_L g4660 ( 
.A1(n_4562),
.A2(n_617),
.B1(n_618),
.B2(n_616),
.Y(n_4660)
);

NAND2xp5_ASAP7_75t_L g4661 ( 
.A(n_4522),
.B(n_617),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4502),
.Y(n_4662)
);

INVx4_ASAP7_75t_L g4663 ( 
.A(n_4541),
.Y(n_4663)
);

HB1xp67_ASAP7_75t_L g4664 ( 
.A(n_4554),
.Y(n_4664)
);

INVx1_ASAP7_75t_SL g4665 ( 
.A(n_4569),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4505),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4503),
.Y(n_4667)
);

OAI22xp5_ASAP7_75t_L g4668 ( 
.A1(n_4526),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4484),
.B(n_235),
.Y(n_4669)
);

AOI221xp5_ASAP7_75t_SL g4670 ( 
.A1(n_4539),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.C(n_239),
.Y(n_4670)
);

AOI22xp33_ASAP7_75t_L g4671 ( 
.A1(n_4565),
.A2(n_621),
.B1(n_622),
.B2(n_619),
.Y(n_4671)
);

OAI22xp5_ASAP7_75t_L g4672 ( 
.A1(n_4570),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_4672)
);

NAND3xp33_ASAP7_75t_L g4673 ( 
.A(n_4582),
.B(n_623),
.C(n_622),
.Y(n_4673)
);

AOI221xp5_ASAP7_75t_L g4674 ( 
.A1(n_4560),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_4674)
);

OAI22xp33_ASAP7_75t_L g4675 ( 
.A1(n_4545),
.A2(n_625),
.B1(n_626),
.B2(n_624),
.Y(n_4675)
);

AOI22xp33_ASAP7_75t_L g4676 ( 
.A1(n_4513),
.A2(n_4591),
.B1(n_4533),
.B2(n_4497),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4496),
.Y(n_4677)
);

OAI221xp5_ASAP7_75t_L g4678 ( 
.A1(n_4578),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.C(n_246),
.Y(n_4678)
);

AOI221xp5_ASAP7_75t_L g4679 ( 
.A1(n_4501),
.A2(n_4595),
.B1(n_4571),
.B2(n_4572),
.C(n_4540),
.Y(n_4679)
);

HB1xp67_ASAP7_75t_L g4680 ( 
.A(n_4532),
.Y(n_4680)
);

INVx5_ASAP7_75t_L g4681 ( 
.A(n_4568),
.Y(n_4681)
);

INVx3_ASAP7_75t_L g4682 ( 
.A(n_4541),
.Y(n_4682)
);

HB1xp67_ASAP7_75t_L g4683 ( 
.A(n_4535),
.Y(n_4683)
);

AOI221xp5_ASAP7_75t_L g4684 ( 
.A1(n_4538),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.C(n_248),
.Y(n_4684)
);

AOI22xp33_ASAP7_75t_L g4685 ( 
.A1(n_4548),
.A2(n_628),
.B1(n_629),
.B2(n_627),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4506),
.Y(n_4686)
);

AND2x2_ASAP7_75t_SL g4687 ( 
.A(n_4507),
.B(n_627),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4519),
.Y(n_4688)
);

AOI221xp5_ASAP7_75t_L g4689 ( 
.A1(n_4553),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_4689)
);

BUFx2_ASAP7_75t_L g4690 ( 
.A(n_4520),
.Y(n_4690)
);

OAI22xp5_ASAP7_75t_L g4691 ( 
.A1(n_4598),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_4691)
);

BUFx6f_ASAP7_75t_L g4692 ( 
.A(n_4598),
.Y(n_4692)
);

BUFx2_ASAP7_75t_L g4693 ( 
.A(n_4534),
.Y(n_4693)
);

OAI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4527),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4491),
.B(n_253),
.Y(n_4695)
);

HB1xp67_ASAP7_75t_L g4696 ( 
.A(n_4518),
.Y(n_4696)
);

AOI22xp33_ASAP7_75t_L g4697 ( 
.A1(n_4564),
.A2(n_632),
.B1(n_634),
.B2(n_630),
.Y(n_4697)
);

BUFx8_ASAP7_75t_SL g4698 ( 
.A(n_4557),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4510),
.B(n_253),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4523),
.B(n_632),
.Y(n_4700)
);

AOI22xp33_ASAP7_75t_SL g4701 ( 
.A1(n_4594),
.A2(n_635),
.B1(n_636),
.B2(n_634),
.Y(n_4701)
);

AND2x6_ASAP7_75t_L g4702 ( 
.A(n_4500),
.B(n_636),
.Y(n_4702)
);

AOI22xp33_ASAP7_75t_L g4703 ( 
.A1(n_4515),
.A2(n_639),
.B1(n_640),
.B2(n_637),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4500),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4511),
.B(n_254),
.Y(n_4705)
);

NOR2xp33_ASAP7_75t_SL g4706 ( 
.A(n_4544),
.B(n_639),
.Y(n_4706)
);

A2O1A1Ixp33_ASAP7_75t_L g4707 ( 
.A1(n_4567),
.A2(n_641),
.B(n_642),
.C(n_640),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4504),
.Y(n_4708)
);

OAI21x1_ASAP7_75t_L g4709 ( 
.A1(n_4492),
.A2(n_254),
.B(n_255),
.Y(n_4709)
);

CKINVDCx5p33_ASAP7_75t_R g4710 ( 
.A(n_4544),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4529),
.Y(n_4711)
);

OAI221xp5_ASAP7_75t_L g4712 ( 
.A1(n_4567),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.C(n_258),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4511),
.B(n_255),
.Y(n_4713)
);

AND2x4_ASAP7_75t_SL g4714 ( 
.A(n_4552),
.B(n_644),
.Y(n_4714)
);

OAI22xp33_ASAP7_75t_L g4715 ( 
.A1(n_4536),
.A2(n_646),
.B1(n_648),
.B2(n_645),
.Y(n_4715)
);

OAI21x1_ASAP7_75t_L g4716 ( 
.A1(n_4492),
.A2(n_256),
.B(n_259),
.Y(n_4716)
);

OR2x2_ASAP7_75t_L g4717 ( 
.A(n_4509),
.B(n_259),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4529),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4511),
.B(n_260),
.Y(n_4719)
);

OAI22xp5_ASAP7_75t_SL g4720 ( 
.A1(n_4589),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4720)
);

AOI22xp33_ASAP7_75t_L g4721 ( 
.A1(n_4589),
.A2(n_646),
.B1(n_648),
.B2(n_645),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4529),
.Y(n_4722)
);

OAI21x1_ASAP7_75t_L g4723 ( 
.A1(n_4492),
.A2(n_262),
.B(n_264),
.Y(n_4723)
);

AOI22xp33_ASAP7_75t_L g4724 ( 
.A1(n_4589),
.A2(n_650),
.B1(n_651),
.B2(n_649),
.Y(n_4724)
);

NAND4xp25_ASAP7_75t_L g4725 ( 
.A(n_4567),
.B(n_267),
.C(n_265),
.D(n_266),
.Y(n_4725)
);

AOI211xp5_ASAP7_75t_L g4726 ( 
.A1(n_4567),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4537),
.B(n_649),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4529),
.Y(n_4728)
);

BUFx2_ASAP7_75t_L g4729 ( 
.A(n_4489),
.Y(n_4729)
);

OAI21x1_ASAP7_75t_L g4730 ( 
.A1(n_4492),
.A2(n_269),
.B(n_270),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4537),
.B(n_650),
.Y(n_4731)
);

BUFx6f_ASAP7_75t_L g4732 ( 
.A(n_4541),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4613),
.Y(n_4733)
);

HB1xp67_ASAP7_75t_L g4734 ( 
.A(n_4664),
.Y(n_4734)
);

HB1xp67_ASAP7_75t_L g4735 ( 
.A(n_4680),
.Y(n_4735)
);

AOI22xp33_ASAP7_75t_L g4736 ( 
.A1(n_4725),
.A2(n_652),
.B1(n_653),
.B2(n_651),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4602),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4729),
.B(n_270),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4620),
.B(n_270),
.Y(n_4739)
);

AOI22xp33_ASAP7_75t_L g4740 ( 
.A1(n_4712),
.A2(n_653),
.B1(n_654),
.B2(n_652),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4711),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4718),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4633),
.B(n_4665),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4722),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4728),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4640),
.B(n_271),
.Y(n_4746)
);

AND2x2_ASAP7_75t_L g4747 ( 
.A(n_4690),
.B(n_4659),
.Y(n_4747)
);

NOR2x1_ASAP7_75t_R g4748 ( 
.A(n_4681),
.B(n_272),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4622),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4683),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4624),
.Y(n_4751)
);

HB1xp67_ASAP7_75t_L g4752 ( 
.A(n_4696),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4634),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4626),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4693),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4679),
.B(n_656),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4635),
.Y(n_4757)
);

INVx2_ASAP7_75t_L g4758 ( 
.A(n_4606),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4677),
.B(n_4667),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4618),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4708),
.Y(n_4761)
);

NAND3xp33_ASAP7_75t_L g4762 ( 
.A(n_4726),
.B(n_273),
.C(n_274),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4638),
.Y(n_4763)
);

AND2x4_ASAP7_75t_L g4764 ( 
.A(n_4658),
.B(n_4682),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4619),
.Y(n_4765)
);

OR2x2_ASAP7_75t_L g4766 ( 
.A(n_4688),
.B(n_273),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4652),
.B(n_658),
.Y(n_4767)
);

INVx3_ASAP7_75t_L g4768 ( 
.A(n_4663),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4662),
.B(n_658),
.Y(n_4769)
);

AND2x4_ASAP7_75t_L g4770 ( 
.A(n_4666),
.B(n_4686),
.Y(n_4770)
);

AOI22xp33_ASAP7_75t_SL g4771 ( 
.A1(n_4608),
.A2(n_660),
.B1(n_661),
.B2(n_659),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4704),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4654),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4625),
.Y(n_4774)
);

INVx1_ASAP7_75t_SL g4775 ( 
.A(n_4698),
.Y(n_4775)
);

INVx2_ASAP7_75t_SL g4776 ( 
.A(n_4681),
.Y(n_4776)
);

BUFx6f_ASAP7_75t_L g4777 ( 
.A(n_4692),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4661),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4705),
.B(n_4713),
.Y(n_4779)
);

OR2x2_ASAP7_75t_L g4780 ( 
.A(n_4605),
.B(n_274),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4669),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4643),
.B(n_660),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4719),
.B(n_661),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4604),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4717),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4647),
.B(n_275),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4681),
.B(n_275),
.Y(n_4787)
);

OR2x2_ASAP7_75t_L g4788 ( 
.A(n_4676),
.B(n_275),
.Y(n_4788)
);

INVx1_ASAP7_75t_SL g4789 ( 
.A(n_4612),
.Y(n_4789)
);

HB1xp67_ASAP7_75t_L g4790 ( 
.A(n_4601),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4727),
.B(n_662),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4657),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4709),
.Y(n_4793)
);

OR2x2_ASAP7_75t_L g4794 ( 
.A(n_4731),
.B(n_276),
.Y(n_4794)
);

OR2x2_ASAP7_75t_L g4795 ( 
.A(n_4632),
.B(n_277),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4609),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4702),
.B(n_663),
.Y(n_4797)
);

NOR2xp33_ASAP7_75t_L g4798 ( 
.A(n_4655),
.B(n_1665),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4716),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4702),
.Y(n_4800)
);

INVx2_ASAP7_75t_L g4801 ( 
.A(n_4723),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4702),
.Y(n_4802)
);

AND2x2_ASAP7_75t_L g4803 ( 
.A(n_4732),
.B(n_278),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4730),
.Y(n_4804)
);

BUFx2_ASAP7_75t_L g4805 ( 
.A(n_4732),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4695),
.B(n_278),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4656),
.B(n_278),
.Y(n_4807)
);

HB1xp67_ASAP7_75t_L g4808 ( 
.A(n_4615),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4699),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_L g4810 ( 
.A(n_4710),
.B(n_1667),
.Y(n_4810)
);

INVx4_ASAP7_75t_L g4811 ( 
.A(n_4714),
.Y(n_4811)
);

AND2x2_ASAP7_75t_L g4812 ( 
.A(n_4687),
.B(n_4621),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4700),
.Y(n_4813)
);

HB1xp67_ASAP7_75t_L g4814 ( 
.A(n_4639),
.Y(n_4814)
);

OAI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4673),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_4815)
);

INVx4_ASAP7_75t_L g4816 ( 
.A(n_4706),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4675),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4694),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4611),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4641),
.Y(n_4820)
);

AND2x2_ASAP7_75t_L g4821 ( 
.A(n_4653),
.B(n_281),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4623),
.A2(n_665),
.B1(n_666),
.B2(n_664),
.Y(n_4822)
);

NOR2xp33_ASAP7_75t_L g4823 ( 
.A(n_4678),
.B(n_1671),
.Y(n_4823)
);

INVx2_ASAP7_75t_SL g4824 ( 
.A(n_4614),
.Y(n_4824)
);

AND2x2_ASAP7_75t_L g4825 ( 
.A(n_4670),
.B(n_282),
.Y(n_4825)
);

AOI22xp33_ASAP7_75t_L g4826 ( 
.A1(n_4616),
.A2(n_665),
.B1(n_666),
.B2(n_664),
.Y(n_4826)
);

AND2x2_ASAP7_75t_L g4827 ( 
.A(n_4701),
.B(n_283),
.Y(n_4827)
);

AND2x4_ASAP7_75t_L g4828 ( 
.A(n_4707),
.B(n_667),
.Y(n_4828)
);

INVx1_ASAP7_75t_SL g4829 ( 
.A(n_4720),
.Y(n_4829)
);

NOR2xp33_ASAP7_75t_L g4830 ( 
.A(n_4651),
.B(n_1680),
.Y(n_4830)
);

NAND2x1p5_ASAP7_75t_L g4831 ( 
.A(n_4610),
.B(n_669),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4645),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4617),
.Y(n_4833)
);

AND2x4_ASAP7_75t_L g4834 ( 
.A(n_4627),
.B(n_670),
.Y(n_4834)
);

OR2x2_ASAP7_75t_L g4835 ( 
.A(n_4644),
.B(n_283),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4703),
.B(n_283),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4685),
.B(n_284),
.Y(n_4837)
);

INVx1_ASAP7_75t_SL g4838 ( 
.A(n_4646),
.Y(n_4838)
);

AND2x2_ASAP7_75t_L g4839 ( 
.A(n_4649),
.B(n_284),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_4650),
.B(n_284),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4629),
.B(n_285),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4668),
.Y(n_4842)
);

NAND3xp33_ASAP7_75t_L g4843 ( 
.A(n_4684),
.B(n_285),
.C(n_286),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4697),
.B(n_285),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4672),
.Y(n_4845)
);

BUFx3_ASAP7_75t_L g4846 ( 
.A(n_4691),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4636),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4715),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4637),
.B(n_286),
.Y(n_4849)
);

NOR2xp33_ASAP7_75t_L g4850 ( 
.A(n_4689),
.B(n_1669),
.Y(n_4850)
);

HB1xp67_ASAP7_75t_L g4851 ( 
.A(n_4674),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4631),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4642),
.B(n_287),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4660),
.B(n_671),
.Y(n_4854)
);

AND2x4_ASAP7_75t_L g4855 ( 
.A(n_4671),
.B(n_672),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4628),
.B(n_672),
.Y(n_4856)
);

INVx2_ASAP7_75t_SL g4857 ( 
.A(n_4648),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4603),
.Y(n_4858)
);

AND2x4_ASAP7_75t_L g4859 ( 
.A(n_4724),
.B(n_673),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4721),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4630),
.B(n_288),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4607),
.B(n_674),
.Y(n_4862)
);

INVxp67_ASAP7_75t_SL g4863 ( 
.A(n_4664),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4613),
.Y(n_4864)
);

OAI22xp5_ASAP7_75t_L g4865 ( 
.A1(n_4608),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4630),
.B(n_289),
.Y(n_4866)
);

INVxp67_ASAP7_75t_SL g4867 ( 
.A(n_4664),
.Y(n_4867)
);

INVx1_ASAP7_75t_SL g4868 ( 
.A(n_4698),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4613),
.Y(n_4869)
);

BUFx3_ASAP7_75t_L g4870 ( 
.A(n_4612),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4607),
.B(n_675),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4613),
.Y(n_4872)
);

BUFx3_ASAP7_75t_L g4873 ( 
.A(n_4612),
.Y(n_4873)
);

BUFx2_ASAP7_75t_L g4874 ( 
.A(n_4630),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4613),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4613),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4613),
.Y(n_4877)
);

INVxp33_ASAP7_75t_SL g4878 ( 
.A(n_4655),
.Y(n_4878)
);

INVx2_ASAP7_75t_L g4879 ( 
.A(n_4874),
.Y(n_4879)
);

AND2x2_ASAP7_75t_L g4880 ( 
.A(n_4800),
.B(n_291),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4802),
.B(n_4747),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4772),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4809),
.B(n_292),
.Y(n_4883)
);

AND2x2_ASAP7_75t_L g4884 ( 
.A(n_4743),
.B(n_292),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4733),
.Y(n_4885)
);

AND2x2_ASAP7_75t_L g4886 ( 
.A(n_4805),
.B(n_294),
.Y(n_4886)
);

AND2x4_ASAP7_75t_L g4887 ( 
.A(n_4768),
.B(n_294),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4737),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4741),
.Y(n_4889)
);

INVx2_ASAP7_75t_L g4890 ( 
.A(n_4770),
.Y(n_4890)
);

HB1xp67_ASAP7_75t_L g4891 ( 
.A(n_4774),
.Y(n_4891)
);

AND2x4_ASAP7_75t_L g4892 ( 
.A(n_4764),
.B(n_295),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4773),
.B(n_295),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4744),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4758),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4745),
.Y(n_4896)
);

AND2x4_ASAP7_75t_L g4897 ( 
.A(n_4792),
.B(n_4781),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4749),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4760),
.Y(n_4899)
);

AND2x4_ASAP7_75t_L g4900 ( 
.A(n_4784),
.B(n_296),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4754),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4757),
.Y(n_4902)
);

OR2x2_ASAP7_75t_L g4903 ( 
.A(n_4785),
.B(n_296),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4779),
.B(n_297),
.Y(n_4904)
);

AND2x4_ASAP7_75t_L g4905 ( 
.A(n_4750),
.B(n_297),
.Y(n_4905)
);

INVx2_ASAP7_75t_L g4906 ( 
.A(n_4761),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4735),
.B(n_297),
.Y(n_4907)
);

NOR2x1_ASAP7_75t_L g4908 ( 
.A(n_4796),
.B(n_299),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4814),
.B(n_676),
.Y(n_4909)
);

OR2x2_ASAP7_75t_L g4910 ( 
.A(n_4778),
.B(n_299),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4763),
.Y(n_4911)
);

OR2x2_ASAP7_75t_L g4912 ( 
.A(n_4734),
.B(n_300),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4863),
.B(n_300),
.Y(n_4913)
);

AND2x2_ASAP7_75t_L g4914 ( 
.A(n_4867),
.B(n_300),
.Y(n_4914)
);

INVx4_ASAP7_75t_L g4915 ( 
.A(n_4870),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4790),
.B(n_301),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4812),
.B(n_301),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4864),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4759),
.B(n_302),
.Y(n_4919)
);

AND2x2_ASAP7_75t_L g4920 ( 
.A(n_4752),
.B(n_302),
.Y(n_4920)
);

NOR2xp67_ASAP7_75t_L g4921 ( 
.A(n_4816),
.B(n_303),
.Y(n_4921)
);

INVx1_ASAP7_75t_SL g4922 ( 
.A(n_4775),
.Y(n_4922)
);

NOR2x1_ASAP7_75t_L g4923 ( 
.A(n_4795),
.B(n_304),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4808),
.B(n_677),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4765),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4793),
.B(n_678),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4869),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4751),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4799),
.B(n_4801),
.Y(n_4929)
);

HB1xp67_ASAP7_75t_L g4930 ( 
.A(n_4755),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4872),
.Y(n_4931)
);

AND2x2_ASAP7_75t_L g4932 ( 
.A(n_4804),
.B(n_305),
.Y(n_4932)
);

OR2x6_ASAP7_75t_L g4933 ( 
.A(n_4811),
.B(n_678),
.Y(n_4933)
);

NOR2xp33_ASAP7_75t_L g4934 ( 
.A(n_4878),
.B(n_679),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4746),
.B(n_679),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4753),
.B(n_305),
.Y(n_4936)
);

BUFx2_ASAP7_75t_L g4937 ( 
.A(n_4787),
.Y(n_4937)
);

INVx4_ASAP7_75t_L g4938 ( 
.A(n_4873),
.Y(n_4938)
);

HB1xp67_ASAP7_75t_L g4939 ( 
.A(n_4742),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4875),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4738),
.B(n_306),
.Y(n_4941)
);

NAND3xp33_ASAP7_75t_L g4942 ( 
.A(n_4830),
.B(n_307),
.C(n_308),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4876),
.Y(n_4943)
);

INVx2_ASAP7_75t_L g4944 ( 
.A(n_4877),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4766),
.Y(n_4945)
);

AND2x4_ASAP7_75t_SL g4946 ( 
.A(n_4777),
.B(n_308),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4739),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4848),
.B(n_309),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4767),
.Y(n_4949)
);

NAND3xp33_ASAP7_75t_L g4950 ( 
.A(n_4851),
.B(n_309),
.C(n_310),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4769),
.Y(n_4951)
);

OR2x2_ASAP7_75t_L g4952 ( 
.A(n_4817),
.B(n_310),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4862),
.Y(n_4953)
);

INVx2_ASAP7_75t_SL g4954 ( 
.A(n_4868),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4819),
.B(n_680),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4871),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4818),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4833),
.B(n_310),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4847),
.B(n_681),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4861),
.B(n_311),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4832),
.B(n_681),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4866),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4756),
.Y(n_4963)
);

OR2x2_ASAP7_75t_L g4964 ( 
.A(n_4824),
.B(n_312),
.Y(n_4964)
);

HB1xp67_ASAP7_75t_L g4965 ( 
.A(n_4842),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4820),
.B(n_682),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4845),
.B(n_682),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4846),
.B(n_313),
.Y(n_4968)
);

NOR2xp67_ASAP7_75t_L g4969 ( 
.A(n_4797),
.B(n_4762),
.Y(n_4969)
);

INVx3_ASAP7_75t_L g4970 ( 
.A(n_4789),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4806),
.B(n_314),
.Y(n_4971)
);

AND2x4_ASAP7_75t_L g4972 ( 
.A(n_4803),
.B(n_314),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4794),
.Y(n_4973)
);

AND2x2_ASAP7_75t_L g4974 ( 
.A(n_4786),
.B(n_4807),
.Y(n_4974)
);

HB1xp67_ASAP7_75t_L g4975 ( 
.A(n_4780),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4838),
.B(n_683),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4788),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4857),
.Y(n_4978)
);

OR2x2_ASAP7_75t_L g4979 ( 
.A(n_4783),
.B(n_315),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_SL g4980 ( 
.A(n_4771),
.B(n_315),
.Y(n_4980)
);

AND2x2_ASAP7_75t_L g4981 ( 
.A(n_4829),
.B(n_315),
.Y(n_4981)
);

AND2x2_ASAP7_75t_L g4982 ( 
.A(n_4858),
.B(n_316),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4860),
.B(n_316),
.Y(n_4983)
);

INVx2_ASAP7_75t_L g4984 ( 
.A(n_4782),
.Y(n_4984)
);

NAND2xp33_ASAP7_75t_L g4985 ( 
.A(n_4825),
.B(n_316),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4791),
.Y(n_4986)
);

BUFx2_ASAP7_75t_L g4987 ( 
.A(n_4831),
.Y(n_4987)
);

AND2x2_ASAP7_75t_L g4988 ( 
.A(n_4798),
.B(n_317),
.Y(n_4988)
);

INVx3_ASAP7_75t_L g4989 ( 
.A(n_4835),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4810),
.B(n_318),
.Y(n_4990)
);

AOI21xp5_ASAP7_75t_SL g4991 ( 
.A1(n_4828),
.A2(n_318),
.B(n_319),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4852),
.B(n_319),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4827),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_4823),
.B(n_684),
.Y(n_4994)
);

INVxp67_ASAP7_75t_SL g4995 ( 
.A(n_4865),
.Y(n_4995)
);

INVx2_ASAP7_75t_L g4996 ( 
.A(n_4821),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4836),
.Y(n_4997)
);

NOR2x1_ASAP7_75t_L g4998 ( 
.A(n_4843),
.B(n_319),
.Y(n_4998)
);

AND2x4_ASAP7_75t_L g4999 ( 
.A(n_4853),
.B(n_320),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4815),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4840),
.B(n_320),
.Y(n_5001)
);

NOR3xp33_ASAP7_75t_L g5002 ( 
.A(n_4850),
.B(n_320),
.C(n_321),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4837),
.B(n_321),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4844),
.B(n_321),
.Y(n_5004)
);

OR2x2_ASAP7_75t_L g5005 ( 
.A(n_4856),
.B(n_322),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4841),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4849),
.B(n_323),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4839),
.Y(n_5008)
);

INVx2_ASAP7_75t_SL g5009 ( 
.A(n_4859),
.Y(n_5009)
);

INVxp67_ASAP7_75t_SL g5010 ( 
.A(n_4854),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4834),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4822),
.B(n_4740),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_4855),
.B(n_323),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4736),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4826),
.B(n_323),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_SL g5016 ( 
.A(n_4776),
.B(n_324),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4772),
.Y(n_5017)
);

AND2x4_ASAP7_75t_L g5018 ( 
.A(n_4776),
.B(n_325),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4813),
.B(n_685),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_4813),
.B(n_686),
.Y(n_5020)
);

AND2x4_ASAP7_75t_L g5021 ( 
.A(n_4776),
.B(n_325),
.Y(n_5021)
);

AOI22xp33_ASAP7_75t_L g5022 ( 
.A1(n_4830),
.A2(n_688),
.B1(n_689),
.B2(n_687),
.Y(n_5022)
);

OAI21xp33_ASAP7_75t_L g5023 ( 
.A1(n_4830),
.A2(n_326),
.B(n_327),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_4874),
.B(n_326),
.Y(n_5024)
);

OR2x2_ASAP7_75t_L g5025 ( 
.A(n_4809),
.B(n_326),
.Y(n_5025)
);

INVx3_ASAP7_75t_L g5026 ( 
.A(n_4764),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4772),
.Y(n_5027)
);

OR2x2_ASAP7_75t_L g5028 ( 
.A(n_4809),
.B(n_327),
.Y(n_5028)
);

HB1xp67_ASAP7_75t_L g5029 ( 
.A(n_4774),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_SL g5030 ( 
.A(n_4776),
.B(n_327),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4772),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4772),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4772),
.Y(n_5033)
);

AND2x2_ASAP7_75t_L g5034 ( 
.A(n_4874),
.B(n_328),
.Y(n_5034)
);

AND2x2_ASAP7_75t_L g5035 ( 
.A(n_4874),
.B(n_328),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4772),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_4772),
.Y(n_5037)
);

AND2x2_ASAP7_75t_L g5038 ( 
.A(n_4874),
.B(n_329),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4874),
.B(n_330),
.Y(n_5039)
);

HB1xp67_ASAP7_75t_L g5040 ( 
.A(n_4774),
.Y(n_5040)
);

INVxp67_ASAP7_75t_L g5041 ( 
.A(n_4748),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4772),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4874),
.B(n_331),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4874),
.B(n_331),
.Y(n_5044)
);

NOR2x1p5_ASAP7_75t_L g5045 ( 
.A(n_4816),
.B(n_332),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4772),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4813),
.B(n_690),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4772),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_4874),
.B(n_333),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4813),
.B(n_691),
.Y(n_5050)
);

AOI33xp33_ASAP7_75t_L g5051 ( 
.A1(n_5022),
.A2(n_335),
.A3(n_337),
.B1(n_333),
.B2(n_334),
.B3(n_336),
.Y(n_5051)
);

NOR3xp33_ASAP7_75t_L g5052 ( 
.A(n_4942),
.B(n_334),
.C(n_335),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4891),
.Y(n_5053)
);

OR2x2_ASAP7_75t_L g5054 ( 
.A(n_4978),
.B(n_338),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_5029),
.Y(n_5055)
);

INVx2_ASAP7_75t_L g5056 ( 
.A(n_4970),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_5026),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4963),
.B(n_338),
.Y(n_5058)
);

AND2x2_ASAP7_75t_L g5059 ( 
.A(n_4937),
.B(n_4881),
.Y(n_5059)
);

HB1xp67_ASAP7_75t_L g5060 ( 
.A(n_4930),
.Y(n_5060)
);

AND2x2_ASAP7_75t_L g5061 ( 
.A(n_4879),
.B(n_339),
.Y(n_5061)
);

AND2x2_ASAP7_75t_L g5062 ( 
.A(n_4975),
.B(n_341),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_5040),
.Y(n_5063)
);

NOR2xp33_ASAP7_75t_L g5064 ( 
.A(n_4915),
.B(n_342),
.Y(n_5064)
);

AND2x2_ASAP7_75t_L g5065 ( 
.A(n_4989),
.B(n_343),
.Y(n_5065)
);

AO21x2_ASAP7_75t_L g5066 ( 
.A1(n_4924),
.A2(n_344),
.B(n_345),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_4987),
.B(n_344),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_5010),
.B(n_346),
.Y(n_5068)
);

AOI33xp33_ASAP7_75t_L g5069 ( 
.A1(n_5000),
.A2(n_350),
.A3(n_352),
.B1(n_347),
.B2(n_349),
.B3(n_351),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4973),
.B(n_352),
.Y(n_5070)
);

AO22x1_ASAP7_75t_L g5071 ( 
.A1(n_4908),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4882),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_5017),
.Y(n_5073)
);

INVxp67_ASAP7_75t_SL g5074 ( 
.A(n_4921),
.Y(n_5074)
);

OR2x2_ASAP7_75t_L g5075 ( 
.A(n_4957),
.B(n_4977),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_4984),
.B(n_353),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_4954),
.Y(n_5077)
);

OAI22xp5_ASAP7_75t_L g5078 ( 
.A1(n_4995),
.A2(n_4969),
.B1(n_4965),
.B2(n_4923),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4890),
.B(n_354),
.Y(n_5079)
);

NAND4xp25_ASAP7_75t_L g5080 ( 
.A(n_5023),
.B(n_356),
.C(n_354),
.D(n_355),
.Y(n_5080)
);

NOR3xp33_ASAP7_75t_L g5081 ( 
.A(n_4985),
.B(n_355),
.C(n_356),
.Y(n_5081)
);

AOI222xp33_ASAP7_75t_L g5082 ( 
.A1(n_4980),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.C1(n_693),
.C2(n_692),
.Y(n_5082)
);

INVx4_ASAP7_75t_L g5083 ( 
.A(n_4938),
.Y(n_5083)
);

AOI22xp33_ASAP7_75t_L g5084 ( 
.A1(n_5002),
.A2(n_359),
.B1(n_693),
.B2(n_692),
.Y(n_5084)
);

HB1xp67_ASAP7_75t_L g5085 ( 
.A(n_4939),
.Y(n_5085)
);

OAI221xp5_ASAP7_75t_L g5086 ( 
.A1(n_4998),
.A2(n_5012),
.B1(n_5041),
.B2(n_4991),
.C(n_4950),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_5027),
.Y(n_5087)
);

AND2x2_ASAP7_75t_L g5088 ( 
.A(n_4986),
.B(n_694),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4917),
.B(n_698),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_5031),
.Y(n_5090)
);

AND2x4_ASAP7_75t_L g5091 ( 
.A(n_4897),
.B(n_699),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4945),
.B(n_4916),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_4953),
.B(n_702),
.Y(n_5093)
);

AOI22xp33_ASAP7_75t_L g5094 ( 
.A1(n_5014),
.A2(n_706),
.B1(n_703),
.B2(n_705),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_5032),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5033),
.Y(n_5096)
);

INVx3_ASAP7_75t_L g5097 ( 
.A(n_4892),
.Y(n_5097)
);

INVx3_ASAP7_75t_L g5098 ( 
.A(n_4922),
.Y(n_5098)
);

INVx4_ASAP7_75t_L g5099 ( 
.A(n_4933),
.Y(n_5099)
);

AND2x4_ASAP7_75t_L g5100 ( 
.A(n_4947),
.B(n_707),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4929),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_4956),
.B(n_4996),
.Y(n_5102)
);

NAND2xp33_ASAP7_75t_SL g5103 ( 
.A(n_5045),
.B(n_708),
.Y(n_5103)
);

AND2x2_ASAP7_75t_L g5104 ( 
.A(n_4949),
.B(n_708),
.Y(n_5104)
);

AOI221xp5_ASAP7_75t_L g5105 ( 
.A1(n_4994),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.C(n_712),
.Y(n_5105)
);

OAI31xp33_ASAP7_75t_L g5106 ( 
.A1(n_5016),
.A2(n_1674),
.A3(n_1675),
.B(n_1673),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_5036),
.Y(n_5107)
);

AOI22xp33_ASAP7_75t_L g5108 ( 
.A1(n_4993),
.A2(n_714),
.B1(n_711),
.B2(n_713),
.Y(n_5108)
);

AOI221xp5_ASAP7_75t_SL g5109 ( 
.A1(n_5030),
.A2(n_1678),
.B1(n_717),
.B2(n_715),
.C(n_716),
.Y(n_5109)
);

AOI22xp33_ASAP7_75t_L g5110 ( 
.A1(n_4997),
.A2(n_5006),
.B1(n_5008),
.B2(n_4951),
.Y(n_5110)
);

NOR3xp33_ASAP7_75t_SL g5111 ( 
.A(n_4909),
.B(n_718),
.C(n_719),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_4962),
.B(n_722),
.Y(n_5112)
);

NOR3xp33_ASAP7_75t_L g5113 ( 
.A(n_4926),
.B(n_723),
.C(n_724),
.Y(n_5113)
);

AND2x2_ASAP7_75t_L g5114 ( 
.A(n_4974),
.B(n_724),
.Y(n_5114)
);

OAI22xp5_ASAP7_75t_L g5115 ( 
.A1(n_4952),
.A2(n_728),
.B1(n_725),
.B2(n_727),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_5037),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_4884),
.B(n_730),
.Y(n_5117)
);

AO21x2_ASAP7_75t_L g5118 ( 
.A1(n_4913),
.A2(n_730),
.B(n_731),
.Y(n_5118)
);

INVx4_ASAP7_75t_L g5119 ( 
.A(n_4887),
.Y(n_5119)
);

AOI33xp33_ASAP7_75t_L g5120 ( 
.A1(n_4992),
.A2(n_734),
.A3(n_736),
.B1(n_732),
.B2(n_733),
.B3(n_735),
.Y(n_5120)
);

INVx2_ASAP7_75t_L g5121 ( 
.A(n_4895),
.Y(n_5121)
);

INVx5_ASAP7_75t_L g5122 ( 
.A(n_4981),
.Y(n_5122)
);

OAI221xp5_ASAP7_75t_L g5123 ( 
.A1(n_5005),
.A2(n_737),
.B1(n_732),
.B2(n_735),
.C(n_738),
.Y(n_5123)
);

INVx2_ASAP7_75t_L g5124 ( 
.A(n_4899),
.Y(n_5124)
);

OAI211xp5_ASAP7_75t_SL g5125 ( 
.A1(n_4966),
.A2(n_739),
.B(n_737),
.C(n_738),
.Y(n_5125)
);

INVx2_ASAP7_75t_L g5126 ( 
.A(n_4906),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_SL g5127 ( 
.A(n_5009),
.B(n_4905),
.Y(n_5127)
);

INVx2_ASAP7_75t_L g5128 ( 
.A(n_4925),
.Y(n_5128)
);

AND2x4_ASAP7_75t_SL g5129 ( 
.A(n_5018),
.B(n_740),
.Y(n_5129)
);

OAI211xp5_ASAP7_75t_L g5130 ( 
.A1(n_5015),
.A2(n_742),
.B(n_740),
.C(n_741),
.Y(n_5130)
);

AND2x2_ASAP7_75t_L g5131 ( 
.A(n_5011),
.B(n_742),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_4883),
.B(n_743),
.Y(n_5132)
);

OR2x2_ASAP7_75t_L g5133 ( 
.A(n_4928),
.B(n_744),
.Y(n_5133)
);

INVx2_ASAP7_75t_SL g5134 ( 
.A(n_5021),
.Y(n_5134)
);

INVx2_ASAP7_75t_L g5135 ( 
.A(n_4943),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4944),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_4919),
.B(n_744),
.Y(n_5137)
);

OAI31xp33_ASAP7_75t_L g5138 ( 
.A1(n_5001),
.A2(n_1677),
.A3(n_1678),
.B(n_1676),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_5042),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_5046),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5048),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_4885),
.Y(n_5142)
);

OR2x2_ASAP7_75t_L g5143 ( 
.A(n_4903),
.B(n_750),
.Y(n_5143)
);

OR2x2_ASAP7_75t_L g5144 ( 
.A(n_4888),
.B(n_750),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_5024),
.B(n_751),
.Y(n_5145)
);

AOI22xp33_ASAP7_75t_L g5146 ( 
.A1(n_4934),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_5146)
);

NAND3xp33_ASAP7_75t_L g5147 ( 
.A(n_4955),
.B(n_754),
.C(n_755),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4889),
.Y(n_5148)
);

HB1xp67_ASAP7_75t_L g5149 ( 
.A(n_4894),
.Y(n_5149)
);

OR2x2_ASAP7_75t_L g5150 ( 
.A(n_4896),
.B(n_756),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_4898),
.Y(n_5151)
);

INVx3_ASAP7_75t_L g5152 ( 
.A(n_4900),
.Y(n_5152)
);

INVx2_ASAP7_75t_SL g5153 ( 
.A(n_4886),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_4901),
.Y(n_5154)
);

OAI211xp5_ASAP7_75t_L g5155 ( 
.A1(n_4961),
.A2(n_761),
.B(n_757),
.C(n_759),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4902),
.Y(n_5156)
);

INVxp67_ASAP7_75t_L g5157 ( 
.A(n_4964),
.Y(n_5157)
);

AOI221xp5_ASAP7_75t_L g5158 ( 
.A1(n_4976),
.A2(n_763),
.B1(n_759),
.B2(n_761),
.C(n_764),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4911),
.Y(n_5159)
);

NAND2xp5_ASAP7_75t_L g5160 ( 
.A(n_4932),
.B(n_764),
.Y(n_5160)
);

OAI221xp5_ASAP7_75t_L g5161 ( 
.A1(n_4935),
.A2(n_767),
.B1(n_765),
.B2(n_766),
.C(n_768),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4918),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4927),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4931),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4940),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_4936),
.Y(n_5166)
);

CKINVDCx5p33_ASAP7_75t_R g5167 ( 
.A(n_4946),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5034),
.B(n_5035),
.Y(n_5168)
);

INVx4_ASAP7_75t_L g5169 ( 
.A(n_4972),
.Y(n_5169)
);

NOR2xp33_ASAP7_75t_L g5170 ( 
.A(n_4967),
.B(n_770),
.Y(n_5170)
);

OAI31xp33_ASAP7_75t_L g5171 ( 
.A1(n_4968),
.A2(n_1668),
.A3(n_1670),
.B(n_1667),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_5038),
.B(n_771),
.Y(n_5172)
);

AND2x4_ASAP7_75t_L g5173 ( 
.A(n_5039),
.B(n_771),
.Y(n_5173)
);

AOI22xp33_ASAP7_75t_L g5174 ( 
.A1(n_5052),
.A2(n_4959),
.B1(n_4999),
.B2(n_4983),
.Y(n_5174)
);

NOR2xp33_ASAP7_75t_L g5175 ( 
.A(n_5083),
.B(n_5047),
.Y(n_5175)
);

NAND2x1p5_ASAP7_75t_L g5176 ( 
.A(n_5098),
.B(n_5043),
.Y(n_5176)
);

INVx3_ASAP7_75t_L g5177 ( 
.A(n_5169),
.Y(n_5177)
);

HB1xp67_ASAP7_75t_L g5178 ( 
.A(n_5122),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5060),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5085),
.Y(n_5180)
);

INVx2_ASAP7_75t_SL g5181 ( 
.A(n_5122),
.Y(n_5181)
);

AND2x2_ASAP7_75t_L g5182 ( 
.A(n_5122),
.B(n_4948),
.Y(n_5182)
);

AOI22xp33_ASAP7_75t_L g5183 ( 
.A1(n_5081),
.A2(n_4982),
.B1(n_4990),
.B2(n_4988),
.Y(n_5183)
);

INVxp67_ASAP7_75t_L g5184 ( 
.A(n_5074),
.Y(n_5184)
);

NAND4xp25_ASAP7_75t_SL g5185 ( 
.A(n_5082),
.B(n_5069),
.C(n_5051),
.D(n_5109),
.Y(n_5185)
);

NOR3xp33_ASAP7_75t_L g5186 ( 
.A(n_5078),
.B(n_5020),
.C(n_5019),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5149),
.Y(n_5187)
);

INVx1_ASAP7_75t_SL g5188 ( 
.A(n_5103),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_5153),
.B(n_4914),
.Y(n_5189)
);

CKINVDCx14_ASAP7_75t_R g5190 ( 
.A(n_5167),
.Y(n_5190)
);

OR2x2_ASAP7_75t_L g5191 ( 
.A(n_5092),
.B(n_5025),
.Y(n_5191)
);

NOR2x1_ASAP7_75t_L g5192 ( 
.A(n_5099),
.B(n_4912),
.Y(n_5192)
);

AND2x4_ASAP7_75t_L g5193 ( 
.A(n_5119),
.B(n_4880),
.Y(n_5193)
);

INVx3_ASAP7_75t_L g5194 ( 
.A(n_5097),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5102),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_5053),
.Y(n_5196)
);

AND2x2_ASAP7_75t_L g5197 ( 
.A(n_5056),
.B(n_4958),
.Y(n_5197)
);

AND2x2_ASAP7_75t_L g5198 ( 
.A(n_5059),
.B(n_5077),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_5057),
.B(n_5044),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_5055),
.Y(n_5200)
);

AND2x2_ASAP7_75t_L g5201 ( 
.A(n_5168),
.B(n_5049),
.Y(n_5201)
);

AND2x4_ASAP7_75t_L g5202 ( 
.A(n_5152),
.B(n_5134),
.Y(n_5202)
);

INVx3_ASAP7_75t_L g5203 ( 
.A(n_5091),
.Y(n_5203)
);

OR2x2_ASAP7_75t_L g5204 ( 
.A(n_5157),
.B(n_5028),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5063),
.Y(n_5205)
);

AND2x2_ASAP7_75t_L g5206 ( 
.A(n_5166),
.B(n_4904),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5133),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_5066),
.B(n_4907),
.Y(n_5208)
);

NOR2x1_ASAP7_75t_L g5209 ( 
.A(n_5118),
.B(n_4910),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_5075),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_5139),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_5054),
.Y(n_5212)
);

NAND2x1_ASAP7_75t_L g5213 ( 
.A(n_5101),
.B(n_4920),
.Y(n_5213)
);

AOI22xp33_ASAP7_75t_L g5214 ( 
.A1(n_5086),
.A2(n_5007),
.B1(n_5003),
.B2(n_5004),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5127),
.B(n_4893),
.Y(n_5215)
);

AND2x2_ASAP7_75t_L g5216 ( 
.A(n_5110),
.B(n_4941),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_5071),
.B(n_5050),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_5067),
.B(n_4971),
.Y(n_5218)
);

OR2x2_ASAP7_75t_L g5219 ( 
.A(n_5121),
.B(n_4979),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5142),
.Y(n_5220)
);

AND2x2_ASAP7_75t_L g5221 ( 
.A(n_5114),
.B(n_4960),
.Y(n_5221)
);

OAI21xp5_ASAP7_75t_L g5222 ( 
.A1(n_5111),
.A2(n_5013),
.B(n_772),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_5112),
.B(n_773),
.Y(n_5223)
);

INVx4_ASAP7_75t_L g5224 ( 
.A(n_5173),
.Y(n_5224)
);

OR2x2_ASAP7_75t_L g5225 ( 
.A(n_5124),
.B(n_1675),
.Y(n_5225)
);

AO21x1_ASAP7_75t_L g5226 ( 
.A1(n_5113),
.A2(n_774),
.B(n_775),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5151),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_5062),
.B(n_776),
.Y(n_5228)
);

NOR2x1_ASAP7_75t_L g5229 ( 
.A(n_5147),
.B(n_776),
.Y(n_5229)
);

OR2x2_ASAP7_75t_L g5230 ( 
.A(n_5126),
.B(n_1658),
.Y(n_5230)
);

INVx1_ASAP7_75t_SL g5231 ( 
.A(n_5129),
.Y(n_5231)
);

OR2x2_ASAP7_75t_L g5232 ( 
.A(n_5128),
.B(n_1659),
.Y(n_5232)
);

AND2x2_ASAP7_75t_L g5233 ( 
.A(n_5104),
.B(n_777),
.Y(n_5233)
);

INVxp67_ASAP7_75t_SL g5234 ( 
.A(n_5064),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_5072),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5073),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_5061),
.Y(n_5237)
);

HB1xp67_ASAP7_75t_L g5238 ( 
.A(n_5135),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_5079),
.Y(n_5239)
);

AND2x4_ASAP7_75t_SL g5240 ( 
.A(n_5100),
.B(n_1660),
.Y(n_5240)
);

OR2x2_ASAP7_75t_L g5241 ( 
.A(n_5136),
.B(n_1660),
.Y(n_5241)
);

CKINVDCx10_ASAP7_75t_R g5242 ( 
.A(n_5138),
.Y(n_5242)
);

AND2x2_ASAP7_75t_L g5243 ( 
.A(n_5131),
.B(n_5065),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5087),
.Y(n_5244)
);

AND2x2_ASAP7_75t_L g5245 ( 
.A(n_5117),
.B(n_778),
.Y(n_5245)
);

INVx2_ASAP7_75t_L g5246 ( 
.A(n_5144),
.Y(n_5246)
);

BUFx2_ASAP7_75t_L g5247 ( 
.A(n_5150),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5090),
.Y(n_5248)
);

HB1xp67_ASAP7_75t_L g5249 ( 
.A(n_5095),
.Y(n_5249)
);

INVx2_ASAP7_75t_L g5250 ( 
.A(n_5088),
.Y(n_5250)
);

OR2x2_ASAP7_75t_L g5251 ( 
.A(n_5076),
.B(n_1664),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5096),
.Y(n_5252)
);

AND2x2_ASAP7_75t_L g5253 ( 
.A(n_5145),
.B(n_5172),
.Y(n_5253)
);

AND2x2_ASAP7_75t_L g5254 ( 
.A(n_5137),
.B(n_780),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5132),
.B(n_781),
.Y(n_5255)
);

INVx1_ASAP7_75t_SL g5256 ( 
.A(n_5143),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_5070),
.B(n_782),
.Y(n_5257)
);

OAI221xp5_ASAP7_75t_L g5258 ( 
.A1(n_5106),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.C(n_787),
.Y(n_5258)
);

AND2x2_ASAP7_75t_L g5259 ( 
.A(n_5058),
.B(n_786),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_5068),
.B(n_788),
.Y(n_5260)
);

AND2x4_ASAP7_75t_L g5261 ( 
.A(n_5107),
.B(n_1655),
.Y(n_5261)
);

OR2x2_ASAP7_75t_L g5262 ( 
.A(n_5093),
.B(n_1655),
.Y(n_5262)
);

INVxp67_ASAP7_75t_SL g5263 ( 
.A(n_5089),
.Y(n_5263)
);

OR2x2_ASAP7_75t_L g5264 ( 
.A(n_5116),
.B(n_1656),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_5170),
.B(n_789),
.Y(n_5265)
);

AOI31xp33_ASAP7_75t_L g5266 ( 
.A1(n_5190),
.A2(n_5226),
.A3(n_5192),
.B(n_5188),
.Y(n_5266)
);

AND2x2_ASAP7_75t_L g5267 ( 
.A(n_5201),
.B(n_5140),
.Y(n_5267)
);

INVxp67_ASAP7_75t_SL g5268 ( 
.A(n_5176),
.Y(n_5268)
);

AND2x2_ASAP7_75t_L g5269 ( 
.A(n_5177),
.B(n_5141),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5178),
.Y(n_5270)
);

INVx2_ASAP7_75t_SL g5271 ( 
.A(n_5193),
.Y(n_5271)
);

NOR3xp33_ASAP7_75t_L g5272 ( 
.A(n_5184),
.B(n_5161),
.C(n_5130),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_L g5273 ( 
.A(n_5218),
.B(n_5171),
.Y(n_5273)
);

AND2x2_ASAP7_75t_L g5274 ( 
.A(n_5253),
.B(n_5148),
.Y(n_5274)
);

AND2x2_ASAP7_75t_L g5275 ( 
.A(n_5215),
.B(n_5154),
.Y(n_5275)
);

OR2x2_ASAP7_75t_L g5276 ( 
.A(n_5208),
.B(n_5156),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_5179),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5202),
.B(n_5198),
.Y(n_5278)
);

AND2x2_ASAP7_75t_L g5279 ( 
.A(n_5194),
.B(n_5159),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_SL g5280 ( 
.A(n_5209),
.B(n_5120),
.Y(n_5280)
);

OR2x2_ASAP7_75t_L g5281 ( 
.A(n_5189),
.B(n_5256),
.Y(n_5281)
);

AND2x2_ASAP7_75t_L g5282 ( 
.A(n_5224),
.B(n_5162),
.Y(n_5282)
);

NAND2xp5_ASAP7_75t_L g5283 ( 
.A(n_5216),
.B(n_5163),
.Y(n_5283)
);

NAND4xp25_ASAP7_75t_L g5284 ( 
.A(n_5214),
.B(n_5080),
.C(n_5105),
.D(n_5084),
.Y(n_5284)
);

INVx2_ASAP7_75t_L g5285 ( 
.A(n_5203),
.Y(n_5285)
);

INVx2_ASAP7_75t_SL g5286 ( 
.A(n_5240),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_5199),
.B(n_5164),
.Y(n_5287)
);

HB1xp67_ASAP7_75t_L g5288 ( 
.A(n_5213),
.Y(n_5288)
);

OR2x2_ASAP7_75t_L g5289 ( 
.A(n_5239),
.B(n_5165),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_5247),
.Y(n_5290)
);

OR2x2_ASAP7_75t_L g5291 ( 
.A(n_5237),
.B(n_5204),
.Y(n_5291)
);

INVxp67_ASAP7_75t_L g5292 ( 
.A(n_5229),
.Y(n_5292)
);

AND2x2_ASAP7_75t_L g5293 ( 
.A(n_5243),
.B(n_5160),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5219),
.Y(n_5294)
);

OR2x2_ASAP7_75t_L g5295 ( 
.A(n_5191),
.B(n_5115),
.Y(n_5295)
);

INVxp67_ASAP7_75t_L g5296 ( 
.A(n_5221),
.Y(n_5296)
);

INVx2_ASAP7_75t_L g5297 ( 
.A(n_5197),
.Y(n_5297)
);

HB1xp67_ASAP7_75t_L g5298 ( 
.A(n_5231),
.Y(n_5298)
);

AND3x1_ASAP7_75t_L g5299 ( 
.A(n_5186),
.B(n_5158),
.C(n_5146),
.Y(n_5299)
);

AND2x2_ASAP7_75t_L g5300 ( 
.A(n_5206),
.B(n_5094),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_5180),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_5249),
.Y(n_5302)
);

AND2x4_ASAP7_75t_L g5303 ( 
.A(n_5250),
.B(n_5108),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5234),
.B(n_5212),
.Y(n_5304)
);

AND2x4_ASAP7_75t_L g5305 ( 
.A(n_5195),
.B(n_5155),
.Y(n_5305)
);

AND2x2_ASAP7_75t_L g5306 ( 
.A(n_5263),
.B(n_790),
.Y(n_5306)
);

NAND2xp5_ASAP7_75t_L g5307 ( 
.A(n_5207),
.B(n_5123),
.Y(n_5307)
);

NOR2xp67_ASAP7_75t_L g5308 ( 
.A(n_5187),
.B(n_790),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_5225),
.Y(n_5309)
);

NAND2x1p5_ASAP7_75t_L g5310 ( 
.A(n_5261),
.B(n_5125),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_5230),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_5246),
.B(n_791),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_5183),
.B(n_791),
.Y(n_5313)
);

NAND2x1p5_ASAP7_75t_L g5314 ( 
.A(n_5232),
.B(n_793),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_5241),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_L g5316 ( 
.A(n_5217),
.B(n_792),
.Y(n_5316)
);

NAND2xp5_ASAP7_75t_L g5317 ( 
.A(n_5174),
.B(n_795),
.Y(n_5317)
);

AND2x2_ASAP7_75t_L g5318 ( 
.A(n_5175),
.B(n_795),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5264),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_5210),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_5238),
.B(n_796),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_5211),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_5220),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_5227),
.Y(n_5324)
);

INVxp67_ASAP7_75t_SL g5325 ( 
.A(n_5228),
.Y(n_5325)
);

NOR2xp33_ASAP7_75t_L g5326 ( 
.A(n_5242),
.B(n_5185),
.Y(n_5326)
);

AND2x2_ASAP7_75t_L g5327 ( 
.A(n_5259),
.B(n_798),
.Y(n_5327)
);

NOR2xp33_ASAP7_75t_L g5328 ( 
.A(n_5251),
.B(n_1671),
.Y(n_5328)
);

OR2x2_ASAP7_75t_L g5329 ( 
.A(n_5196),
.B(n_798),
.Y(n_5329)
);

AND2x2_ASAP7_75t_L g5330 ( 
.A(n_5255),
.B(n_800),
.Y(n_5330)
);

OR2x6_ASAP7_75t_L g5331 ( 
.A(n_5222),
.B(n_5245),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_5235),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_5254),
.B(n_801),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_5200),
.B(n_801),
.Y(n_5334)
);

OR2x2_ASAP7_75t_L g5335 ( 
.A(n_5205),
.B(n_803),
.Y(n_5335)
);

OR2x6_ASAP7_75t_L g5336 ( 
.A(n_5233),
.B(n_803),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_5236),
.Y(n_5337)
);

INVx1_ASAP7_75t_SL g5338 ( 
.A(n_5223),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_5260),
.B(n_804),
.Y(n_5339)
);

NOR4xp25_ASAP7_75t_L g5340 ( 
.A(n_5258),
.B(n_806),
.C(n_804),
.D(n_805),
.Y(n_5340)
);

OR2x2_ASAP7_75t_L g5341 ( 
.A(n_5262),
.B(n_805),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_5244),
.Y(n_5342)
);

NOR2xp33_ASAP7_75t_L g5343 ( 
.A(n_5257),
.B(n_1657),
.Y(n_5343)
);

OR2x2_ASAP7_75t_L g5344 ( 
.A(n_5248),
.B(n_807),
.Y(n_5344)
);

AND2x2_ASAP7_75t_L g5345 ( 
.A(n_5252),
.B(n_807),
.Y(n_5345)
);

INVxp67_ASAP7_75t_SL g5346 ( 
.A(n_5265),
.Y(n_5346)
);

AND2x2_ASAP7_75t_L g5347 ( 
.A(n_5182),
.B(n_808),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_5182),
.B(n_808),
.Y(n_5348)
);

INVx2_ASAP7_75t_L g5349 ( 
.A(n_5181),
.Y(n_5349)
);

INVx1_ASAP7_75t_SL g5350 ( 
.A(n_5188),
.Y(n_5350)
);

NAND3xp33_ASAP7_75t_SL g5351 ( 
.A(n_5280),
.B(n_809),
.C(n_810),
.Y(n_5351)
);

OAI21xp5_ASAP7_75t_L g5352 ( 
.A1(n_5266),
.A2(n_809),
.B(n_810),
.Y(n_5352)
);

AOI32xp33_ASAP7_75t_L g5353 ( 
.A1(n_5299),
.A2(n_813),
.A3(n_811),
.B1(n_812),
.B2(n_814),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_5298),
.B(n_5350),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5290),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5291),
.Y(n_5356)
);

OAI21xp33_ASAP7_75t_L g5357 ( 
.A1(n_5326),
.A2(n_817),
.B(n_818),
.Y(n_5357)
);

AND2x2_ASAP7_75t_L g5358 ( 
.A(n_5286),
.B(n_1653),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_5268),
.B(n_1654),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_5270),
.Y(n_5360)
);

NOR2xp33_ASAP7_75t_L g5361 ( 
.A(n_5292),
.B(n_1661),
.Y(n_5361)
);

INVxp67_ASAP7_75t_SL g5362 ( 
.A(n_5308),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5304),
.Y(n_5363)
);

A2O1A1Ixp33_ASAP7_75t_L g5364 ( 
.A1(n_5272),
.A2(n_824),
.B(n_822),
.C(n_823),
.Y(n_5364)
);

OAI22xp5_ASAP7_75t_L g5365 ( 
.A1(n_5310),
.A2(n_827),
.B1(n_828),
.B2(n_826),
.Y(n_5365)
);

NAND2xp5_ASAP7_75t_L g5366 ( 
.A(n_5349),
.B(n_5347),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_5348),
.B(n_825),
.Y(n_5367)
);

AOI22xp5_ASAP7_75t_L g5368 ( 
.A1(n_5284),
.A2(n_829),
.B1(n_827),
.B2(n_828),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_5345),
.Y(n_5369)
);

AOI222xp33_ASAP7_75t_L g5370 ( 
.A1(n_5307),
.A2(n_832),
.B1(n_835),
.B2(n_836),
.C1(n_831),
.C2(n_833),
.Y(n_5370)
);

AND2x2_ASAP7_75t_L g5371 ( 
.A(n_5271),
.B(n_1663),
.Y(n_5371)
);

AOI22xp5_ASAP7_75t_L g5372 ( 
.A1(n_5305),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_5372)
);

AOI22xp33_ASAP7_75t_L g5373 ( 
.A1(n_5285),
.A2(n_837),
.B1(n_833),
.B2(n_836),
.Y(n_5373)
);

AOI21xp33_ASAP7_75t_SL g5374 ( 
.A1(n_5340),
.A2(n_1676),
.B(n_838),
.Y(n_5374)
);

OAI21xp33_ASAP7_75t_L g5375 ( 
.A1(n_5273),
.A2(n_839),
.B(n_840),
.Y(n_5375)
);

OR2x2_ASAP7_75t_L g5376 ( 
.A(n_5338),
.B(n_840),
.Y(n_5376)
);

OAI21xp5_ASAP7_75t_SL g5377 ( 
.A1(n_5296),
.A2(n_5300),
.B(n_5313),
.Y(n_5377)
);

AOI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_5303),
.A2(n_844),
.B1(n_842),
.B2(n_843),
.Y(n_5378)
);

INVxp67_ASAP7_75t_L g5379 ( 
.A(n_5288),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_5281),
.Y(n_5380)
);

OAI22xp5_ASAP7_75t_L g5381 ( 
.A1(n_5295),
.A2(n_846),
.B1(n_847),
.B2(n_845),
.Y(n_5381)
);

AOI21xp5_ASAP7_75t_L g5382 ( 
.A1(n_5316),
.A2(n_847),
.B(n_848),
.Y(n_5382)
);

NAND2xp5_ASAP7_75t_L g5383 ( 
.A(n_5293),
.B(n_849),
.Y(n_5383)
);

INVx2_ASAP7_75t_L g5384 ( 
.A(n_5314),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5341),
.Y(n_5385)
);

OAI21xp5_ASAP7_75t_L g5386 ( 
.A1(n_5317),
.A2(n_850),
.B(n_851),
.Y(n_5386)
);

AOI22xp33_ASAP7_75t_SL g5387 ( 
.A1(n_5346),
.A2(n_1673),
.B1(n_853),
.B2(n_851),
.Y(n_5387)
);

NAND3xp33_ASAP7_75t_L g5388 ( 
.A(n_5277),
.B(n_5301),
.C(n_5302),
.Y(n_5388)
);

AND2x2_ASAP7_75t_L g5389 ( 
.A(n_5274),
.B(n_5331),
.Y(n_5389)
);

AOI22xp5_ASAP7_75t_L g5390 ( 
.A1(n_5297),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.Y(n_5390)
);

BUFx2_ASAP7_75t_L g5391 ( 
.A(n_5336),
.Y(n_5391)
);

OAI22xp5_ASAP7_75t_L g5392 ( 
.A1(n_5283),
.A2(n_855),
.B1(n_856),
.B2(n_854),
.Y(n_5392)
);

CKINVDCx20_ASAP7_75t_R g5393 ( 
.A(n_5336),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_5306),
.B(n_852),
.Y(n_5394)
);

AND2x2_ASAP7_75t_L g5395 ( 
.A(n_5275),
.B(n_1651),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_5344),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5282),
.Y(n_5397)
);

AND2x2_ASAP7_75t_L g5398 ( 
.A(n_5267),
.B(n_1652),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_5269),
.B(n_855),
.Y(n_5399)
);

OAI21xp33_ASAP7_75t_L g5400 ( 
.A1(n_5325),
.A2(n_857),
.B(n_858),
.Y(n_5400)
);

AO22x1_ASAP7_75t_L g5401 ( 
.A1(n_5294),
.A2(n_5319),
.B1(n_5311),
.B2(n_5315),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_L g5402 ( 
.A(n_5279),
.B(n_859),
.Y(n_5402)
);

AOI22xp5_ASAP7_75t_L g5403 ( 
.A1(n_5287),
.A2(n_861),
.B1(n_859),
.B2(n_860),
.Y(n_5403)
);

OR2x2_ASAP7_75t_L g5404 ( 
.A(n_5309),
.B(n_5320),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5321),
.Y(n_5405)
);

OAI22xp33_ASAP7_75t_L g5406 ( 
.A1(n_5276),
.A2(n_865),
.B1(n_863),
.B2(n_864),
.Y(n_5406)
);

INVxp67_ASAP7_75t_L g5407 ( 
.A(n_5318),
.Y(n_5407)
);

OAI22xp33_ASAP7_75t_L g5408 ( 
.A1(n_5334),
.A2(n_866),
.B1(n_864),
.B2(n_865),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_5328),
.B(n_867),
.Y(n_5409)
);

AOI22xp5_ASAP7_75t_L g5410 ( 
.A1(n_5343),
.A2(n_869),
.B1(n_867),
.B2(n_868),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5329),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5335),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5289),
.Y(n_5413)
);

AND2x2_ASAP7_75t_L g5414 ( 
.A(n_5327),
.B(n_1647),
.Y(n_5414)
);

AND2x2_ASAP7_75t_SL g5415 ( 
.A(n_5312),
.B(n_870),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5330),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5333),
.Y(n_5417)
);

OAI221xp5_ASAP7_75t_SL g5418 ( 
.A1(n_5322),
.A2(n_874),
.B1(n_872),
.B2(n_873),
.C(n_875),
.Y(n_5418)
);

AOI222xp33_ASAP7_75t_L g5419 ( 
.A1(n_5332),
.A2(n_874),
.B1(n_876),
.B2(n_877),
.C1(n_873),
.C2(n_875),
.Y(n_5419)
);

AND2x4_ASAP7_75t_L g5420 ( 
.A(n_5323),
.B(n_5324),
.Y(n_5420)
);

AND2x2_ASAP7_75t_L g5421 ( 
.A(n_5339),
.B(n_1657),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_5337),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5342),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5290),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5290),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5278),
.Y(n_5426)
);

AND2x2_ASAP7_75t_L g5427 ( 
.A(n_5278),
.B(n_1642),
.Y(n_5427)
);

HB1xp67_ASAP7_75t_L g5428 ( 
.A(n_5308),
.Y(n_5428)
);

NAND2xp5_ASAP7_75t_L g5429 ( 
.A(n_5298),
.B(n_878),
.Y(n_5429)
);

O2A1O1Ixp33_ASAP7_75t_L g5430 ( 
.A1(n_5266),
.A2(n_881),
.B(n_879),
.C(n_880),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_5278),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_5362),
.B(n_883),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_5428),
.Y(n_5433)
);

NOR2x1p5_ASAP7_75t_SL g5434 ( 
.A(n_5355),
.B(n_884),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5424),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_5425),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5389),
.B(n_887),
.Y(n_5437)
);

INVxp67_ASAP7_75t_L g5438 ( 
.A(n_5391),
.Y(n_5438)
);

AOI222xp33_ASAP7_75t_L g5439 ( 
.A1(n_5401),
.A2(n_910),
.B1(n_893),
.B2(n_918),
.C1(n_903),
.C2(n_888),
.Y(n_5439)
);

AOI21xp5_ASAP7_75t_L g5440 ( 
.A1(n_5430),
.A2(n_889),
.B(n_890),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_L g5441 ( 
.A(n_5379),
.B(n_891),
.Y(n_5441)
);

AND2x2_ASAP7_75t_L g5442 ( 
.A(n_5426),
.B(n_891),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5414),
.Y(n_5443)
);

AOI21xp33_ASAP7_75t_L g5444 ( 
.A1(n_5380),
.A2(n_1650),
.B(n_1648),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5358),
.Y(n_5445)
);

OAI22xp5_ASAP7_75t_L g5446 ( 
.A1(n_5368),
.A2(n_897),
.B1(n_894),
.B2(n_895),
.Y(n_5446)
);

NOR2xp33_ASAP7_75t_L g5447 ( 
.A(n_5357),
.B(n_898),
.Y(n_5447)
);

INVx1_ASAP7_75t_SL g5448 ( 
.A(n_5359),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5376),
.Y(n_5449)
);

AOI21x1_ASAP7_75t_L g5450 ( 
.A1(n_5382),
.A2(n_899),
.B(n_900),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_5431),
.B(n_900),
.Y(n_5451)
);

AOI31xp33_ASAP7_75t_SL g5452 ( 
.A1(n_5407),
.A2(n_906),
.A3(n_904),
.B(n_905),
.Y(n_5452)
);

NAND2xp5_ASAP7_75t_L g5453 ( 
.A(n_5353),
.B(n_5415),
.Y(n_5453)
);

INVx2_ASAP7_75t_SL g5454 ( 
.A(n_5371),
.Y(n_5454)
);

INVx2_ASAP7_75t_L g5455 ( 
.A(n_5397),
.Y(n_5455)
);

OAI322xp33_ASAP7_75t_L g5456 ( 
.A1(n_5388),
.A2(n_911),
.A3(n_909),
.B1(n_907),
.B2(n_904),
.C1(n_905),
.C2(n_908),
.Y(n_5456)
);

OAI31xp33_ASAP7_75t_L g5457 ( 
.A1(n_5364),
.A2(n_912),
.A3(n_907),
.B(n_909),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_5429),
.Y(n_5458)
);

OAI321xp33_ASAP7_75t_L g5459 ( 
.A1(n_5356),
.A2(n_916),
.A3(n_918),
.B1(n_913),
.B2(n_915),
.C(n_917),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5404),
.Y(n_5460)
);

AOI221xp5_ASAP7_75t_L g5461 ( 
.A1(n_5377),
.A2(n_934),
.B1(n_943),
.B2(n_924),
.C(n_913),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5398),
.Y(n_5462)
);

OAI21xp33_ASAP7_75t_L g5463 ( 
.A1(n_5366),
.A2(n_920),
.B(n_921),
.Y(n_5463)
);

NAND2xp5_ASAP7_75t_SL g5464 ( 
.A(n_5384),
.B(n_921),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5416),
.Y(n_5465)
);

INVx2_ASAP7_75t_L g5466 ( 
.A(n_5427),
.Y(n_5466)
);

NOR2xp33_ASAP7_75t_SL g5467 ( 
.A(n_5418),
.B(n_922),
.Y(n_5467)
);

BUFx2_ASAP7_75t_L g5468 ( 
.A(n_5395),
.Y(n_5468)
);

NAND3xp33_ASAP7_75t_L g5469 ( 
.A(n_5370),
.B(n_923),
.C(n_924),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_5417),
.Y(n_5470)
);

AOI221xp5_ASAP7_75t_L g5471 ( 
.A1(n_5360),
.A2(n_944),
.B1(n_950),
.B2(n_935),
.C(n_925),
.Y(n_5471)
);

OAI22xp5_ASAP7_75t_L g5472 ( 
.A1(n_5372),
.A2(n_928),
.B1(n_926),
.B2(n_927),
.Y(n_5472)
);

OAI31xp33_ASAP7_75t_L g5473 ( 
.A1(n_5408),
.A2(n_931),
.A3(n_929),
.B(n_930),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5367),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5369),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5385),
.Y(n_5476)
);

OAI21xp5_ASAP7_75t_L g5477 ( 
.A1(n_5361),
.A2(n_931),
.B(n_934),
.Y(n_5477)
);

NAND2xp5_ASAP7_75t_L g5478 ( 
.A(n_5396),
.B(n_936),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5399),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5402),
.Y(n_5480)
);

NAND2xp33_ASAP7_75t_SL g5481 ( 
.A(n_5413),
.B(n_937),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5411),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_5412),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_5421),
.B(n_936),
.Y(n_5484)
);

INVx2_ASAP7_75t_SL g5485 ( 
.A(n_5420),
.Y(n_5485)
);

OAI221xp5_ASAP7_75t_L g5486 ( 
.A1(n_5375),
.A2(n_940),
.B1(n_937),
.B2(n_938),
.C(n_941),
.Y(n_5486)
);

NOR3xp33_ASAP7_75t_L g5487 ( 
.A(n_5363),
.B(n_938),
.C(n_942),
.Y(n_5487)
);

INVxp67_ASAP7_75t_L g5488 ( 
.A(n_5394),
.Y(n_5488)
);

INVxp67_ASAP7_75t_L g5489 ( 
.A(n_5383),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_5387),
.B(n_943),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5420),
.Y(n_5491)
);

AOI21xp33_ASAP7_75t_L g5492 ( 
.A1(n_5405),
.A2(n_1639),
.B(n_1638),
.Y(n_5492)
);

NAND2xp5_ASAP7_75t_L g5493 ( 
.A(n_5378),
.B(n_947),
.Y(n_5493)
);

AND2x2_ASAP7_75t_L g5494 ( 
.A(n_5386),
.B(n_948),
.Y(n_5494)
);

INVxp67_ASAP7_75t_L g5495 ( 
.A(n_5365),
.Y(n_5495)
);

INVx1_ASAP7_75t_SL g5496 ( 
.A(n_5409),
.Y(n_5496)
);

OAI22xp33_ASAP7_75t_L g5497 ( 
.A1(n_5403),
.A2(n_954),
.B1(n_951),
.B2(n_952),
.Y(n_5497)
);

NAND2xp5_ASAP7_75t_L g5498 ( 
.A(n_5406),
.B(n_952),
.Y(n_5498)
);

NAND2x1_ASAP7_75t_L g5499 ( 
.A(n_5422),
.B(n_1643),
.Y(n_5499)
);

AND2x2_ASAP7_75t_L g5500 ( 
.A(n_5423),
.B(n_955),
.Y(n_5500)
);

AND2x2_ASAP7_75t_L g5501 ( 
.A(n_5400),
.B(n_957),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_SL g5502 ( 
.A(n_5381),
.B(n_5419),
.Y(n_5502)
);

NAND2xp5_ASAP7_75t_L g5503 ( 
.A(n_5392),
.B(n_5410),
.Y(n_5503)
);

AOI21xp33_ASAP7_75t_L g5504 ( 
.A1(n_5373),
.A2(n_1647),
.B(n_1646),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_5390),
.B(n_958),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_5389),
.B(n_959),
.Y(n_5506)
);

OAI211xp5_ASAP7_75t_L g5507 ( 
.A1(n_5352),
.A2(n_968),
.B(n_965),
.C(n_967),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_5362),
.B(n_967),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5428),
.Y(n_5509)
);

NAND2xp5_ASAP7_75t_L g5510 ( 
.A(n_5362),
.B(n_969),
.Y(n_5510)
);

NOR2xp33_ASAP7_75t_L g5511 ( 
.A(n_5354),
.B(n_972),
.Y(n_5511)
);

BUFx2_ASAP7_75t_L g5512 ( 
.A(n_5362),
.Y(n_5512)
);

OAI322xp33_ASAP7_75t_L g5513 ( 
.A1(n_5374),
.A2(n_978),
.A3(n_977),
.B1(n_975),
.B2(n_973),
.C1(n_974),
.C2(n_976),
.Y(n_5513)
);

OAI221xp5_ASAP7_75t_L g5514 ( 
.A1(n_5352),
.A2(n_975),
.B1(n_973),
.B2(n_974),
.C(n_976),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_5362),
.B(n_979),
.Y(n_5515)
);

AOI221xp5_ASAP7_75t_L g5516 ( 
.A1(n_5352),
.A2(n_997),
.B1(n_1005),
.B2(n_987),
.C(n_980),
.Y(n_5516)
);

NOR2x1_ASAP7_75t_L g5517 ( 
.A(n_5351),
.B(n_981),
.Y(n_5517)
);

OAI211xp5_ASAP7_75t_SL g5518 ( 
.A1(n_5352),
.A2(n_984),
.B(n_982),
.C(n_983),
.Y(n_5518)
);

INVx2_ASAP7_75t_L g5519 ( 
.A(n_5393),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5428),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_5393),
.Y(n_5521)
);

AOI21xp33_ASAP7_75t_L g5522 ( 
.A1(n_5362),
.A2(n_1641),
.B(n_1640),
.Y(n_5522)
);

AOI21xp33_ASAP7_75t_L g5523 ( 
.A1(n_5362),
.A2(n_1645),
.B(n_1644),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5393),
.Y(n_5524)
);

AOI22xp5_ASAP7_75t_L g5525 ( 
.A1(n_5393),
.A2(n_988),
.B1(n_985),
.B2(n_986),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5428),
.Y(n_5526)
);

AOI211xp5_ASAP7_75t_L g5527 ( 
.A1(n_5374),
.A2(n_989),
.B(n_985),
.C(n_986),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5428),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_5428),
.Y(n_5529)
);

NAND2xp5_ASAP7_75t_L g5530 ( 
.A(n_5362),
.B(n_990),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5428),
.Y(n_5531)
);

NAND2xp5_ASAP7_75t_L g5532 ( 
.A(n_5362),
.B(n_991),
.Y(n_5532)
);

OAI322xp33_ASAP7_75t_L g5533 ( 
.A1(n_5374),
.A2(n_1000),
.A3(n_999),
.B1(n_996),
.B2(n_992),
.C1(n_993),
.C2(n_998),
.Y(n_5533)
);

OAI21xp33_ASAP7_75t_SL g5534 ( 
.A1(n_5352),
.A2(n_992),
.B(n_996),
.Y(n_5534)
);

AOI211xp5_ASAP7_75t_L g5535 ( 
.A1(n_5374),
.A2(n_1002),
.B(n_999),
.C(n_1001),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5362),
.B(n_1001),
.Y(n_5536)
);

NOR2xp33_ASAP7_75t_L g5537 ( 
.A(n_5354),
.B(n_1006),
.Y(n_5537)
);

INVx1_ASAP7_75t_SL g5538 ( 
.A(n_5393),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_5428),
.Y(n_5539)
);

OAI322xp33_ASAP7_75t_L g5540 ( 
.A1(n_5374),
.A2(n_1014),
.A3(n_1013),
.B1(n_1011),
.B2(n_1009),
.C1(n_1010),
.C2(n_1012),
.Y(n_5540)
);

NOR2xp33_ASAP7_75t_L g5541 ( 
.A(n_5354),
.B(n_1013),
.Y(n_5541)
);

INVx1_ASAP7_75t_L g5542 ( 
.A(n_5428),
.Y(n_5542)
);

NOR2xp67_ASAP7_75t_L g5543 ( 
.A(n_5485),
.B(n_1017),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5512),
.Y(n_5544)
);

AND2x2_ASAP7_75t_L g5545 ( 
.A(n_5538),
.B(n_5519),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5468),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5433),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_5509),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_5521),
.B(n_1018),
.Y(n_5549)
);

OR2x2_ASAP7_75t_L g5550 ( 
.A(n_5448),
.B(n_1018),
.Y(n_5550)
);

AOI221xp5_ASAP7_75t_L g5551 ( 
.A1(n_5502),
.A2(n_1664),
.B1(n_1663),
.B2(n_1646),
.C(n_1022),
.Y(n_5551)
);

AND2x2_ASAP7_75t_L g5552 ( 
.A(n_5524),
.B(n_1019),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5520),
.Y(n_5553)
);

NAND3xp33_ASAP7_75t_L g5554 ( 
.A(n_5439),
.B(n_1019),
.C(n_1020),
.Y(n_5554)
);

OAI22xp33_ASAP7_75t_SL g5555 ( 
.A1(n_5467),
.A2(n_5491),
.B1(n_5438),
.B2(n_5453),
.Y(n_5555)
);

AND2x2_ASAP7_75t_L g5556 ( 
.A(n_5437),
.B(n_5506),
.Y(n_5556)
);

XNOR2xp5_ASAP7_75t_L g5557 ( 
.A(n_5527),
.B(n_1023),
.Y(n_5557)
);

OAI22xp5_ASAP7_75t_L g5558 ( 
.A1(n_5469),
.A2(n_1026),
.B1(n_1024),
.B2(n_1025),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5526),
.Y(n_5559)
);

CKINVDCx16_ASAP7_75t_R g5560 ( 
.A(n_5481),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5528),
.Y(n_5561)
);

AND2x4_ASAP7_75t_L g5562 ( 
.A(n_5434),
.B(n_1637),
.Y(n_5562)
);

OAI32xp33_ASAP7_75t_L g5563 ( 
.A1(n_5534),
.A2(n_1040),
.A3(n_1047),
.B1(n_1035),
.B2(n_1028),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5529),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5531),
.Y(n_5565)
);

NOR2xp33_ASAP7_75t_L g5566 ( 
.A(n_5513),
.B(n_1029),
.Y(n_5566)
);

AND2x2_ASAP7_75t_L g5567 ( 
.A(n_5466),
.B(n_1030),
.Y(n_5567)
);

INVx2_ASAP7_75t_SL g5568 ( 
.A(n_5499),
.Y(n_5568)
);

AND2x2_ASAP7_75t_L g5569 ( 
.A(n_5454),
.B(n_1030),
.Y(n_5569)
);

NAND2xp5_ASAP7_75t_L g5570 ( 
.A(n_5539),
.B(n_1031),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5542),
.Y(n_5571)
);

NOR2xp33_ASAP7_75t_L g5572 ( 
.A(n_5533),
.B(n_1031),
.Y(n_5572)
);

AND2x2_ASAP7_75t_L g5573 ( 
.A(n_5445),
.B(n_1033),
.Y(n_5573)
);

OAI221xp5_ASAP7_75t_L g5574 ( 
.A1(n_5457),
.A2(n_1632),
.B1(n_1633),
.B2(n_1628),
.C(n_1626),
.Y(n_5574)
);

O2A1O1Ixp33_ASAP7_75t_SL g5575 ( 
.A1(n_5535),
.A2(n_1036),
.B(n_1034),
.C(n_1035),
.Y(n_5575)
);

NOR2xp33_ASAP7_75t_L g5576 ( 
.A(n_5540),
.B(n_1034),
.Y(n_5576)
);

AND2x4_ASAP7_75t_L g5577 ( 
.A(n_5460),
.B(n_1635),
.Y(n_5577)
);

OAI31xp33_ASAP7_75t_L g5578 ( 
.A1(n_5507),
.A2(n_1039),
.A3(n_1037),
.B(n_1038),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5432),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5508),
.Y(n_5580)
);

AND2x2_ASAP7_75t_L g5581 ( 
.A(n_5443),
.B(n_1042),
.Y(n_5581)
);

OAI32xp33_ASAP7_75t_L g5582 ( 
.A1(n_5503),
.A2(n_1058),
.A3(n_1061),
.B1(n_1049),
.B2(n_1043),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5510),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_5515),
.Y(n_5584)
);

NOR2x1_ASAP7_75t_L g5585 ( 
.A(n_5452),
.B(n_1046),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5462),
.B(n_1048),
.Y(n_5586)
);

OAI21xp5_ASAP7_75t_L g5587 ( 
.A1(n_5440),
.A2(n_1051),
.B(n_1050),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_SL g5588 ( 
.A(n_5517),
.B(n_1049),
.Y(n_5588)
);

AOI22xp33_ASAP7_75t_L g5589 ( 
.A1(n_5474),
.A2(n_5480),
.B1(n_5479),
.B2(n_5495),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5530),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5532),
.Y(n_5591)
);

OAI322xp33_ASAP7_75t_L g5592 ( 
.A1(n_5435),
.A2(n_1058),
.A3(n_1056),
.B1(n_1054),
.B2(n_1052),
.C1(n_1053),
.C2(n_1055),
.Y(n_5592)
);

AOI221xp5_ASAP7_75t_L g5593 ( 
.A1(n_5436),
.A2(n_1628),
.B1(n_1634),
.B2(n_1621),
.C(n_1620),
.Y(n_5593)
);

NAND2x1p5_ASAP7_75t_L g5594 ( 
.A(n_5464),
.B(n_1059),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5536),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_5442),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_5484),
.Y(n_5597)
);

AOI21xp33_ASAP7_75t_SL g5598 ( 
.A1(n_5449),
.A2(n_1613),
.B(n_1612),
.Y(n_5598)
);

AOI211xp5_ASAP7_75t_SL g5599 ( 
.A1(n_5476),
.A2(n_1071),
.B(n_1081),
.C(n_1062),
.Y(n_5599)
);

NAND3xp33_ASAP7_75t_L g5600 ( 
.A(n_5461),
.B(n_1062),
.C(n_1063),
.Y(n_5600)
);

AOI22xp5_ASAP7_75t_L g5601 ( 
.A1(n_5511),
.A2(n_5537),
.B1(n_5541),
.B2(n_5455),
.Y(n_5601)
);

AOI221xp5_ASAP7_75t_L g5602 ( 
.A1(n_5456),
.A2(n_1635),
.B1(n_1636),
.B2(n_1621),
.C(n_1618),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5441),
.Y(n_5603)
);

AOI22xp5_ASAP7_75t_L g5604 ( 
.A1(n_5470),
.A2(n_5518),
.B1(n_5496),
.B2(n_5487),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5500),
.Y(n_5605)
);

OAI32xp33_ASAP7_75t_L g5606 ( 
.A1(n_5490),
.A2(n_1086),
.A3(n_1089),
.B1(n_1080),
.B2(n_1068),
.Y(n_5606)
);

NAND2xp5_ASAP7_75t_L g5607 ( 
.A(n_5494),
.B(n_1068),
.Y(n_5607)
);

NOR2xp33_ASAP7_75t_L g5608 ( 
.A(n_5463),
.B(n_1070),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_L g5609 ( 
.A(n_5465),
.B(n_1070),
.Y(n_5609)
);

A2O1A1Ixp33_ASAP7_75t_L g5610 ( 
.A1(n_5459),
.A2(n_1075),
.B(n_1073),
.C(n_1074),
.Y(n_5610)
);

INVxp67_ASAP7_75t_L g5611 ( 
.A(n_5447),
.Y(n_5611)
);

NAND3xp33_ASAP7_75t_L g5612 ( 
.A(n_5482),
.B(n_5483),
.C(n_5516),
.Y(n_5612)
);

AOI22xp5_ASAP7_75t_L g5613 ( 
.A1(n_5489),
.A2(n_1610),
.B1(n_1611),
.B2(n_1609),
.Y(n_5613)
);

OR2x2_ASAP7_75t_L g5614 ( 
.A(n_5451),
.B(n_1075),
.Y(n_5614)
);

BUFx3_ASAP7_75t_L g5615 ( 
.A(n_5475),
.Y(n_5615)
);

OAI21xp33_ASAP7_75t_L g5616 ( 
.A1(n_5488),
.A2(n_1076),
.B(n_1077),
.Y(n_5616)
);

OAI32xp33_ASAP7_75t_L g5617 ( 
.A1(n_5498),
.A2(n_1089),
.A3(n_1097),
.B1(n_1086),
.B2(n_1078),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_5478),
.Y(n_5618)
);

NAND2xp5_ASAP7_75t_L g5619 ( 
.A(n_5473),
.B(n_5501),
.Y(n_5619)
);

OAI221xp5_ASAP7_75t_L g5620 ( 
.A1(n_5504),
.A2(n_5471),
.B1(n_5514),
.B2(n_5477),
.C(n_5458),
.Y(n_5620)
);

AND2x2_ASAP7_75t_L g5621 ( 
.A(n_5450),
.B(n_1087),
.Y(n_5621)
);

AOI22xp33_ASAP7_75t_L g5622 ( 
.A1(n_5545),
.A2(n_5446),
.B1(n_5486),
.B2(n_5522),
.Y(n_5622)
);

AOI211xp5_ASAP7_75t_SL g5623 ( 
.A1(n_5555),
.A2(n_5523),
.B(n_5444),
.C(n_5497),
.Y(n_5623)
);

AOI221x1_ASAP7_75t_L g5624 ( 
.A1(n_5544),
.A2(n_5492),
.B1(n_5493),
.B2(n_5472),
.C(n_5505),
.Y(n_5624)
);

AND2x2_ASAP7_75t_L g5625 ( 
.A(n_5556),
.B(n_5525),
.Y(n_5625)
);

AOI22xp33_ASAP7_75t_L g5626 ( 
.A1(n_5546),
.A2(n_1091),
.B1(n_1088),
.B2(n_1090),
.Y(n_5626)
);

AOI221xp5_ASAP7_75t_L g5627 ( 
.A1(n_5612),
.A2(n_1095),
.B1(n_1092),
.B2(n_1093),
.C(n_1096),
.Y(n_5627)
);

OAI211xp5_ASAP7_75t_L g5628 ( 
.A1(n_5604),
.A2(n_1104),
.B(n_1101),
.C(n_1103),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5543),
.Y(n_5629)
);

OAI211xp5_ASAP7_75t_SL g5630 ( 
.A1(n_5601),
.A2(n_1105),
.B(n_1103),
.C(n_1104),
.Y(n_5630)
);

OAI221xp5_ASAP7_75t_SL g5631 ( 
.A1(n_5578),
.A2(n_1604),
.B1(n_1605),
.B2(n_1603),
.C(n_1602),
.Y(n_5631)
);

O2A1O1Ixp33_ASAP7_75t_L g5632 ( 
.A1(n_5610),
.A2(n_1111),
.B(n_1109),
.C(n_1110),
.Y(n_5632)
);

AOI221xp5_ASAP7_75t_L g5633 ( 
.A1(n_5620),
.A2(n_1112),
.B1(n_1110),
.B2(n_1111),
.C(n_1113),
.Y(n_5633)
);

NOR2xp33_ASAP7_75t_L g5634 ( 
.A(n_5568),
.B(n_1112),
.Y(n_5634)
);

AOI221x1_ASAP7_75t_L g5635 ( 
.A1(n_5558),
.A2(n_1116),
.B1(n_1113),
.B2(n_1115),
.C(n_1117),
.Y(n_5635)
);

NAND2xp5_ASAP7_75t_SL g5636 ( 
.A(n_5585),
.B(n_1115),
.Y(n_5636)
);

XNOR2xp5_ASAP7_75t_L g5637 ( 
.A(n_5557),
.B(n_1116),
.Y(n_5637)
);

O2A1O1Ixp33_ASAP7_75t_SL g5638 ( 
.A1(n_5588),
.A2(n_1120),
.B(n_1118),
.C(n_1119),
.Y(n_5638)
);

NAND4xp25_ASAP7_75t_L g5639 ( 
.A(n_5619),
.B(n_1122),
.C(n_1119),
.D(n_1121),
.Y(n_5639)
);

AOI221xp5_ASAP7_75t_L g5640 ( 
.A1(n_5554),
.A2(n_1125),
.B1(n_1121),
.B2(n_1122),
.C(n_1126),
.Y(n_5640)
);

OAI21xp33_ASAP7_75t_L g5641 ( 
.A1(n_5611),
.A2(n_1128),
.B(n_1129),
.Y(n_5641)
);

AOI211xp5_ASAP7_75t_L g5642 ( 
.A1(n_5563),
.A2(n_1637),
.B(n_1617),
.C(n_1132),
.Y(n_5642)
);

NAND4xp75_ASAP7_75t_L g5643 ( 
.A(n_5547),
.B(n_1133),
.C(n_1130),
.D(n_1131),
.Y(n_5643)
);

INVxp67_ASAP7_75t_SL g5644 ( 
.A(n_5594),
.Y(n_5644)
);

NOR4xp25_ASAP7_75t_SL g5645 ( 
.A(n_5575),
.B(n_1140),
.C(n_1138),
.D(n_1139),
.Y(n_5645)
);

NOR2xp33_ASAP7_75t_L g5646 ( 
.A(n_5616),
.B(n_1138),
.Y(n_5646)
);

OAI211xp5_ASAP7_75t_L g5647 ( 
.A1(n_5602),
.A2(n_1144),
.B(n_1142),
.C(n_1143),
.Y(n_5647)
);

AOI221xp5_ASAP7_75t_L g5648 ( 
.A1(n_5548),
.A2(n_1146),
.B1(n_1142),
.B2(n_1145),
.C(n_1147),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5599),
.B(n_1147),
.Y(n_5649)
);

AOI21xp5_ASAP7_75t_L g5650 ( 
.A1(n_5587),
.A2(n_1148),
.B(n_1149),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5569),
.Y(n_5651)
);

AOI22xp5_ASAP7_75t_L g5652 ( 
.A1(n_5566),
.A2(n_1151),
.B1(n_1149),
.B2(n_1150),
.Y(n_5652)
);

AOI322xp5_ASAP7_75t_L g5653 ( 
.A1(n_5572),
.A2(n_5576),
.A3(n_5551),
.B1(n_5553),
.B2(n_5559),
.C1(n_5564),
.C2(n_5561),
.Y(n_5653)
);

NAND2xp5_ASAP7_75t_L g5654 ( 
.A(n_5552),
.B(n_1152),
.Y(n_5654)
);

O2A1O1Ixp33_ASAP7_75t_L g5655 ( 
.A1(n_5582),
.A2(n_1157),
.B(n_1155),
.C(n_1156),
.Y(n_5655)
);

AOI221xp5_ASAP7_75t_L g5656 ( 
.A1(n_5565),
.A2(n_1161),
.B1(n_1158),
.B2(n_1159),
.C(n_1162),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_5577),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5550),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5581),
.Y(n_5659)
);

AOI221xp5_ASAP7_75t_L g5660 ( 
.A1(n_5571),
.A2(n_1168),
.B1(n_1166),
.B2(n_1167),
.C(n_1169),
.Y(n_5660)
);

AOI221xp5_ASAP7_75t_L g5661 ( 
.A1(n_5606),
.A2(n_1170),
.B1(n_1167),
.B2(n_1168),
.C(n_1171),
.Y(n_5661)
);

AOI211xp5_ASAP7_75t_L g5662 ( 
.A1(n_5574),
.A2(n_1614),
.B(n_1608),
.C(n_1172),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_5586),
.Y(n_5663)
);

AOI311xp33_ASAP7_75t_L g5664 ( 
.A1(n_5605),
.A2(n_1174),
.A3(n_1170),
.B(n_1173),
.C(n_1175),
.Y(n_5664)
);

NOR3xp33_ASAP7_75t_L g5665 ( 
.A(n_5579),
.B(n_1175),
.C(n_1176),
.Y(n_5665)
);

OR2x2_ASAP7_75t_L g5666 ( 
.A(n_5596),
.B(n_5570),
.Y(n_5666)
);

AOI32xp33_ASAP7_75t_L g5667 ( 
.A1(n_5615),
.A2(n_1179),
.A3(n_1177),
.B1(n_1178),
.B2(n_1180),
.Y(n_5667)
);

AOI221xp5_ASAP7_75t_L g5668 ( 
.A1(n_5600),
.A2(n_1184),
.B1(n_1182),
.B2(n_1183),
.C(n_1185),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5567),
.Y(n_5669)
);

AOI21xp5_ASAP7_75t_L g5670 ( 
.A1(n_5607),
.A2(n_5621),
.B(n_5549),
.Y(n_5670)
);

AOI322xp5_ASAP7_75t_L g5671 ( 
.A1(n_5608),
.A2(n_1614),
.A3(n_1188),
.B1(n_1185),
.B2(n_1187),
.C1(n_1183),
.C2(n_1184),
.Y(n_5671)
);

HB1xp67_ASAP7_75t_L g5672 ( 
.A(n_5577),
.Y(n_5672)
);

AOI221xp5_ASAP7_75t_L g5673 ( 
.A1(n_5617),
.A2(n_1193),
.B1(n_1191),
.B2(n_1192),
.C(n_1194),
.Y(n_5673)
);

NAND2xp5_ASAP7_75t_L g5674 ( 
.A(n_5598),
.B(n_1191),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5573),
.Y(n_5675)
);

OAI21xp33_ASAP7_75t_L g5676 ( 
.A1(n_5597),
.A2(n_1195),
.B(n_1196),
.Y(n_5676)
);

AOI211x1_ASAP7_75t_L g5677 ( 
.A1(n_5609),
.A2(n_1202),
.B(n_1200),
.C(n_1201),
.Y(n_5677)
);

NOR3xp33_ASAP7_75t_L g5678 ( 
.A(n_5580),
.B(n_1202),
.C(n_1203),
.Y(n_5678)
);

NAND4xp25_ASAP7_75t_SL g5679 ( 
.A(n_5583),
.B(n_1205),
.C(n_1203),
.D(n_1204),
.Y(n_5679)
);

AOI211xp5_ASAP7_75t_L g5680 ( 
.A1(n_5592),
.A2(n_1598),
.B(n_1601),
.C(n_1597),
.Y(n_5680)
);

OAI221xp5_ASAP7_75t_L g5681 ( 
.A1(n_5584),
.A2(n_1208),
.B1(n_1206),
.B2(n_1207),
.C(n_1209),
.Y(n_5681)
);

NOR3xp33_ASAP7_75t_L g5682 ( 
.A(n_5590),
.B(n_1212),
.C(n_1213),
.Y(n_5682)
);

OAI221xp5_ASAP7_75t_L g5683 ( 
.A1(n_5591),
.A2(n_5595),
.B1(n_5603),
.B2(n_5618),
.C(n_5593),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5614),
.Y(n_5684)
);

OAI211xp5_ASAP7_75t_SL g5685 ( 
.A1(n_5613),
.A2(n_1215),
.B(n_1213),
.C(n_1214),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5543),
.Y(n_5686)
);

OAI211xp5_ASAP7_75t_SL g5687 ( 
.A1(n_5589),
.A2(n_1223),
.B(n_1221),
.C(n_1222),
.Y(n_5687)
);

OAI22xp5_ASAP7_75t_L g5688 ( 
.A1(n_5560),
.A2(n_1223),
.B1(n_1221),
.B2(n_1222),
.Y(n_5688)
);

AOI221x1_ASAP7_75t_L g5689 ( 
.A1(n_5555),
.A2(n_1232),
.B1(n_1230),
.B2(n_1231),
.C(n_1233),
.Y(n_5689)
);

NOR2xp33_ASAP7_75t_L g5690 ( 
.A(n_5560),
.B(n_1236),
.Y(n_5690)
);

AOI21xp5_ASAP7_75t_L g5691 ( 
.A1(n_5562),
.A2(n_1239),
.B(n_1240),
.Y(n_5691)
);

OAI21xp33_ASAP7_75t_L g5692 ( 
.A1(n_5545),
.A2(n_1243),
.B(n_1244),
.Y(n_5692)
);

AOI211xp5_ASAP7_75t_L g5693 ( 
.A1(n_5555),
.A2(n_1594),
.B(n_1595),
.C(n_1593),
.Y(n_5693)
);

AOI211xp5_ASAP7_75t_L g5694 ( 
.A1(n_5555),
.A2(n_1596),
.B(n_1606),
.C(n_1595),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_SL g5695 ( 
.A(n_5562),
.B(n_1247),
.Y(n_5695)
);

AOI21xp5_ASAP7_75t_L g5696 ( 
.A1(n_5562),
.A2(n_1248),
.B(n_1249),
.Y(n_5696)
);

NAND2xp5_ASAP7_75t_L g5697 ( 
.A(n_5562),
.B(n_1250),
.Y(n_5697)
);

NOR2xp33_ASAP7_75t_L g5698 ( 
.A(n_5560),
.B(n_1251),
.Y(n_5698)
);

OAI22xp5_ASAP7_75t_L g5699 ( 
.A1(n_5622),
.A2(n_1257),
.B1(n_1255),
.B2(n_1256),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_L g5700 ( 
.A(n_5672),
.B(n_1258),
.Y(n_5700)
);

AOI21xp5_ASAP7_75t_L g5701 ( 
.A1(n_5695),
.A2(n_1261),
.B(n_1263),
.Y(n_5701)
);

NAND5xp2_ASAP7_75t_L g5702 ( 
.A(n_5653),
.B(n_1266),
.C(n_1264),
.D(n_1265),
.E(n_1267),
.Y(n_5702)
);

AOI221xp5_ASAP7_75t_SL g5703 ( 
.A1(n_5693),
.A2(n_1269),
.B1(n_1265),
.B2(n_1268),
.C(n_1270),
.Y(n_5703)
);

INVx3_ASAP7_75t_L g5704 ( 
.A(n_5657),
.Y(n_5704)
);

OR2x2_ASAP7_75t_L g5705 ( 
.A(n_5629),
.B(n_1271),
.Y(n_5705)
);

AOI21xp5_ASAP7_75t_L g5706 ( 
.A1(n_5636),
.A2(n_1272),
.B(n_1273),
.Y(n_5706)
);

HB1xp67_ASAP7_75t_L g5707 ( 
.A(n_5686),
.Y(n_5707)
);

OAI21xp5_ASAP7_75t_SL g5708 ( 
.A1(n_5623),
.A2(n_1274),
.B(n_1276),
.Y(n_5708)
);

OAI22xp5_ASAP7_75t_L g5709 ( 
.A1(n_5652),
.A2(n_5631),
.B1(n_5694),
.B2(n_5644),
.Y(n_5709)
);

AOI222xp33_ASAP7_75t_L g5710 ( 
.A1(n_5627),
.A2(n_1282),
.B1(n_1284),
.B2(n_1278),
.C1(n_1281),
.C2(n_1283),
.Y(n_5710)
);

OAI32xp33_ASAP7_75t_L g5711 ( 
.A1(n_5690),
.A2(n_1290),
.A3(n_1285),
.B1(n_1287),
.B2(n_1292),
.Y(n_5711)
);

OAI21xp5_ASAP7_75t_SL g5712 ( 
.A1(n_5647),
.A2(n_1292),
.B(n_1294),
.Y(n_5712)
);

NAND2xp5_ASAP7_75t_L g5713 ( 
.A(n_5698),
.B(n_1298),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5697),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_5625),
.B(n_1300),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_5634),
.Y(n_5716)
);

NAND2xp5_ASAP7_75t_L g5717 ( 
.A(n_5691),
.B(n_1300),
.Y(n_5717)
);

OAI21xp5_ASAP7_75t_SL g5718 ( 
.A1(n_5632),
.A2(n_1304),
.B(n_1305),
.Y(n_5718)
);

AOI22xp5_ASAP7_75t_L g5719 ( 
.A1(n_5651),
.A2(n_1308),
.B1(n_1306),
.B2(n_1307),
.Y(n_5719)
);

OAI22xp5_ASAP7_75t_L g5720 ( 
.A1(n_5680),
.A2(n_1310),
.B1(n_1308),
.B2(n_1309),
.Y(n_5720)
);

NOR2xp67_ASAP7_75t_SL g5721 ( 
.A(n_5643),
.B(n_1311),
.Y(n_5721)
);

NAND3xp33_ASAP7_75t_L g5722 ( 
.A(n_5689),
.B(n_1587),
.C(n_1586),
.Y(n_5722)
);

XOR2x2_ASAP7_75t_L g5723 ( 
.A(n_5637),
.B(n_1312),
.Y(n_5723)
);

AOI22xp33_ASAP7_75t_L g5724 ( 
.A1(n_5659),
.A2(n_1315),
.B1(n_1313),
.B2(n_1314),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5654),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5663),
.Y(n_5726)
);

AOI21xp5_ASAP7_75t_SL g5727 ( 
.A1(n_5635),
.A2(n_1314),
.B(n_1315),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5675),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5674),
.Y(n_5729)
);

AOI21xp5_ASAP7_75t_L g5730 ( 
.A1(n_5696),
.A2(n_1316),
.B(n_1317),
.Y(n_5730)
);

OAI221xp5_ASAP7_75t_SL g5731 ( 
.A1(n_5683),
.A2(n_1319),
.B1(n_1317),
.B2(n_1318),
.C(n_1320),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5649),
.Y(n_5732)
);

HB1xp67_ASAP7_75t_L g5733 ( 
.A(n_5679),
.Y(n_5733)
);

NAND2xp5_ASAP7_75t_L g5734 ( 
.A(n_5642),
.B(n_1322),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5669),
.Y(n_5735)
);

AOI211xp5_ASAP7_75t_L g5736 ( 
.A1(n_5628),
.A2(n_1328),
.B(n_1326),
.C(n_1327),
.Y(n_5736)
);

AND4x1_ASAP7_75t_L g5737 ( 
.A(n_5664),
.B(n_1331),
.C(n_1329),
.D(n_1330),
.Y(n_5737)
);

AND2x2_ASAP7_75t_L g5738 ( 
.A(n_5658),
.B(n_1332),
.Y(n_5738)
);

AOI222xp33_ASAP7_75t_L g5739 ( 
.A1(n_5633),
.A2(n_1337),
.B1(n_1340),
.B2(n_1335),
.C1(n_1336),
.C2(n_1338),
.Y(n_5739)
);

AOI21xp5_ASAP7_75t_L g5740 ( 
.A1(n_5638),
.A2(n_1340),
.B(n_1341),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5688),
.Y(n_5741)
);

AOI221xp5_ASAP7_75t_L g5742 ( 
.A1(n_5655),
.A2(n_1344),
.B1(n_1347),
.B2(n_1343),
.C(n_1346),
.Y(n_5742)
);

NAND2xp5_ASAP7_75t_L g5743 ( 
.A(n_5645),
.B(n_1342),
.Y(n_5743)
);

OAI21xp33_ASAP7_75t_L g5744 ( 
.A1(n_5684),
.A2(n_1348),
.B(n_1349),
.Y(n_5744)
);

BUFx2_ASAP7_75t_L g5745 ( 
.A(n_5704),
.Y(n_5745)
);

AOI322xp5_ASAP7_75t_L g5746 ( 
.A1(n_5733),
.A2(n_5640),
.A3(n_5668),
.B1(n_5682),
.B2(n_5678),
.C1(n_5665),
.C2(n_5646),
.Y(n_5746)
);

INVx2_ASAP7_75t_L g5747 ( 
.A(n_5704),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5707),
.Y(n_5748)
);

AOI21xp5_ASAP7_75t_L g5749 ( 
.A1(n_5727),
.A2(n_5670),
.B(n_5650),
.Y(n_5749)
);

AOI22xp33_ASAP7_75t_L g5750 ( 
.A1(n_5702),
.A2(n_5666),
.B1(n_5687),
.B2(n_5639),
.Y(n_5750)
);

OAI211xp5_ASAP7_75t_L g5751 ( 
.A1(n_5708),
.A2(n_5624),
.B(n_5677),
.C(n_5661),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5715),
.Y(n_5752)
);

AOI22xp5_ASAP7_75t_L g5753 ( 
.A1(n_5741),
.A2(n_5673),
.B1(n_5630),
.B2(n_5685),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5700),
.Y(n_5754)
);

CKINVDCx5p33_ASAP7_75t_R g5755 ( 
.A(n_5723),
.Y(n_5755)
);

AOI221xp5_ASAP7_75t_L g5756 ( 
.A1(n_5731),
.A2(n_5667),
.B1(n_5660),
.B2(n_5656),
.C(n_5648),
.Y(n_5756)
);

OR2x2_ASAP7_75t_L g5757 ( 
.A(n_5743),
.B(n_5692),
.Y(n_5757)
);

AOI22xp5_ASAP7_75t_L g5758 ( 
.A1(n_5709),
.A2(n_5662),
.B1(n_5641),
.B2(n_5676),
.Y(n_5758)
);

CKINVDCx6p67_ASAP7_75t_R g5759 ( 
.A(n_5738),
.Y(n_5759)
);

A2O1A1Ixp33_ASAP7_75t_L g5760 ( 
.A1(n_5722),
.A2(n_5671),
.B(n_5626),
.C(n_5681),
.Y(n_5760)
);

OAI211xp5_ASAP7_75t_SL g5761 ( 
.A1(n_5732),
.A2(n_5716),
.B(n_5735),
.C(n_5728),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5705),
.Y(n_5762)
);

NAND2xp5_ASAP7_75t_L g5763 ( 
.A(n_5721),
.B(n_1351),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5713),
.Y(n_5764)
);

INVxp67_ASAP7_75t_SL g5765 ( 
.A(n_5740),
.Y(n_5765)
);

AOI221xp5_ASAP7_75t_L g5766 ( 
.A1(n_5720),
.A2(n_1355),
.B1(n_1352),
.B2(n_1354),
.C(n_1356),
.Y(n_5766)
);

A2O1A1Ixp33_ASAP7_75t_SL g5767 ( 
.A1(n_5726),
.A2(n_1357),
.B(n_1355),
.C(n_1356),
.Y(n_5767)
);

OAI22xp33_ASAP7_75t_SL g5768 ( 
.A1(n_5729),
.A2(n_1360),
.B1(n_1358),
.B2(n_1359),
.Y(n_5768)
);

AOI22xp5_ASAP7_75t_L g5769 ( 
.A1(n_5699),
.A2(n_1363),
.B1(n_1361),
.B2(n_1362),
.Y(n_5769)
);

OAI21xp5_ASAP7_75t_L g5770 ( 
.A1(n_5706),
.A2(n_1365),
.B(n_1366),
.Y(n_5770)
);

OR2x2_ASAP7_75t_L g5771 ( 
.A(n_5734),
.B(n_1365),
.Y(n_5771)
);

OAI21xp5_ASAP7_75t_L g5772 ( 
.A1(n_5712),
.A2(n_1366),
.B(n_1367),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5717),
.Y(n_5773)
);

XOR2x2_ASAP7_75t_L g5774 ( 
.A(n_5737),
.B(n_5703),
.Y(n_5774)
);

AOI322xp5_ASAP7_75t_L g5775 ( 
.A1(n_5742),
.A2(n_1592),
.A3(n_1374),
.B1(n_1371),
.B2(n_1373),
.C1(n_1369),
.C2(n_1370),
.Y(n_5775)
);

OAI21xp5_ASAP7_75t_SL g5776 ( 
.A1(n_5718),
.A2(n_1372),
.B(n_1374),
.Y(n_5776)
);

NAND3xp33_ASAP7_75t_L g5777 ( 
.A(n_5745),
.B(n_5739),
.C(n_5736),
.Y(n_5777)
);

OAI21xp5_ASAP7_75t_L g5778 ( 
.A1(n_5749),
.A2(n_5701),
.B(n_5730),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5747),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_5748),
.Y(n_5780)
);

XNOR2x1_ASAP7_75t_L g5781 ( 
.A(n_5774),
.B(n_5755),
.Y(n_5781)
);

AOI22xp33_ASAP7_75t_L g5782 ( 
.A1(n_5759),
.A2(n_5725),
.B1(n_5714),
.B2(n_5710),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5765),
.Y(n_5783)
);

INVx2_ASAP7_75t_L g5784 ( 
.A(n_5771),
.Y(n_5784)
);

NAND2xp5_ASAP7_75t_SL g5785 ( 
.A(n_5768),
.B(n_5744),
.Y(n_5785)
);

OAI21xp5_ASAP7_75t_L g5786 ( 
.A1(n_5760),
.A2(n_5719),
.B(n_5724),
.Y(n_5786)
);

OAI211xp5_ASAP7_75t_L g5787 ( 
.A1(n_5758),
.A2(n_5711),
.B(n_1378),
.C(n_1376),
.Y(n_5787)
);

O2A1O1Ixp33_ASAP7_75t_L g5788 ( 
.A1(n_5767),
.A2(n_1379),
.B(n_1377),
.C(n_1378),
.Y(n_5788)
);

BUFx3_ASAP7_75t_L g5789 ( 
.A(n_5752),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5762),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_L g5791 ( 
.A(n_5750),
.B(n_1383),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_5757),
.Y(n_5792)
);

XNOR2xp5_ASAP7_75t_L g5793 ( 
.A(n_5753),
.B(n_1384),
.Y(n_5793)
);

INVx6_ASAP7_75t_L g5794 ( 
.A(n_5761),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5763),
.Y(n_5795)
);

NAND2xp5_ASAP7_75t_L g5796 ( 
.A(n_5775),
.B(n_1387),
.Y(n_5796)
);

AOI22xp5_ASAP7_75t_L g5797 ( 
.A1(n_5751),
.A2(n_1390),
.B1(n_1388),
.B2(n_1389),
.Y(n_5797)
);

OAI21xp33_ASAP7_75t_SL g5798 ( 
.A1(n_5746),
.A2(n_1393),
.B(n_1394),
.Y(n_5798)
);

OAI211xp5_ASAP7_75t_L g5799 ( 
.A1(n_5776),
.A2(n_1395),
.B(n_1393),
.C(n_1394),
.Y(n_5799)
);

AO22x2_ASAP7_75t_L g5800 ( 
.A1(n_5781),
.A2(n_5773),
.B1(n_5754),
.B2(n_5764),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_5793),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5789),
.Y(n_5802)
);

NOR2xp33_ASAP7_75t_L g5803 ( 
.A(n_5798),
.B(n_5799),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5791),
.Y(n_5804)
);

INVx2_ASAP7_75t_L g5805 ( 
.A(n_5794),
.Y(n_5805)
);

NOR2x1_ASAP7_75t_L g5806 ( 
.A(n_5783),
.B(n_5772),
.Y(n_5806)
);

NOR2x1_ASAP7_75t_L g5807 ( 
.A(n_5777),
.B(n_5770),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5780),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5797),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5792),
.Y(n_5810)
);

AOI22xp5_ASAP7_75t_L g5811 ( 
.A1(n_5790),
.A2(n_5756),
.B1(n_5766),
.B2(n_5769),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5779),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5796),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_5810),
.Y(n_5814)
);

XOR2xp5_ASAP7_75t_L g5815 ( 
.A(n_5811),
.B(n_5786),
.Y(n_5815)
);

OR2x2_ASAP7_75t_L g5816 ( 
.A(n_5802),
.B(n_5785),
.Y(n_5816)
);

XNOR2x1_ASAP7_75t_L g5817 ( 
.A(n_5807),
.B(n_5778),
.Y(n_5817)
);

INVx3_ASAP7_75t_L g5818 ( 
.A(n_5805),
.Y(n_5818)
);

XNOR2x1_ASAP7_75t_L g5819 ( 
.A(n_5800),
.B(n_5784),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_5803),
.B(n_5788),
.Y(n_5820)
);

OAI21xp5_ASAP7_75t_L g5821 ( 
.A1(n_5806),
.A2(n_5787),
.B(n_5782),
.Y(n_5821)
);

NOR2x1_ASAP7_75t_L g5822 ( 
.A(n_5808),
.B(n_5795),
.Y(n_5822)
);

AND4x1_ASAP7_75t_L g5823 ( 
.A(n_5821),
.B(n_5812),
.C(n_5813),
.D(n_5801),
.Y(n_5823)
);

AOI21xp33_ASAP7_75t_SL g5824 ( 
.A1(n_5819),
.A2(n_5809),
.B(n_5804),
.Y(n_5824)
);

OAI21xp33_ASAP7_75t_L g5825 ( 
.A1(n_5817),
.A2(n_1396),
.B(n_1397),
.Y(n_5825)
);

AOI21xp5_ASAP7_75t_L g5826 ( 
.A1(n_5820),
.A2(n_5815),
.B(n_5822),
.Y(n_5826)
);

OAI22xp33_ASAP7_75t_L g5827 ( 
.A1(n_5816),
.A2(n_1400),
.B1(n_1398),
.B2(n_1399),
.Y(n_5827)
);

HB1xp67_ASAP7_75t_L g5828 ( 
.A(n_5818),
.Y(n_5828)
);

NAND3xp33_ASAP7_75t_L g5829 ( 
.A(n_5814),
.B(n_1399),
.C(n_1400),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5828),
.Y(n_5830)
);

NOR3xp33_ASAP7_75t_L g5831 ( 
.A(n_5824),
.B(n_1402),
.C(n_1403),
.Y(n_5831)
);

XNOR2xp5_ASAP7_75t_L g5832 ( 
.A(n_5830),
.B(n_5823),
.Y(n_5832)
);

AND2x4_ASAP7_75t_SL g5833 ( 
.A(n_5831),
.B(n_5826),
.Y(n_5833)
);

OA21x2_ASAP7_75t_L g5834 ( 
.A1(n_5832),
.A2(n_5825),
.B(n_5829),
.Y(n_5834)
);

AND2x2_ASAP7_75t_SL g5835 ( 
.A(n_5834),
.B(n_5833),
.Y(n_5835)
);

INVx3_ASAP7_75t_L g5836 ( 
.A(n_5835),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5836),
.Y(n_5837)
);

XNOR2x1_ASAP7_75t_L g5838 ( 
.A(n_5837),
.B(n_5827),
.Y(n_5838)
);

AOI22xp33_ASAP7_75t_SL g5839 ( 
.A1(n_5838),
.A2(n_1407),
.B1(n_1404),
.B2(n_1406),
.Y(n_5839)
);

OAI221xp5_ASAP7_75t_R g5840 ( 
.A1(n_5839),
.A2(n_1410),
.B1(n_1408),
.B2(n_1409),
.C(n_1411),
.Y(n_5840)
);

AO21x2_ASAP7_75t_L g5841 ( 
.A1(n_5840),
.A2(n_1412),
.B(n_1413),
.Y(n_5841)
);

OAI22xp5_ASAP7_75t_L g5842 ( 
.A1(n_5841),
.A2(n_1417),
.B1(n_1414),
.B2(n_1416),
.Y(n_5842)
);

AOI211xp5_ASAP7_75t_L g5843 ( 
.A1(n_5842),
.A2(n_1589),
.B(n_1419),
.C(n_1418),
.Y(n_5843)
);


endmodule