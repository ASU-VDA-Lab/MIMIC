module fake_jpeg_327_n_58 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_17),
.B(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_18),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_23),
.Y(n_32)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_0),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_35),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_31),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.C(n_47),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_31),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_7),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI21x1_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_52),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_52),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_54),
.A3(n_50),
.B1(n_51),
.B2(n_5),
.C1(n_6),
.C2(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_6),
.Y(n_58)
);


endmodule