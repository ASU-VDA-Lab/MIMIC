module fake_netlist_5_530_n_1786 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1786);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1786;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_314;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_130),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_54),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_17),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_52),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_25),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_45),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_81),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_71),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_17),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_49),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_7),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_50),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_170),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_174),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_136),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_147),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_22),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_59),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_91),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_35),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_87),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_115),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_112),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_32),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_98),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_153),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_70),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_121),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_83),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_78),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_47),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_124),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_54),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_64),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_12),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_66),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_32),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_46),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_157),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_36),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_116),
.Y(n_265)
);

INVxp33_ASAP7_75t_R g266 ( 
.A(n_126),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_105),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_74),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_51),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_155),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_102),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_62),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_167),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_113),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_186),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_29),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_79),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_168),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_159),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_88),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_109),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_97),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_185),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_119),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_90),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_58),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_183),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_44),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_65),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_92),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_33),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_158),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_55),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_33),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_77),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_184),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_76),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_143),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_94),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_57),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_179),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_100),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_137),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_2),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_43),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_89),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_72),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_151),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_110),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_15),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_19),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_29),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_10),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_47),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_55),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_108),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_42),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_31),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_42),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_34),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_93),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_9),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_38),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_118),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_164),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_75),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_35),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_31),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_34),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_58),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_11),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_172),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_41),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_39),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_53),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_37),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_27),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_175),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_150),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_60),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_86),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_43),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_128),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_37),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_23),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_4),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_48),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_13),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_139),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_36),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_156),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_45),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_20),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_46),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_123),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_161),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_16),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_1),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_1),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_39),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_23),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_19),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_85),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_68),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_22),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_212),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_286),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_212),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_254),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_217),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_212),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_241),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_191),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_205),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_283),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_221),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_272),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_212),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_219),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_212),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_321),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_226),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_226),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_226),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_222),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_226),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_233),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_226),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_317),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_368),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_317),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_224),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_317),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_191),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_234),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_235),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_239),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_237),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_242),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_243),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_244),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_237),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_245),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_248),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_194),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_199),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_187),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_210),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_250),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_215),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_252),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_256),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_197),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_259),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_262),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_274),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_197),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_295),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_297),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_233),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_233),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_303),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_258),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_322),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_306),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_316),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_322),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_260),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_204),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_323),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_325),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_329),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_263),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_330),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_334),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_346),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_324),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_355),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_267),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_361),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_200),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_209),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_200),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_270),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_214),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_271),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_211),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_214),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_L g475 ( 
.A(n_382),
.B(n_357),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_384),
.B(n_192),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_390),
.B(n_459),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_192),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_381),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_398),
.B(n_198),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_198),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_428),
.B(n_350),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_386),
.B(n_357),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_450),
.B(n_350),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_409),
.B(n_315),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_408),
.B(n_315),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_396),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_390),
.B(n_459),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_218),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_391),
.Y(n_502)
);

CKINVDCx8_ASAP7_75t_R g503 ( 
.A(n_388),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_413),
.B(n_218),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_389),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_396),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_415),
.B(n_419),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_399),
.A2(n_265),
.B(n_255),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_473),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_389),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_389),
.B(n_205),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_420),
.B(n_255),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_422),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_406),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_265),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_454),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_465),
.B(n_281),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_392),
.A2(n_327),
.B1(n_261),
.B2(n_374),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_468),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_412),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_472),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_380),
.A2(n_378),
.B1(n_374),
.B2(n_373),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_473),
.B(n_370),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_393),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_471),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_432),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_432),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_387),
.B(n_281),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_414),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_397),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_463),
.B(n_338),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_407),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_463),
.B(n_338),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_470),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_388),
.A2(n_378),
.B1(n_373),
.B2(n_367),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_418),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_417),
.B(n_351),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_411),
.B(n_351),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_421),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_421),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_487),
.B(n_411),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_515),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_515),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_485),
.B(n_383),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_485),
.B(n_403),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_486),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_551),
.B(n_438),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_478),
.Y(n_563)
);

OAI21xp33_ASAP7_75t_SL g564 ( 
.A1(n_551),
.A2(n_370),
.B(n_424),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_482),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_511),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_485),
.B(n_403),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_498),
.B(n_441),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_478),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_551),
.Y(n_571)
);

AND3x2_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_445),
.C(n_404),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_507),
.A2(n_430),
.B1(n_444),
.B2(n_423),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_464),
.C(n_448),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_517),
.B(n_462),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_441),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_498),
.B(n_442),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_523),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_493),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_477),
.B(n_266),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_486),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_528),
.B(n_442),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_493),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_498),
.B(n_216),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_495),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_476),
.B(n_466),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_521),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_519),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_481),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_519),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_530),
.B(n_466),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_497),
.B(n_480),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_491),
.B(n_188),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_483),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_504),
.B(n_220),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_540),
.B(n_474),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_529),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_529),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_483),
.Y(n_607)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_492),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_SL g610 ( 
.A(n_547),
.B(n_358),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_512),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_489),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_489),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_537),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_490),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_490),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_516),
.B(n_236),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_496),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_496),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_506),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_522),
.B(n_296),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_513),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_495),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_531),
.A2(n_332),
.B1(n_294),
.B2(n_268),
.Y(n_627)
);

INVx6_ASAP7_75t_L g628 ( 
.A(n_479),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_533),
.Y(n_629)
);

AO21x2_ASAP7_75t_L g630 ( 
.A1(n_492),
.A2(n_231),
.B(n_225),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_494),
.B(n_531),
.C(n_533),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_479),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_538),
.B(n_313),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_506),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_541),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_508),
.Y(n_636)
);

NOR2x1p5_ASAP7_75t_L g637 ( 
.A(n_537),
.B(n_358),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_503),
.B(n_188),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_521),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_501),
.B(n_223),
.C(n_213),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_538),
.B(n_344),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_508),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_510),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_501),
.B(n_189),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_538),
.B(n_275),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_510),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

NOR2x1p5_ASAP7_75t_L g649 ( 
.A(n_501),
.B(n_359),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_514),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_518),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_518),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_543),
.A2(n_205),
.B1(n_208),
.B2(n_307),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_543),
.A2(n_205),
.B1(n_208),
.B2(n_307),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_512),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_538),
.B(n_277),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_520),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_532),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_501),
.B(n_426),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_525),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_535),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_547),
.A2(n_189),
.B1(n_190),
.B2(n_376),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_502),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g669 ( 
.A(n_526),
.B(n_359),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_525),
.B(n_190),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_525),
.B(n_278),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_512),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_521),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_521),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_524),
.Y(n_675)
);

BUFx6f_ASAP7_75t_SL g676 ( 
.A(n_525),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_549),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_512),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_486),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_526),
.A2(n_193),
.B1(n_207),
.B2(n_376),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_524),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_486),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_505),
.B(n_280),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_SL g684 ( 
.A(n_545),
.B(n_363),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_512),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_505),
.B(n_282),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_545),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_539),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_524),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_505),
.B(n_284),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_505),
.B(n_285),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_479),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_552),
.B(n_424),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_550),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_524),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_524),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_550),
.A2(n_276),
.B1(n_208),
.B2(n_229),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_524),
.Y(n_699)
);

INVxp67_ASAP7_75t_SL g700 ( 
.A(n_527),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_527),
.B(n_536),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_527),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_663),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_608),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_591),
.B(n_193),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_608),
.B(n_287),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_663),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_568),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_571),
.A2(n_292),
.B1(n_288),
.B2(n_289),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_571),
.A2(n_293),
.B1(n_291),
.B2(n_299),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_591),
.B(n_205),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_688),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_592),
.B(n_195),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_600),
.B(n_556),
.Y(n_714)
);

AO22x2_ASAP7_75t_L g715 ( 
.A1(n_631),
.A2(n_298),
.B1(n_251),
.B2(n_257),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_626),
.B(n_536),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_589),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_562),
.A2(n_302),
.B1(n_308),
.B2(n_309),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_667),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_668),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_565),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_668),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_626),
.B(n_536),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_629),
.B(n_527),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_629),
.A2(n_290),
.B1(n_333),
.B2(n_320),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_556),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_565),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_573),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_573),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_603),
.B(n_195),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_SL g731 ( 
.A1(n_669),
.A2(n_544),
.B1(n_542),
.B2(n_534),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_527),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_564),
.B(n_269),
.C(n_246),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_608),
.B(n_527),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_620),
.B(n_509),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_662),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_554),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_624),
.B(n_566),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_630),
.A2(n_509),
.B1(n_276),
.B2(n_229),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_578),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_604),
.B(n_471),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_578),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_637),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_635),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_558),
.B(n_509),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_559),
.B(n_196),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_662),
.B(n_426),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_579),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_574),
.B(n_539),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_581),
.B(n_196),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_560),
.B(n_201),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_555),
.B(n_546),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_555),
.B(n_546),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_630),
.A2(n_229),
.B1(n_208),
.B2(n_276),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_557),
.B(n_548),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_692),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_567),
.A2(n_328),
.B1(n_356),
.B2(n_354),
.Y(n_758)
);

O2A1O1Ixp5_ASAP7_75t_L g759 ( 
.A1(n_563),
.A2(n_377),
.B(n_369),
.C(n_273),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_569),
.B(n_201),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_557),
.B(n_687),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_687),
.B(n_548),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_583),
.B(n_474),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_694),
.B(n_336),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_616),
.B(n_324),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_649),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_694),
.B(n_353),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_579),
.Y(n_768)
);

AND2x2_ASAP7_75t_SL g769 ( 
.A(n_698),
.B(n_208),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_695),
.B(n_552),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_695),
.B(n_553),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_577),
.B(n_202),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_580),
.A2(n_314),
.B1(n_352),
.B2(n_348),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_635),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_617),
.B(n_202),
.Y(n_775)
);

OR2x6_ASAP7_75t_L g776 ( 
.A(n_583),
.B(n_427),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_662),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_644),
.B(n_203),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_633),
.B(n_553),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_630),
.A2(n_307),
.B1(n_276),
.B2(n_229),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_641),
.B(n_310),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_582),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_666),
.B(n_318),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_563),
.B(n_319),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_575),
.B(n_203),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_581),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_604),
.B(n_206),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_570),
.B(n_337),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_654),
.A2(n_229),
.B1(n_276),
.B2(n_307),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_601),
.B(n_206),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_570),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_588),
.B(n_513),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_596),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_596),
.A2(n_439),
.B(n_469),
.C(n_467),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_597),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_611),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_602),
.B(n_513),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_611),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_640),
.B(n_207),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_677),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_671),
.B(n_362),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_611),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_602),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_585),
.B(n_362),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_576),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_655),
.B(n_513),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_599),
.B(n_324),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_638),
.B(n_364),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_680),
.A2(n_365),
.B1(n_363),
.B2(n_367),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_676),
.A2(n_364),
.B1(n_307),
.B2(n_513),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_693),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_582),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_607),
.B(n_609),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_607),
.B(n_513),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_693),
.B(n_427),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_676),
.A2(n_341),
.B1(n_227),
.B2(n_228),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_676),
.A2(n_335),
.B1(n_230),
.B2(n_232),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_609),
.B(n_615),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_611),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_586),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_583),
.B(n_339),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_611),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_590),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_645),
.B(n_238),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_610),
.A2(n_365),
.B1(n_339),
.B2(n_467),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_590),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_615),
.B(n_513),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_618),
.B(n_429),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_593),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_618),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_619),
.B(n_429),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_619),
.B(n_431),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_622),
.B(n_431),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_622),
.B(n_433),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_627),
.B(n_240),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_583),
.B(n_339),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_247),
.C(n_249),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_643),
.B(n_647),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_643),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_647),
.B(n_433),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_665),
.B(n_253),
.Y(n_841)
);

AO221x1_ASAP7_75t_L g842 ( 
.A1(n_692),
.A2(n_469),
.B1(n_461),
.B2(n_460),
.C(n_458),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_684),
.B(n_264),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_595),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_648),
.B(n_279),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_648),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_653),
.B(n_435),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_653),
.B(n_435),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_661),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_661),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_595),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_598),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_612),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_670),
.B(n_436),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_572),
.B(n_300),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_683),
.B(n_436),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_625),
.B(n_301),
.Y(n_857)
);

AND2x6_ASAP7_75t_L g858 ( 
.A(n_681),
.B(n_437),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_692),
.B(n_437),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_646),
.B(n_304),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_708),
.B(n_625),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_757),
.B(n_657),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_719),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_757),
.B(n_612),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_614),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_811),
.B(n_614),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_726),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_769),
.A2(n_610),
.B1(n_669),
.B2(n_650),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_769),
.A2(n_642),
.B1(n_658),
.B2(n_659),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_739),
.B(n_621),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_748),
.B(n_623),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_733),
.B(n_686),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_713),
.B(n_690),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_800),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_713),
.B(n_691),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_726),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_730),
.B(n_634),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_SL g878 ( 
.A(n_809),
.B(n_841),
.C(n_837),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_714),
.B(n_634),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_733),
.B(n_636),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_714),
.B(n_636),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_720),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_745),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_860),
.A2(n_700),
.B1(n_664),
.B2(n_651),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_738),
.B(n_642),
.Y(n_885)
);

AND2x4_ASAP7_75t_SL g886 ( 
.A(n_708),
.B(n_650),
.Y(n_886)
);

OAI221xp5_ASAP7_75t_L g887 ( 
.A1(n_825),
.A2(n_326),
.B1(n_312),
.B2(n_331),
.C(n_342),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_846),
.B(n_651),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_730),
.B(n_658),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_SL g890 ( 
.A(n_809),
.B(n_305),
.C(n_345),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_747),
.B(n_860),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_708),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_708),
.B(n_625),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_722),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_786),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_737),
.B(n_625),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_737),
.B(n_625),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_774),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_737),
.B(n_659),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_747),
.B(n_791),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_777),
.B(n_660),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_793),
.B(n_660),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_755),
.A2(n_597),
.B1(n_632),
.B2(n_628),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_853),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_721),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_736),
.A2(n_701),
.B(n_664),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_776),
.B(n_439),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_742),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_803),
.B(n_673),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_830),
.B(n_673),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_750),
.A2(n_632),
.B1(n_628),
.B2(n_597),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_777),
.B(n_674),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_839),
.B(n_674),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_849),
.B(n_850),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_777),
.B(n_681),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_727),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_825),
.A2(n_347),
.B(n_455),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_712),
.B(n_597),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_795),
.B(n_689),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_703),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_766),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_728),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_707),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_R g924 ( 
.A(n_704),
.B(n_61),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_765),
.B(n_440),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_753),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_787),
.B(n_628),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_729),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_746),
.A2(n_702),
.B(n_699),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_741),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_856),
.A2(n_632),
.B1(n_628),
.B2(n_689),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_SL g932 ( 
.A(n_731),
.B(n_443),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_743),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_744),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_749),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_704),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_768),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_815),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_795),
.A2(n_594),
.B(n_613),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_752),
.B(n_685),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_754),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_815),
.B(n_443),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_813),
.B(n_696),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_752),
.B(n_685),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_854),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_796),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_756),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_796),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_835),
.B(n_632),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_858),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_807),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_782),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_762),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_854),
.Y(n_954)
);

NOR2x2_ASAP7_75t_L g955 ( 
.A(n_776),
.B(n_696),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_705),
.B(n_446),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_772),
.B(n_685),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_772),
.B(n_818),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_761),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_838),
.B(n_561),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_848),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_770),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_755),
.A2(n_697),
.B1(n_598),
.B2(n_605),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_771),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_751),
.B(n_594),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_812),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_781),
.B(n_697),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_715),
.A2(n_605),
.B1(n_606),
.B2(n_447),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_820),
.Y(n_969)
);

NAND2x1p5_ASAP7_75t_L g970 ( 
.A(n_796),
.B(n_594),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_796),
.Y(n_971)
);

BUFx8_ASAP7_75t_L g972 ( 
.A(n_821),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_715),
.A2(n_606),
.B1(n_446),
.B2(n_447),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_848),
.B(n_451),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_763),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_823),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_785),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_836),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_785),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_845),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_715),
.A2(n_780),
.B1(n_789),
.B2(n_842),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_826),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_780),
.A2(n_456),
.B1(n_451),
.B2(n_452),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_829),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_858),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_763),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_716),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_779),
.B(n_656),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_789),
.A2(n_456),
.B1(n_452),
.B2(n_453),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_856),
.B(n_453),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_858),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_723),
.B(n_682),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_798),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_844),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_851),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_858),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_859),
.B(n_682),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_763),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_740),
.B(n_682),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_SL g1000 ( 
.A(n_843),
.B(n_455),
.C(n_457),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_852),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_724),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_828),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_824),
.B(n_613),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_709),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_740),
.B(n_679),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_734),
.B1(n_824),
.B2(n_801),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_734),
.A2(n_767),
.B1(n_764),
.B2(n_788),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_855),
.B(n_457),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_855),
.B(n_613),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_798),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_831),
.Y(n_1012)
);

INVx8_ASAP7_75t_L g1013 ( 
.A(n_858),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_775),
.B(n_679),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_832),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_833),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_834),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_784),
.B(n_639),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_775),
.B(n_778),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_799),
.B(n_458),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_778),
.B(n_561),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_840),
.B(n_460),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_798),
.B(n_656),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_847),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_802),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_792),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_808),
.Y(n_1027)
);

AND2x6_ASAP7_75t_L g1028 ( 
.A(n_810),
.B(n_587),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_797),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_802),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_711),
.B(n_561),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_891),
.B(n_783),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_1005),
.A2(n_710),
.B1(n_817),
.B2(n_816),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1019),
.B(n_760),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_983),
.A2(n_711),
.B1(n_725),
.B2(n_790),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_958),
.B(n_718),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_971),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_936),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_873),
.A2(n_758),
.B(n_773),
.C(n_827),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_959),
.B(n_732),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_983),
.A2(n_814),
.B1(n_804),
.B2(n_735),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_977),
.B(n_802),
.Y(n_1043)
);

O2A1O1Ixp5_ASAP7_75t_SL g1044 ( 
.A1(n_967),
.A2(n_857),
.B(n_461),
.C(n_425),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_873),
.A2(n_857),
.B(n_759),
.C(n_639),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_979),
.B(n_706),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_903),
.A2(n_862),
.B(n_948),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_948),
.A2(n_1018),
.B(n_911),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_984),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_876),
.B(n_802),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_863),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_867),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_984),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_874),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_867),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_900),
.A2(n_794),
.B(n_759),
.C(n_806),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_925),
.B(n_794),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1007),
.A2(n_822),
.B1(n_819),
.B2(n_584),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_948),
.A2(n_822),
.B(n_819),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_948),
.A2(n_822),
.B(n_819),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_954),
.B(n_819),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_895),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1018),
.A2(n_639),
.B(n_675),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_962),
.B(n_652),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_964),
.B(n_652),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_938),
.B(n_678),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_961),
.B(n_425),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_879),
.B(n_587),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_864),
.A2(n_675),
.B(n_678),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_882),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_945),
.B(n_678),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_999),
.A2(n_675),
.B(n_678),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_905),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_SL g1074 ( 
.A(n_932),
.B(n_0),
.C(n_2),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_951),
.B(n_584),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_945),
.B(n_584),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1006),
.A2(n_939),
.B(n_1004),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_894),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_906),
.A2(n_678),
.B(n_672),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_SL g1080 ( 
.A(n_936),
.B(n_672),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1004),
.A2(n_672),
.B(n_656),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_880),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_883),
.Y(n_1083)
);

AO32x1_ASAP7_75t_L g1084 ( 
.A1(n_963),
.A2(n_0),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_936),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_883),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_908),
.B(n_672),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_888),
.B(n_166),
.Y(n_1088)
);

NAND2x1_ASAP7_75t_L g1089 ( 
.A(n_946),
.B(n_163),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_888),
.B(n_162),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_879),
.B(n_154),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_865),
.B(n_3),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_SL g1093 ( 
.A1(n_881),
.A2(n_5),
.B(n_7),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_898),
.B(n_138),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_881),
.B(n_131),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_SL g1096 ( 
.A1(n_875),
.A2(n_120),
.B(n_117),
.C(n_114),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_890),
.B(n_14),
.C(n_15),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_902),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1009),
.B(n_974),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1012),
.B(n_14),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_898),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_907),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_890),
.B(n_16),
.C(n_18),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1003),
.B(n_18),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_SL g1105 ( 
.A(n_924),
.B(n_20),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1012),
.B(n_21),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_981),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_875),
.A2(n_1010),
.B1(n_980),
.B2(n_927),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_916),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_889),
.A2(n_111),
.B(n_106),
.C(n_103),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_904),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1015),
.B(n_1016),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_SL g1113 ( 
.A(n_971),
.B(n_28),
.Y(n_1113)
);

O2A1O1Ixp5_ASAP7_75t_SL g1114 ( 
.A1(n_967),
.A2(n_28),
.B(n_30),
.C(n_38),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_1010),
.A2(n_101),
.B(n_96),
.C(n_95),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_998),
.B(n_84),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_914),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_922),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_871),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_981),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_921),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_953),
.B(n_69),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_993),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_907),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_909),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_910),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_949),
.A2(n_67),
.B(n_52),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_878),
.A2(n_51),
.B(n_53),
.C(n_56),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_942),
.B(n_57),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_949),
.A2(n_997),
.B(n_944),
.Y(n_1130)
);

OAI21xp33_ASAP7_75t_SL g1131 ( 
.A1(n_889),
.A2(n_1024),
.B(n_1017),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_926),
.B(n_941),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_907),
.B(n_975),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_868),
.A2(n_878),
.B1(n_869),
.B2(n_989),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_921),
.B(n_866),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_913),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_872),
.B(n_978),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_995),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_940),
.A2(n_957),
.B(n_960),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_868),
.A2(n_869),
.B1(n_989),
.B2(n_877),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_885),
.B(n_920),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_990),
.B(n_885),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_993),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_987),
.A2(n_947),
.B1(n_1022),
.B2(n_990),
.Y(n_1145)
);

CKINVDCx10_ASAP7_75t_R g1146 ( 
.A(n_972),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_870),
.B(n_1002),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1022),
.B(n_920),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_L g1149 ( 
.A1(n_988),
.A2(n_927),
.B(n_965),
.C(n_943),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_SL g1150 ( 
.A(n_965),
.B(n_946),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_928),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_968),
.A2(n_1008),
.B1(n_923),
.B2(n_973),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1001),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_887),
.A2(n_917),
.B1(n_1027),
.B2(n_986),
.C(n_973),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1020),
.B(n_956),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_943),
.A2(n_1000),
.B(n_901),
.C(n_899),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_930),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_919),
.A2(n_918),
.B(n_970),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_933),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1020),
.B(n_934),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_935),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_937),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_919),
.A2(n_918),
.B(n_970),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_952),
.Y(n_1164)
);

XOR2x2_ASAP7_75t_SL g1165 ( 
.A(n_972),
.B(n_1021),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_892),
.B(n_991),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_1026),
.A2(n_1029),
.B(n_899),
.C(n_901),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1117),
.B(n_982),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1077),
.A2(n_1014),
.B(n_988),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1128),
.A2(n_912),
.B(n_915),
.C(n_976),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1134),
.A2(n_931),
.B1(n_884),
.B2(n_886),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1051),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1131),
.A2(n_992),
.B(n_1031),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1112),
.B(n_994),
.Y(n_1174)
);

AOI211x1_ASAP7_75t_L g1175 ( 
.A1(n_1107),
.A2(n_1023),
.B(n_912),
.C(n_915),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1149),
.A2(n_1028),
.B(n_1023),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1137),
.B(n_924),
.Y(n_1177)
);

AOI221x1_ASAP7_75t_L g1178 ( 
.A1(n_1134),
.A2(n_1011),
.B1(n_969),
.B2(n_966),
.C(n_1028),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1132),
.B(n_1033),
.Y(n_1179)
);

BUFx4_ASAP7_75t_SL g1180 ( 
.A(n_1062),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1146),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1132),
.B(n_886),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1049),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_L g1184 ( 
.A(n_1083),
.B(n_896),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1140),
.A2(n_1011),
.B1(n_991),
.B2(n_985),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1143),
.B(n_985),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_1040),
.A2(n_896),
.B(n_897),
.C(n_861),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1130),
.A2(n_1028),
.A3(n_1013),
.B(n_950),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1147),
.B(n_1098),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1034),
.A2(n_950),
.B1(n_996),
.B2(n_1028),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1054),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1072),
.A2(n_893),
.B(n_897),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1139),
.A2(n_1028),
.B(n_996),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1032),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_1032),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1140),
.A2(n_1011),
.B1(n_1025),
.B2(n_1013),
.Y(n_1196)
);

AO21x2_ASAP7_75t_L g1197 ( 
.A1(n_1079),
.A2(n_1048),
.B(n_1047),
.Y(n_1197)
);

O2A1O1Ixp5_ASAP7_75t_L g1198 ( 
.A1(n_1091),
.A2(n_1095),
.B(n_1046),
.C(n_1036),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1158),
.A2(n_1163),
.B(n_1069),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1035),
.B(n_1057),
.Y(n_1200)
);

NOR2xp67_ASAP7_75t_SL g1201 ( 
.A(n_1032),
.B(n_1121),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1063),
.A2(n_1041),
.B(n_1081),
.Y(n_1202)
);

BUFx10_ASAP7_75t_L g1203 ( 
.A(n_1106),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1055),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1045),
.A2(n_1068),
.B(n_1091),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1145),
.B(n_1082),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1167),
.A2(n_1095),
.B(n_1150),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1150),
.A2(n_1068),
.B(n_1042),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1082),
.B(n_1125),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1115),
.A2(n_1058),
.B(n_1096),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1056),
.A2(n_1044),
.B(n_1042),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1059),
.A2(n_1060),
.B(n_1065),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1142),
.A2(n_1152),
.B(n_1122),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1152),
.A2(n_1122),
.B(n_1136),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_1036),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1135),
.B(n_1160),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1107),
.A2(n_1120),
.A3(n_1127),
.B(n_1064),
.Y(n_1217)
);

AOI221xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1120),
.A2(n_1093),
.B1(n_1104),
.B2(n_1154),
.C(n_1119),
.Y(n_1218)
);

CKINVDCx16_ASAP7_75t_R g1219 ( 
.A(n_1116),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1052),
.B(n_1155),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_SL g1221 ( 
.A(n_1129),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1105),
.B(n_1092),
.C(n_1148),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1126),
.B(n_1100),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1043),
.A2(n_1071),
.B(n_1061),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1053),
.A2(n_1075),
.B(n_1090),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_SL g1226 ( 
.A1(n_1066),
.A2(n_1088),
.B(n_1138),
.C(n_1153),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1111),
.A2(n_1161),
.B(n_1164),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1039),
.B(n_1085),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1162),
.A2(n_1073),
.B1(n_1159),
.B2(n_1118),
.C(n_1157),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_SL g1230 ( 
.A1(n_1109),
.A2(n_1151),
.B(n_1165),
.Y(n_1230)
);

O2A1O1Ixp5_ASAP7_75t_L g1231 ( 
.A1(n_1113),
.A2(n_1089),
.B(n_1080),
.C(n_1087),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1101),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1097),
.A2(n_1103),
.B(n_1129),
.C(n_1094),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1067),
.B(n_1076),
.Y(n_1234)
);

NOR3xp33_ASAP7_75t_L g1235 ( 
.A(n_1141),
.B(n_1124),
.C(n_1102),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1070),
.B(n_1078),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1050),
.B(n_1166),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1094),
.B(n_1038),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1123),
.A2(n_1144),
.B(n_1084),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1144),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1084),
.A2(n_891),
.B(n_1007),
.C(n_873),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1037),
.A2(n_891),
.B(n_1007),
.C(n_873),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1131),
.A2(n_891),
.B(n_1149),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1099),
.B(n_1143),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1099),
.B(n_1143),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1038),
.Y(n_1247)
);

AOI31xp67_ASAP7_75t_L g1248 ( 
.A1(n_1108),
.A2(n_1091),
.A3(n_1095),
.B(n_1008),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1134),
.A2(n_891),
.B1(n_983),
.B2(n_780),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1077),
.A2(n_1130),
.A3(n_1047),
.B(n_1139),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1133),
.B(n_1094),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1128),
.A2(n_891),
.B(n_713),
.C(n_1019),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1099),
.B(n_805),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1077),
.A2(n_1130),
.A3(n_1047),
.B(n_1139),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1134),
.A2(n_891),
.B1(n_983),
.B2(n_780),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1131),
.A2(n_891),
.B(n_1149),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1086),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1121),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1134),
.A2(n_903),
.B(n_795),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1112),
.B(n_391),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1039),
.Y(n_1267)
);

AOI31xp67_ASAP7_75t_L g1268 ( 
.A1(n_1108),
.A2(n_1091),
.A3(n_1095),
.B(n_1008),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1082),
.B(n_677),
.Y(n_1271)
);

CKINVDCx8_ASAP7_75t_R g1272 ( 
.A(n_1146),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1134),
.A2(n_891),
.B1(n_983),
.B2(n_780),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1121),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1277)
);

INVx3_ASAP7_75t_SL g1278 ( 
.A(n_1062),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1039),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1054),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1156),
.A2(n_1122),
.B(n_1128),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1108),
.B(n_891),
.C(n_713),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1062),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1072),
.A2(n_929),
.B(n_1077),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1131),
.A2(n_891),
.B(n_1149),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1082),
.B(n_677),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1083),
.B(n_895),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_L g1290 ( 
.A(n_1112),
.B(n_891),
.Y(n_1290)
);

AND3x4_ASAP7_75t_L g1291 ( 
.A(n_1121),
.B(n_722),
.C(n_720),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1131),
.A2(n_891),
.B(n_1149),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1077),
.A2(n_795),
.B(n_903),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1131),
.A2(n_891),
.B(n_1149),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1107),
.A2(n_1120),
.B1(n_1134),
.B2(n_1128),
.C(n_1140),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1099),
.B(n_805),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1099),
.B(n_805),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1037),
.A2(n_891),
.B(n_1007),
.C(n_873),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1198),
.A2(n_1298),
.B(n_1243),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1179),
.A2(n_1275),
.B1(n_1258),
.B2(n_1250),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1282),
.A2(n_1241),
.B(n_1254),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1250),
.A2(n_1275),
.B1(n_1258),
.B2(n_1282),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1199),
.A2(n_1212),
.B(n_1192),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1293),
.A2(n_1249),
.B(n_1242),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_SL g1307 ( 
.A(n_1253),
.B(n_1222),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1283),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1189),
.A2(n_1200),
.B1(n_1253),
.B2(n_1223),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1180),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1247),
.B(n_1201),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1207),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1195),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1202),
.A2(n_1264),
.B(n_1290),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1244),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1208),
.A2(n_1213),
.B(n_1214),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1233),
.A2(n_1218),
.B(n_1222),
.C(n_1295),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1218),
.A2(n_1295),
.B(n_1286),
.C(n_1292),
.Y(n_1319)
);

INVx5_ASAP7_75t_L g1320 ( 
.A(n_1247),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1251),
.A2(n_1259),
.B(n_1256),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1215),
.A2(n_1244),
.B(n_1294),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1172),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1247),
.B(n_1267),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1220),
.B(n_1209),
.Y(n_1325)
);

NAND2x1_ASAP7_75t_L g1326 ( 
.A(n_1267),
.B(n_1279),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1169),
.A2(n_1193),
.B(n_1260),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1263),
.A2(n_1270),
.B(n_1266),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1216),
.B(n_1186),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1260),
.A2(n_1286),
.B(n_1292),
.C(n_1294),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1273),
.A2(n_1284),
.B(n_1285),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1173),
.B(n_1205),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1265),
.A2(n_1177),
.B1(n_1255),
.B2(n_1296),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1191),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1194),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1281),
.A2(n_1206),
.B1(n_1203),
.B2(n_1171),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1272),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1269),
.A2(n_1300),
.B1(n_1299),
.B2(n_1289),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1181),
.B(n_1219),
.Y(n_1339)
);

INVx8_ASAP7_75t_L g1340 ( 
.A(n_1247),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1176),
.A2(n_1239),
.B(n_1196),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1274),
.A2(n_1277),
.B1(n_1190),
.B2(n_1182),
.Y(n_1342)
);

AO32x2_ASAP7_75t_L g1343 ( 
.A1(n_1171),
.A2(n_1185),
.A3(n_1196),
.B1(n_1248),
.B2(n_1268),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1176),
.A2(n_1226),
.B(n_1185),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1210),
.A2(n_1197),
.A3(n_1205),
.B(n_1257),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1170),
.A2(n_1187),
.B(n_1231),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1280),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1229),
.A2(n_1225),
.B(n_1224),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1204),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1174),
.A2(n_1237),
.B(n_1168),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1228),
.A2(n_1230),
.B(n_1238),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1236),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1252),
.A2(n_1257),
.A3(n_1188),
.B(n_1175),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1184),
.A2(n_1252),
.B(n_1257),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1195),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1229),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1271),
.B(n_1287),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1234),
.A2(n_1297),
.B(n_1188),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1288),
.B(n_1232),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1188),
.A2(n_1235),
.B(n_1217),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1261),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1278),
.B(n_1262),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1221),
.A2(n_1291),
.B1(n_1276),
.B2(n_1240),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1200),
.B(n_1179),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_L g1365 ( 
.A(n_1179),
.B(n_1291),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1282),
.A2(n_1074),
.B1(n_891),
.B2(n_1134),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1191),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1194),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1282),
.A2(n_1074),
.B1(n_891),
.B2(n_1134),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1244),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1178),
.A2(n_1241),
.A3(n_1207),
.B(n_1208),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1265),
.A2(n_549),
.B1(n_391),
.B2(n_393),
.Y(n_1372)
);

AO32x2_ASAP7_75t_L g1373 ( 
.A1(n_1250),
.A2(n_1120),
.A3(n_1107),
.B1(n_1275),
.B2(n_1258),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1227),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_SL g1375 ( 
.A(n_1253),
.B(n_936),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1282),
.A2(n_1074),
.B1(n_891),
.B2(n_1134),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1180),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1244),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1200),
.B(n_891),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1198),
.A2(n_1298),
.B(n_1243),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1282),
.A2(n_1074),
.B1(n_891),
.B2(n_1134),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1227),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1200),
.B(n_891),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1244),
.Y(n_1384)
);

AOI21xp33_ASAP7_75t_L g1385 ( 
.A1(n_1254),
.A2(n_891),
.B(n_1282),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1200),
.B(n_891),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1267),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1254),
.A2(n_891),
.B(n_1298),
.C(n_1243),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1247),
.B(n_1080),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1200),
.B(n_891),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1244),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1195),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1180),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1207),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1244),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1396)
);

NOR2x1_ASAP7_75t_L g1397 ( 
.A(n_1179),
.B(n_1291),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1199),
.A2(n_1212),
.B(n_1192),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1191),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1183),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1178),
.A2(n_1241),
.A3(n_1207),
.B(n_1208),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1282),
.A2(n_1074),
.B1(n_891),
.B2(n_1134),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1194),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1179),
.A2(n_1134),
.B1(n_983),
.B2(n_1250),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1243),
.A2(n_1298),
.B(n_891),
.C(n_1254),
.Y(n_1405)
);

AO32x2_ASAP7_75t_L g1406 ( 
.A1(n_1250),
.A2(n_1120),
.A3(n_1107),
.B1(n_1275),
.B2(n_1258),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1254),
.A2(n_713),
.B1(n_1295),
.B2(n_1134),
.C(n_1282),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1325),
.B(n_1352),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1349),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1366),
.A2(n_1376),
.B1(n_1381),
.B2(n_1369),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1349),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1314),
.A2(n_1327),
.B(n_1388),
.Y(n_1414)
);

O2A1O1Ixp5_ASAP7_75t_L g1415 ( 
.A1(n_1303),
.A2(n_1301),
.B(n_1380),
.C(n_1385),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1361),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1369),
.A2(n_1402),
.B1(n_1376),
.B2(n_1381),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1392),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1304),
.A2(n_1364),
.B1(n_1386),
.B2(n_1390),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1303),
.A2(n_1301),
.B(n_1380),
.C(n_1302),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1386),
.B(n_1390),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1357),
.B(n_1309),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1405),
.A2(n_1311),
.B(n_1375),
.Y(n_1423)
);

AOI211xp5_ASAP7_75t_L g1424 ( 
.A1(n_1407),
.A2(n_1317),
.B(n_1338),
.C(n_1309),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1327),
.A2(n_1316),
.B(n_1330),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1332),
.A2(n_1404),
.B(n_1319),
.Y(n_1426)
);

AND2x4_ASAP7_75t_SL g1427 ( 
.A(n_1308),
.B(n_1359),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1304),
.A2(n_1365),
.B1(n_1397),
.B2(n_1336),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1329),
.B(n_1357),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1311),
.A2(n_1389),
.B(n_1338),
.Y(n_1430)
);

INVx3_ASAP7_75t_SL g1431 ( 
.A(n_1310),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1350),
.A2(n_1332),
.B(n_1344),
.C(n_1358),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1372),
.B(n_1334),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1389),
.A2(n_1359),
.B(n_1307),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1342),
.A2(n_1341),
.B(n_1351),
.C(n_1356),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1342),
.A2(n_1363),
.B1(n_1320),
.B2(n_1395),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1374),
.A2(n_1382),
.B(n_1322),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1320),
.A2(n_1395),
.B1(n_1370),
.B2(n_1378),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1347),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1320),
.A2(n_1391),
.B1(n_1384),
.B2(n_1370),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1337),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1367),
.A2(n_1399),
.B(n_1322),
.C(n_1394),
.Y(n_1442)
);

OR2x2_ASAP7_75t_SL g1443 ( 
.A(n_1400),
.B(n_1368),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1360),
.B(n_1353),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1312),
.A2(n_1355),
.B(n_1313),
.C(n_1362),
.Y(n_1445)
);

O2A1O1Ixp5_ASAP7_75t_L g1446 ( 
.A1(n_1374),
.A2(n_1382),
.B(n_1326),
.C(n_1387),
.Y(n_1446)
);

NOR2xp67_ASAP7_75t_L g1447 ( 
.A(n_1377),
.B(n_1393),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1339),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_L g1449 ( 
.A(n_1335),
.B(n_1403),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1315),
.A2(n_1391),
.B1(n_1384),
.B2(n_1378),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1354),
.A2(n_1324),
.B(n_1348),
.C(n_1373),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1306),
.A2(n_1331),
.B(n_1321),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1373),
.A2(n_1406),
.B1(n_1368),
.B2(n_1348),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1373),
.A2(n_1406),
.B(n_1343),
.C(n_1371),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1406),
.B(n_1401),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1371),
.B(n_1401),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1343),
.A2(n_1345),
.B1(n_1328),
.B2(n_1305),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1343),
.B(n_1345),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1398),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1346),
.A2(n_1303),
.B(n_1301),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1314),
.A2(n_891),
.B(n_1243),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_SL g1464 ( 
.A1(n_1303),
.A2(n_713),
.B(n_1046),
.C(n_1113),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1388),
.A2(n_1298),
.B(n_1243),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1314),
.A2(n_891),
.B(n_1243),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1365),
.A2(n_1397),
.B1(n_1333),
.B2(n_1369),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1323),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1325),
.B(n_1352),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1318),
.B(n_1396),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1325),
.B(n_1352),
.Y(n_1477)
);

NOR2xp67_ASAP7_75t_L g1478 ( 
.A(n_1333),
.B(n_1271),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1388),
.A2(n_1298),
.B(n_1243),
.Y(n_1479)
);

BUFx2_ASAP7_75t_SL g1480 ( 
.A(n_1308),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1346),
.A2(n_1303),
.B(n_1301),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1314),
.A2(n_891),
.B(n_1243),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1340),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_1120),
.B2(n_1134),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1414),
.A2(n_1432),
.B(n_1437),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_SL g1488 ( 
.A(n_1412),
.B(n_1417),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1426),
.A2(n_1425),
.B(n_1438),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1471),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1452),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1438),
.A2(n_1440),
.B(n_1457),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1453),
.Y(n_1493)
);

BUFx4f_ASAP7_75t_L g1494 ( 
.A(n_1462),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1465),
.B(n_1479),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1469),
.A2(n_1428),
.B1(n_1419),
.B2(n_1410),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1435),
.A2(n_1415),
.B(n_1420),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1452),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1441),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1482),
.B(n_1458),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1444),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1459),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1440),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1450),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1446),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1480),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1463),
.A2(n_1483),
.B(n_1468),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1451),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1454),
.B(n_1422),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1419),
.B(n_1409),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1423),
.B(n_1430),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1436),
.A2(n_1417),
.B(n_1412),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1421),
.B(n_1470),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1445),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1442),
.Y(n_1515)
);

INVxp67_ASAP7_75t_R g1516 ( 
.A(n_1428),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1424),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1443),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1411),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1413),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1408),
.B(n_1474),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1477),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1481),
.Y(n_1523)
);

OR2x6_ASAP7_75t_L g1524 ( 
.A(n_1434),
.B(n_1485),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1460),
.A2(n_1485),
.B(n_1461),
.Y(n_1525)
);

OR2x6_ASAP7_75t_SL g1526 ( 
.A(n_1515),
.B(n_1473),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1492),
.A2(n_1464),
.B(n_1460),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1504),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1491),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1500),
.B(n_1475),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1500),
.B(n_1429),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1493),
.B(n_1439),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1494),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1494),
.B(n_1472),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1489),
.B(n_1472),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1501),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1490),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1489),
.B(n_1467),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1489),
.B(n_1467),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1476),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1487),
.B(n_1492),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1511),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1492),
.B(n_1493),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1492),
.B(n_1466),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1502),
.B(n_1484),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1535),
.A2(n_1495),
.B1(n_1525),
.B2(n_1488),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1546),
.A2(n_1517),
.B1(n_1488),
.B2(n_1496),
.C(n_1510),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1546),
.A2(n_1517),
.B1(n_1496),
.B2(n_1510),
.C(n_1461),
.Y(n_1552)
);

INVx3_ASAP7_75t_SL g1553 ( 
.A(n_1547),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1529),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1543),
.B(n_1503),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1547),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1535),
.A2(n_1495),
.B1(n_1525),
.B2(n_1524),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1537),
.B(n_1508),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1547),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1538),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1535),
.A2(n_1495),
.B1(n_1525),
.B2(n_1524),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1535),
.A2(n_1495),
.B1(n_1525),
.B2(n_1524),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1539),
.B(n_1515),
.Y(n_1564)
);

OAI211xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1533),
.A2(n_1433),
.B(n_1523),
.C(n_1448),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1543),
.B(n_1503),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1543),
.B(n_1530),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1527),
.A2(n_1486),
.B(n_1505),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1508),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

AOI211xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1546),
.A2(n_1516),
.B(n_1478),
.C(n_1495),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1531),
.B(n_1486),
.Y(n_1572)
);

AOI33xp33_ASAP7_75t_L g1573 ( 
.A1(n_1546),
.A2(n_1523),
.A3(n_1519),
.B1(n_1520),
.B2(n_1509),
.B3(n_1522),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1526),
.A2(n_1516),
.B1(n_1495),
.B2(n_1524),
.Y(n_1574)
);

OAI211xp5_ASAP7_75t_L g1575 ( 
.A1(n_1546),
.A2(n_1512),
.B(n_1497),
.C(n_1507),
.Y(n_1575)
);

OAI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1536),
.A2(n_1513),
.B(n_1509),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1536),
.A2(n_1512),
.B1(n_1507),
.B2(n_1511),
.C(n_1497),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1528),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1544),
.Y(n_1579)
);

OAI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1536),
.A2(n_1512),
.B1(n_1507),
.B2(n_1511),
.C(n_1497),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1550),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1579),
.B(n_1511),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1576),
.B(n_1531),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1558),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1558),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1549),
.B(n_1552),
.C(n_1571),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1575),
.A2(n_1545),
.B(n_1532),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_SL g1588 ( 
.A(n_1549),
.B(n_1536),
.C(n_1540),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1556),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1560),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1550),
.B(n_1545),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1575),
.A2(n_1545),
.B(n_1532),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1560),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1553),
.B(n_1531),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_SL g1595 ( 
.A(n_1571),
.B(n_1540),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1553),
.B(n_1534),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1579),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_R g1600 ( 
.A(n_1559),
.B(n_1506),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1556),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1553),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1564),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1570),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1534),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1568),
.A2(n_1527),
.B(n_1540),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1554),
.Y(n_1608)
);

NAND4xp25_ASAP7_75t_SL g1609 ( 
.A(n_1586),
.B(n_1552),
.C(n_1573),
.D(n_1548),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1599),
.B(n_1511),
.Y(n_1610)
);

NOR2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1586),
.B(n_1579),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1605),
.B(n_1567),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

AND2x4_ASAP7_75t_SL g1614 ( 
.A(n_1599),
.B(n_1511),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1602),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1584),
.B(n_1569),
.Y(n_1617)
);

CKINVDCx16_ASAP7_75t_R g1618 ( 
.A(n_1600),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1608),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1567),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1581),
.B(n_1572),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1555),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1593),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1593),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1585),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1594),
.B(n_1555),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1598),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1596),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1596),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1555),
.Y(n_1631)
);

AOI211x1_ASAP7_75t_L g1632 ( 
.A1(n_1588),
.A2(n_1566),
.B(n_1574),
.C(n_1577),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1599),
.B(n_1541),
.C(n_1540),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_1541),
.C(n_1540),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1584),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1608),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1602),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1603),
.B(n_1572),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1583),
.B(n_1499),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1595),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1587),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1591),
.A2(n_1580),
.B(n_1577),
.C(n_1563),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1604),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1582),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1582),
.B(n_1541),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.B(n_1566),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1587),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1602),
.B(n_1566),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1642),
.B(n_1595),
.Y(n_1651)
);

OAI31xp67_ASAP7_75t_L g1652 ( 
.A1(n_1609),
.A2(n_1595),
.A3(n_1607),
.B(n_1518),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1648),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1642),
.A2(n_1580),
.B1(n_1541),
.B2(n_1542),
.C(n_1607),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1636),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1625),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1613),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1613),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1611),
.B(n_1606),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1616),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1647),
.B(n_1589),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1617),
.B(n_1569),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1618),
.B(n_1431),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1627),
.Y(n_1665)
);

AND2x4_ASAP7_75t_SL g1666 ( 
.A(n_1646),
.B(n_1582),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1618),
.A2(n_1644),
.B(n_1635),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1633),
.A2(n_1607),
.B(n_1574),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1641),
.Y(n_1669)
);

NOR2xp67_ASAP7_75t_SL g1670 ( 
.A(n_1646),
.B(n_1418),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1632),
.A2(n_1526),
.B1(n_1562),
.B2(n_1557),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1639),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1631),
.B(n_1551),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1650),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1647),
.B(n_1589),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1616),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1650),
.B(n_1648),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1601),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1647),
.B(n_1646),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1647),
.B(n_1601),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1615),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1617),
.B(n_1606),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1615),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1612),
.B(n_1620),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1623),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1623),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1655),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1659),
.B(n_1612),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1657),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1656),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1672),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1684),
.B(n_1620),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1661),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1651),
.B(n_1682),
.Y(n_1695)
);

AOI222xp33_ASAP7_75t_L g1696 ( 
.A1(n_1654),
.A2(n_1541),
.B1(n_1542),
.B2(n_1649),
.C1(n_1643),
.C2(n_1565),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1667),
.A2(n_1542),
.B1(n_1527),
.B2(n_1610),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1684),
.B(n_1639),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1658),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1679),
.B(n_1616),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1681),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1683),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1664),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1679),
.B(n_1622),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1669),
.B(n_1665),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1653),
.B(n_1677),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1653),
.B(n_1622),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1664),
.B(n_1521),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1686),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1660),
.B(n_1626),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1671),
.A2(n_1542),
.B1(n_1527),
.B2(n_1610),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1687),
.B(n_1674),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1692),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1687),
.B(n_1682),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1697),
.A2(n_1668),
.B(n_1660),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1695),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1703),
.B(n_1670),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1712),
.A2(n_1652),
.B(n_1661),
.Y(n_1719)
);

AO22x1_ASAP7_75t_L g1720 ( 
.A1(n_1688),
.A2(n_1676),
.B1(n_1662),
.B2(n_1680),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1690),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1690),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1705),
.B(n_1666),
.Y(n_1723)
);

OAI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1696),
.A2(n_1707),
.B(n_1711),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1688),
.A2(n_1676),
.B(n_1675),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1691),
.A2(n_1649),
.B(n_1643),
.C(n_1607),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1691),
.A2(n_1542),
.B1(n_1666),
.B2(n_1587),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1695),
.A2(n_1675),
.B(n_1662),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1689),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1700),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1709),
.B(n_1698),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1711),
.A2(n_1610),
.B1(n_1680),
.B2(n_1678),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1722),
.Y(n_1733)
);

NAND2xp33_ASAP7_75t_L g1734 ( 
.A(n_1721),
.B(n_1700),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1722),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_L g1736 ( 
.A(n_1718),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1717),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1714),
.B(n_1693),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1723),
.B(n_1693),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1730),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1715),
.Y(n_1741)
);

INVx6_ASAP7_75t_L g1742 ( 
.A(n_1720),
.Y(n_1742)
);

NAND2x1_ASAP7_75t_L g1743 ( 
.A(n_1732),
.B(n_1693),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1729),
.Y(n_1744)
);

NAND2x1_ASAP7_75t_L g1745 ( 
.A(n_1742),
.B(n_1693),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1734),
.B(n_1719),
.C(n_1725),
.Y(n_1746)
);

OAI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1743),
.A2(n_1716),
.B(n_1727),
.C(n_1724),
.Y(n_1747)
);

AOI322xp5_ASAP7_75t_L g1748 ( 
.A1(n_1733),
.A2(n_1727),
.A3(n_1713),
.B1(n_1731),
.B2(n_1708),
.C1(n_1704),
.C2(n_1692),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1735),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1740),
.A2(n_1726),
.B(n_1728),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1740),
.B(n_1694),
.C(n_1689),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_SL g1752 ( 
.A(n_1741),
.B(n_1694),
.C(n_1698),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1739),
.A2(n_1710),
.B(n_1702),
.C(n_1701),
.Y(n_1753)
);

OAI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1742),
.A2(n_1610),
.B1(n_1694),
.B2(n_1592),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1746),
.A2(n_1737),
.B1(n_1610),
.B2(n_1744),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_SL g1756 ( 
.A1(n_1745),
.A2(n_1699),
.B(n_1701),
.C(n_1710),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1750),
.A2(n_1738),
.B(n_1702),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1751),
.Y(n_1758)
);

OAI31xp33_ASAP7_75t_L g1759 ( 
.A1(n_1747),
.A2(n_1736),
.A3(n_1699),
.B(n_1706),
.Y(n_1759)
);

NAND2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1758),
.B(n_1447),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_L g1761 ( 
.A(n_1757),
.B(n_1752),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1759),
.B(n_1749),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1756),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1755),
.B(n_1748),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1758),
.B(n_1753),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1754),
.B1(n_1704),
.B2(n_1706),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_L g1767 ( 
.A1(n_1761),
.A2(n_1708),
.B(n_1678),
.C(n_1592),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1762),
.B(n_1427),
.Y(n_1768)
);

AOI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1764),
.A2(n_1663),
.B(n_1634),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1763),
.A2(n_1527),
.B1(n_1582),
.B2(n_1614),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1767),
.B(n_1763),
.Y(n_1771)
);

NOR2x1p5_ASAP7_75t_L g1772 ( 
.A(n_1768),
.B(n_1760),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1769),
.A2(n_1614),
.B1(n_1527),
.B2(n_1663),
.Y(n_1773)
);

INVx4_ASAP7_75t_L g1774 ( 
.A(n_1772),
.Y(n_1774)
);

OAI22xp33_ASAP7_75t_R g1775 ( 
.A1(n_1774),
.A2(n_1771),
.B1(n_1766),
.B2(n_1770),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1775),
.Y(n_1776)
);

OR3x1_ASAP7_75t_L g1777 ( 
.A(n_1775),
.B(n_1773),
.C(n_1565),
.Y(n_1777)
);

OAI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1776),
.A2(n_1637),
.B1(n_1619),
.B2(n_1634),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1777),
.A2(n_1673),
.B(n_1416),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1779),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1780),
.B(n_1778),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1637),
.B1(n_1619),
.B2(n_1630),
.C(n_1645),
.Y(n_1782)
);

OAI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_1621),
.B(n_1640),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1629),
.B1(n_1645),
.B2(n_1630),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1624),
.B1(n_1628),
.B2(n_1638),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1449),
.B(n_1624),
.C(n_1628),
.Y(n_1786)
);


endmodule