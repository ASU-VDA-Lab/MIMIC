module fake_jpeg_15734_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_2),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_4),
.B1(n_7),
.B2(n_16),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_16),
.B1(n_14),
.B2(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_38),
.B1(n_27),
.B2(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_15),
.B1(n_38),
.B2(n_41),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_9),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_33),
.C(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_7),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx12f_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_48),
.C(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_49),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_43),
.C(n_39),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_45),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.C(n_44),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_53),
.B(n_35),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_36),
.B(n_37),
.Y(n_57)
);


endmodule