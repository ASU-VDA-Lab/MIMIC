module fake_jpeg_9707_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_26),
.Y(n_58)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_30),
.B1(n_31),
.B2(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_18),
.B1(n_26),
.B2(n_15),
.Y(n_66)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_25),
.B(n_16),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_51),
.B(n_15),
.C(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_19),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_28),
.B(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_64),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_68),
.B(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_47),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_14),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_53),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_16),
.B(n_25),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_25),
.B(n_27),
.C(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_67),
.B1(n_70),
.B2(n_45),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_86),
.B1(n_91),
.B2(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_45),
.B1(n_53),
.B2(n_43),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_69),
.C(n_56),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_57),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_47),
.B1(n_52),
.B2(n_49),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_22),
.B(n_61),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_42),
.C(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_100),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_107),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_27),
.B(n_17),
.C(n_22),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_92),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_102),
.Y(n_136)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_94),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_28),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_62),
.B1(n_23),
.B2(n_20),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_129),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_88),
.B1(n_77),
.B2(n_85),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_128),
.B(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_94),
.B1(n_95),
.B2(n_86),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_79),
.B1(n_64),
.B2(n_81),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_90),
.B(n_28),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_62),
.B1(n_54),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_109),
.B1(n_100),
.B2(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_28),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_134),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_116),
.B1(n_108),
.B2(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_150),
.B1(n_23),
.B2(n_20),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_97),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_120),
.B1(n_119),
.B2(n_132),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_104),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_109),
.C(n_98),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_101),
.B1(n_106),
.B2(n_113),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_122),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_28),
.B(n_1),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_0),
.B(n_1),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_128),
.C(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_167),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_136),
.B(n_124),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_165),
.B(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_23),
.B1(n_20),
.B2(n_2),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_23),
.B1(n_20),
.B2(n_12),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_12),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_171),
.A2(n_158),
.B(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_28),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_147),
.CI(n_140),
.CON(n_177),
.SN(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_0),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_151),
.C(n_144),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_182),
.C(n_184),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_138),
.C(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_149),
.C(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_192),
.C(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_159),
.C(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_3),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_198),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_3),
.B(n_4),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_181),
.B1(n_175),
.B2(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_182),
.C(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_207),
.C(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_179),
.C(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_212),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_177),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_204),
.C(n_205),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_8),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_9),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_223),
.A2(n_224),
.B(n_9),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_224),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_227),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_220),
.B(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_10),
.Y(n_230)
);


endmodule