module fake_jpeg_20054_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_37),
.B1(n_18),
.B2(n_32),
.Y(n_54)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_28),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_33),
.B1(n_29),
.B2(n_15),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_42),
.B1(n_40),
.B2(n_22),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_43),
.B1(n_46),
.B2(n_44),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_46),
.B1(n_44),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_40),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_41),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_79),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_32),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_16),
.B1(n_30),
.B2(n_24),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

AO21x1_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_101),
.B(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_46),
.B1(n_44),
.B2(n_40),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_42),
.B1(n_20),
.B2(n_15),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_20),
.B1(n_29),
.B2(n_31),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_16),
.B(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_31),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_38),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_41),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_110),
.A2(n_76),
.B1(n_81),
.B2(n_78),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_41),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_108),
.B1(n_104),
.B2(n_89),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_90),
.C(n_82),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_19),
.C(n_69),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_1),
.B(n_3),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_136),
.Y(n_143)
);

OAI22x1_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_80),
.B1(n_83),
.B2(n_107),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_38),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_147),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_150),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_135),
.B1(n_83),
.B2(n_36),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_102),
.C(n_99),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_167),
.C(n_170),
.Y(n_172)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_155),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_105),
.B1(n_81),
.B2(n_99),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_127),
.B1(n_135),
.B2(n_35),
.Y(n_194)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_136),
.B1(n_131),
.B2(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_159),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_112),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_35),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_127),
.B1(n_125),
.B2(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_95),
.B1(n_87),
.B2(n_36),
.Y(n_197)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_19),
.Y(n_203)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_76),
.C(n_74),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_75),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_113),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_87),
.C(n_41),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_122),
.B(n_128),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_174),
.A2(n_175),
.B(n_195),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_122),
.B(n_123),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_180),
.B(n_181),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_141),
.B(n_123),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_119),
.C(n_129),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_30),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_118),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_144),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_196),
.B1(n_28),
.B2(n_27),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_30),
.B(n_16),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_143),
.A2(n_167),
.B1(n_164),
.B2(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_199),
.A2(n_172),
.B1(n_201),
.B2(n_190),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_229),
.Y(n_251)
);

NAND2x1_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_34),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_206),
.A2(n_211),
.B(n_232),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_221),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_208),
.B(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_34),
.B1(n_28),
.B2(n_27),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_195),
.B(n_198),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_34),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_220),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_27),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_192),
.A2(n_25),
.B1(n_26),
.B2(n_9),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_179),
.B(n_5),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_181),
.A2(n_26),
.B(n_25),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_179),
.C(n_172),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_248),
.C(n_229),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_178),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_209),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_173),
.C(n_188),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_249),
.A2(n_220),
.B1(n_218),
.B2(n_222),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_173),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_254),
.B1(n_194),
.B2(n_211),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_212),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_185),
.B1(n_176),
.B2(n_200),
.Y(n_273)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_260),
.Y(n_282)
);

XOR2x2_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_206),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_255),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_206),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_217),
.C(n_221),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_210),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_232),
.C(n_227),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_246),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_211),
.C(n_188),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_228),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_185),
.Y(n_275)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_284),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_254),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_289),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_280),
.B1(n_239),
.B2(n_290),
.Y(n_300)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_263),
.C(n_260),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_258),
.C(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_278),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_271),
.B1(n_252),
.B2(n_239),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_296),
.B(n_237),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_270),
.C(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_298),
.C(n_282),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_277),
.C(n_241),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_236),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_255),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_306),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_222),
.B1(n_247),
.B2(n_237),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_282),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_314),
.C(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_171),
.Y(n_315)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_303),
.B(n_307),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_317),
.B(n_311),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_323),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_309),
.A2(n_304),
.B1(n_246),
.B2(n_249),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_298),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_314),
.C(n_310),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_318),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_329),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_322),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_328),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

OAI321xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_330),
.A3(n_321),
.B1(n_327),
.B2(n_310),
.C(n_176),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_177),
.C(n_213),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_306),
.B(n_9),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_8),
.Y(n_337)
);


endmodule