module fake_jpeg_2853_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AOI21xp33_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_4),
.B(n_0),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_20),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_0),
.B(n_3),
.C(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_15),
.A2(n_11),
.B1(n_12),
.B2(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_18),
.C(n_16),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_35),
.B1(n_29),
.B2(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_37),
.Y(n_43)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_35),
.B(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_42),
.C(n_39),
.Y(n_45)
);


endmodule