module fake_jpeg_10359_n_230 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_20),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_56),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_20),
.B1(n_17),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_26),
.B1(n_18),
.B2(n_29),
.Y(n_89)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_60),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_23),
.C(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_4),
.Y(n_97)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_34),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_2),
.B(n_4),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_2),
.B(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_93),
.B1(n_76),
.B2(n_97),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_81),
.B1(n_93),
.B2(n_5),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_90),
.Y(n_115)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_39),
.B1(n_46),
.B2(n_36),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_89),
.B1(n_57),
.B2(n_30),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_46),
.B1(n_36),
.B2(n_18),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_80),
.A3(n_72),
.B1(n_71),
.B2(n_74),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_36),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_59),
.C(n_47),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_125),
.C(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_57),
.B1(n_18),
.B2(n_29),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_136)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_72),
.B(n_80),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_53),
.B1(n_30),
.B2(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_89),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_47),
.C(n_30),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_132),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_125),
.B(n_105),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_137),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_83),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_145),
.C(n_102),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_76),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_79),
.Y(n_145)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_103),
.B(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_157),
.B(n_132),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_102),
.B(n_107),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_160),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_164),
.C(n_168),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_85),
.B1(n_75),
.B2(n_91),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_144),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_107),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_123),
.B1(n_99),
.B2(n_85),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_133),
.B1(n_139),
.B2(n_137),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_114),
.C(n_78),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_138),
.B1(n_131),
.B2(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_180),
.B1(n_182),
.B2(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_175),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_167),
.B1(n_160),
.B2(n_158),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_140),
.C(n_128),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_150),
.C(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_134),
.B1(n_136),
.B2(n_126),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_127),
.B1(n_135),
.B2(n_147),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_153),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_164),
.C(n_155),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_168),
.C(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_151),
.C(n_157),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_152),
.Y(n_196)
);

AOI321xp33_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_185),
.A3(n_184),
.B1(n_183),
.B2(n_178),
.C(n_181),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_174),
.B1(n_173),
.B2(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_202),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_189),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_186),
.A2(n_175),
.B(n_179),
.Y(n_202)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_183),
.A3(n_170),
.B1(n_161),
.B2(n_148),
.C1(n_146),
.C2(n_30),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_91),
.B(n_92),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_170),
.B(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_5),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_75),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_191),
.C(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_204),
.C(n_201),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_SL g209 ( 
.A1(n_206),
.A2(n_146),
.A3(n_13),
.B(n_15),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_212),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_205),
.B1(n_12),
.B2(n_15),
.C(n_14),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_218),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_213),
.Y(n_218)
);

OAI321xp33_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_14),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_207),
.B(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_223),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_6),
.B(n_9),
.C(n_10),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_6),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_225),
.B(n_217),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_6),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_10),
.C(n_11),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_11),
.Y(n_230)
);


endmodule