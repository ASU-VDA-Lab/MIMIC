module fake_netlist_1_11662_n_946 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_946);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_946;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_786;
wire n_857;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_638;
wire n_563;
wire n_540;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_771;
wire n_735;
wire n_696;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_805;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_875;
wire n_339;
wire n_657;
wire n_583;
wire n_728;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_831;
wire n_602;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g109 ( .A(n_33), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_57), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_97), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_22), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_55), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_9), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_4), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_25), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_14), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_70), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_24), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_26), .Y(n_124) );
NOR2xp67_ASAP7_75t_L g125 ( .A(n_15), .B(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_104), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_39), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_102), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_37), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_66), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_38), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_93), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_62), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_40), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_86), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_46), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_92), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_9), .Y(n_139) );
NOR2xp67_ASAP7_75t_L g140 ( .A(n_81), .B(n_35), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_100), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_15), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_4), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_10), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_5), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_44), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_108), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_8), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
OAI22x1_ASAP7_75t_L g151 ( .A1(n_120), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_110), .B(n_1), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_110), .B(n_2), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_120), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_113), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_139), .B(n_3), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_113), .Y(n_163) );
INVxp67_ASAP7_75t_L g164 ( .A(n_142), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_124), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_139), .B(n_6), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_142), .B(n_7), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_134), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_117), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_144), .B(n_7), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_121), .B(n_8), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_121), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_157), .B(n_112), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_174), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_150), .B(n_119), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_174), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_157), .B(n_164), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_160), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_174), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
NAND2xp33_ASAP7_75t_L g184 ( .A(n_154), .B(n_118), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_174), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_172), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_157), .B(n_123), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_172), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_172), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_157), .B(n_127), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_154), .B(n_143), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_155), .B(n_149), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_132), .B1(n_131), .B2(n_146), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_155), .B(n_133), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_152), .B(n_126), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_158), .B(n_135), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_158), .B(n_136), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_161), .B(n_122), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_161), .B(n_137), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
NOR2x1p5_ASAP7_75t_L g211 ( .A(n_156), .B(n_168), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_171), .B(n_138), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_156), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
AND3x2_ASAP7_75t_L g216 ( .A(n_168), .B(n_144), .C(n_146), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
INVxp33_ASAP7_75t_SL g222 ( .A(n_166), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_167), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_222), .B(n_214), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_215), .B(n_166), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_214), .B(n_141), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_215), .B(n_147), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_220), .B(n_173), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_177), .B(n_151), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_185), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_195), .Y(n_235) );
NAND3xp33_ASAP7_75t_L g236 ( .A(n_204), .B(n_170), .C(n_169), .Y(n_236) );
AO221x1_ASAP7_75t_L g237 ( .A1(n_201), .A2(n_151), .B1(n_122), .B2(n_130), .C(n_145), .Y(n_237) );
NOR2xp33_ASAP7_75t_R g238 ( .A(n_177), .B(n_10), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_216), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_211), .B(n_125), .Y(n_240) );
INVxp33_ASAP7_75t_L g241 ( .A(n_198), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_195), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_220), .B(n_109), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_199), .B(n_128), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_202), .B(n_128), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_179), .B(n_175), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_210), .B(n_129), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_191), .B(n_129), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_210), .B(n_130), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_211), .B(n_145), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_190), .B(n_148), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_190), .A2(n_170), .B1(n_169), .B2(n_167), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_192), .B(n_148), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_184), .B(n_170), .C(n_169), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_192), .B(n_167), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_208), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_193), .B(n_169), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_194), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g261 ( .A1(n_208), .A2(n_170), .B1(n_169), .B2(n_140), .C(n_14), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_197), .B(n_207), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_203), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_193), .A2(n_11), .B(n_12), .C(n_13), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_185), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_194), .B(n_170), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_194), .B(n_11), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_194), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_203), .B(n_13), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_185), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_203), .B(n_63), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_209), .B(n_61), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_200), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_206), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g277 ( .A1(n_201), .A2(n_16), .B(n_17), .C(n_18), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
INVx8_ASAP7_75t_L g279 ( .A(n_225), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_200), .B(n_19), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_200), .B(n_19), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_225), .B(n_20), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_176), .B(n_68), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_176), .B(n_67), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_225), .B(n_69), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_225), .B(n_20), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_226), .B(n_21), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_178), .B(n_23), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_178), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_181), .B(n_189), .C(n_226), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_255), .A2(n_181), .B(n_189), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_233), .B(n_27), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_260), .B(n_226), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_228), .A2(n_226), .B(n_224), .C(n_223), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_238), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_227), .A2(n_224), .B1(n_223), .B2(n_221), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_260), .A2(n_224), .B(n_223), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_270), .B(n_221), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_241), .B(n_248), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_241), .B(n_221), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_263), .B(n_219), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_274), .B(n_219), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_240), .A2(n_219), .B1(n_218), .B2(n_217), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_240), .B(n_218), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_269), .A2(n_218), .B(n_217), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_269), .A2(n_217), .B(n_213), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_267), .A2(n_213), .B(n_205), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_270), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_238), .B(n_213), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_252), .B(n_205), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_255), .A2(n_205), .B(n_196), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_232), .A2(n_196), .B1(n_188), .B2(n_187), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_235), .A2(n_196), .B(n_188), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_250), .B(n_188), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_230), .B(n_187), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_245), .B(n_187), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_229), .B(n_186), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_280), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_280), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_253), .A2(n_186), .B(n_183), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_257), .A2(n_186), .B(n_183), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_268), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_246), .B(n_183), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_242), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_275), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_247), .B(n_182), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_249), .A2(n_182), .B(n_180), .C(n_31), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_259), .A2(n_182), .B(n_180), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_251), .B(n_28), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_237), .B(n_244), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_277), .B(n_107), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_276), .A2(n_30), .B1(n_32), .B2(n_34), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_273), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_264), .B(n_105), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_289), .A2(n_36), .B(n_41), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_236), .A2(n_42), .B(n_43), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_265), .B(n_45), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_297), .A2(n_272), .B(n_288), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_314), .A2(n_272), .B(n_288), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_309), .B(n_279), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_327), .B(n_279), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_337), .A2(n_283), .B(n_284), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_306), .A2(n_283), .B(n_284), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_266), .B(n_234), .Y(n_347) );
OAI22x1_ASAP7_75t_L g348 ( .A1(n_295), .A2(n_256), .B1(n_261), .B2(n_281), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_317), .A2(n_271), .B(n_234), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_323), .A2(n_271), .B(n_243), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_321), .A2(n_286), .B1(n_282), .B2(n_254), .Y(n_352) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_301), .A2(n_285), .B(n_287), .C(n_278), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_293), .A2(n_266), .B(n_262), .Y(n_354) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_315), .B(n_275), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_293), .A2(n_262), .B(n_243), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
OAI21x1_ASAP7_75t_SL g358 ( .A1(n_333), .A2(n_278), .B(n_231), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_326), .A2(n_231), .B(n_275), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_340), .A2(n_275), .B1(n_48), .B2(n_49), .C(n_50), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_312), .A2(n_47), .B(n_51), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_325), .B(n_322), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_315), .B(n_52), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_308), .A2(n_53), .B(n_54), .Y(n_364) );
BUFx10_ASAP7_75t_L g365 ( .A(n_300), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_294), .A2(n_56), .B(n_58), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_330), .A2(n_59), .B(n_60), .Y(n_367) );
OAI21x1_ASAP7_75t_L g368 ( .A1(n_324), .A2(n_65), .B(n_71), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_331), .A2(n_72), .B(n_73), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_320), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_340), .A2(n_74), .B(n_75), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_339), .A2(n_76), .B(n_77), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_358), .A2(n_338), .B(n_332), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_372), .A2(n_298), .B(n_335), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_353), .A2(n_319), .B(n_298), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_350), .A2(n_292), .B(n_319), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_370), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_366), .A2(n_367), .B(n_342), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_357), .B(n_334), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_361), .Y(n_381) );
AOI21x1_ASAP7_75t_L g382 ( .A1(n_341), .A2(n_310), .B(n_313), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_351), .B(n_301), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_345), .A2(n_328), .B(n_290), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_355), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_367), .A2(n_291), .B(n_318), .Y(n_386) );
AOI22x1_ASAP7_75t_L g387 ( .A1(n_348), .A2(n_336), .B1(n_320), .B2(n_304), .Y(n_387) );
AO31x2_ASAP7_75t_L g388 ( .A1(n_352), .A2(n_311), .A3(n_302), .B(n_329), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_343), .B(n_300), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_370), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_366), .B(n_311), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_368), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_344), .B(n_362), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_316), .B(n_296), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_346), .A2(n_302), .B(n_79), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_371), .A2(n_78), .B(n_80), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_371), .A2(n_352), .B(n_359), .Y(n_399) );
CKINVDCx11_ASAP7_75t_R g400 ( .A(n_365), .Y(n_400) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_349), .A2(n_82), .B(n_83), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_363), .Y(n_402) );
AO21x1_ASAP7_75t_L g403 ( .A1(n_363), .A2(n_85), .B(n_87), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_380), .A2(n_360), .B1(n_362), .B2(n_344), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_388), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_394), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_378), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_394), .Y(n_408) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_397), .A2(n_360), .B(n_356), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_402), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_394), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_373), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_400), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_380), .A2(n_365), .B1(n_303), .B2(n_354), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_389), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_400), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_378), .B(n_88), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_380), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_373), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_373), .Y(n_432) );
OAI21x1_ASAP7_75t_L g433 ( .A1(n_397), .A2(n_98), .B(n_99), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
BUFx2_ASAP7_75t_R g438 ( .A(n_398), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_392), .B(n_101), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_392), .A2(n_376), .B(n_386), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_373), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_373), .Y(n_442) );
AOI21x1_ASAP7_75t_L g443 ( .A1(n_393), .A2(n_395), .B(n_381), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_383), .B(n_390), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
INVx3_ASAP7_75t_SL g447 ( .A(n_385), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_390), .B(n_376), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_385), .A2(n_387), .B1(n_403), .B2(n_399), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_399), .B(n_387), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_385), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_423), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_406), .B(n_399), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_423), .B(n_399), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_406), .A2(n_385), .B1(n_398), .B2(n_399), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_408), .B(n_379), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_408), .B(n_385), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_412), .B(n_379), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_412), .B(n_379), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_429), .B(n_385), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_443), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_445), .B(n_398), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_417), .A2(n_375), .B1(n_386), .B2(n_395), .C1(n_393), .C2(n_397), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_443), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_429), .B(n_379), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_445), .B(n_398), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_404), .A2(n_398), .B1(n_379), .B2(n_401), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_436), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_410), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_437), .B(n_401), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_437), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_405), .B(n_401), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_421), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_413), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_421), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_405), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_424), .B(n_401), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_411), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_415), .B(n_386), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_448), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_413), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_413), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_448), .B(n_377), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_422), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_427), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_444), .B(n_377), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_427), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_434), .B(n_375), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_434), .B(n_375), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_418), .B(n_382), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_435), .B(n_384), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_419), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_377), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_435), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_419), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_435), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_410), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_422), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_411), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_410), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_404), .A2(n_377), .B1(n_395), .B2(n_393), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_410), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_441), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_419), .Y(n_514) );
INVx5_ASAP7_75t_L g515 ( .A(n_416), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_441), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_416), .B(n_377), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_447), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_451), .B(n_384), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_447), .B(n_384), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_420), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_451), .B(n_381), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_451), .B(n_381), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_420), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_420), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_447), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_428), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_440), .B(n_396), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_428), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_428), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_425), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_440), .B(n_396), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_432), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_456), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_479), .B(n_439), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_482), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_459), .B(n_432), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_482), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_490), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_490), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
AND2x4_ASAP7_75t_SL g542 ( .A(n_498), .B(n_439), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_459), .B(n_432), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_479), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_491), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_506), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_491), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_484), .B(n_442), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_518), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_461), .B(n_442), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_518), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_502), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_481), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_483), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_484), .B(n_442), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_461), .B(n_452), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_476), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_453), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_494), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_500), .B(n_439), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_453), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_498), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_489), .A2(n_452), .B1(n_446), .B2(n_426), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_462), .B(n_446), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_462), .B(n_450), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_454), .B(n_450), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_454), .B(n_449), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_496), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_502), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_489), .A2(n_425), .B1(n_409), .B2(n_430), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_471), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_471), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_472), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_472), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_519), .B(n_433), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_505), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_514), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_473), .B(n_438), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_473), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_524), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_474), .B(n_438), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_474), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_529), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_488), .B(n_425), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_478), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_529), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_425), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_478), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_480), .B(n_409), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_493), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_519), .B(n_433), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_493), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_480), .B(n_409), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_477), .B(n_409), .Y(n_600) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_458), .B(n_409), .C(n_396), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_530), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_477), .B(n_433), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_513), .B(n_396), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_513), .B(n_396), .Y(n_605) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_504), .B(n_414), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_530), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_516), .B(n_382), .Y(n_608) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_486), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_522), .B(n_523), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_508), .B(n_374), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g612 ( .A(n_515), .B(n_374), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_526), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_516), .B(n_374), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_508), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_521), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_531), .B(n_512), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_527), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_527), .Y(n_620) );
CKINVDCx6p67_ASAP7_75t_R g621 ( .A(n_515), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_503), .B(n_532), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_503), .B(n_532), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_528), .B(n_517), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_533), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_533), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_525), .Y(n_627) );
BUFx3_ASAP7_75t_L g628 ( .A(n_515), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_468), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_528), .B(n_517), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_464), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_515), .B(n_526), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_460), .B(n_475), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_468), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_464), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_467), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_467), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_463), .B(n_509), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_463), .B(n_523), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_486), .B(n_509), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_629), .B(n_455), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_544), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_544), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_622), .B(n_507), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_622), .B(n_507), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_639), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_550), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_623), .B(n_475), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_550), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_549), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_561), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_554), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_639), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_623), .B(n_510), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_546), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_561), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_624), .B(n_495), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_624), .B(n_510), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_554), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_630), .B(n_512), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_629), .B(n_455), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_555), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_546), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_630), .B(n_515), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_613), .B(n_515), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_534), .B(n_487), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_555), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_610), .B(n_520), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_610), .B(n_520), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_634), .B(n_465), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_610), .B(n_522), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_610), .B(n_522), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_549), .B(n_522), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_552), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_634), .B(n_495), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_541), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_628), .B(n_497), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_552), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_628), .B(n_499), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_568), .B(n_469), .Y(n_680) );
AND2x4_ASAP7_75t_SL g681 ( .A(n_621), .B(n_525), .Y(n_681) );
AND2x4_ASAP7_75t_L g682 ( .A(n_628), .B(n_501), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_541), .B(n_525), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_617), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_559), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_606), .B(n_485), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_638), .B(n_492), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_621), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_557), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_633), .B(n_525), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_557), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_617), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_618), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_596), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_596), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_598), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_568), .B(n_492), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_562), .B(n_485), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_625), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_640), .B(n_525), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_565), .B(n_470), .C(n_466), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_625), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_570), .B(n_511), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_618), .B(n_564), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_558), .B(n_566), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_609), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_598), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_558), .B(n_566), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_615), .Y(n_709) );
OR2x6_ASAP7_75t_L g710 ( .A(n_632), .B(n_612), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_615), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_564), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_567), .B(n_537), .Y(n_713) );
NOR3x1_ASAP7_75t_L g714 ( .A(n_606), .B(n_535), .C(n_601), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_567), .B(n_537), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_543), .B(n_551), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_560), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_618), .B(n_576), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_560), .B(n_578), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_543), .B(n_551), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_601), .B(n_585), .C(n_577), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_564), .Y(n_722) );
NAND2x1p5_ASAP7_75t_L g723 ( .A(n_576), .B(n_593), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_563), .B(n_588), .C(n_578), .Y(n_724) );
AND2x4_ASAP7_75t_SL g725 ( .A(n_576), .B(n_626), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_583), .B(n_587), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_563), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_626), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_583), .B(n_587), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_569), .B(n_542), .Y(n_730) );
AND2x4_ASAP7_75t_SL g731 ( .A(n_616), .B(n_620), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_573), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_548), .B(n_556), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_573), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_542), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_575), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_575), .B(n_591), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_612), .B(n_590), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_548), .B(n_556), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_577), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_585), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_588), .B(n_591), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_594), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_594), .B(n_619), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_536), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_616), .B(n_620), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_619), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_614), .B(n_579), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_650), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_713), .B(n_569), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_742), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_720), .B(n_595), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_680), .B(n_600), .Y(n_753) );
OR2x6_ASAP7_75t_L g754 ( .A(n_710), .B(n_590), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_742), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_668), .B(n_595), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_685), .B(n_572), .C(n_636), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_719), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_719), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_669), .B(n_599), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_648), .B(n_599), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_657), .B(n_536), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_651), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_737), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_715), .B(n_538), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_676), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_651), .Y(n_767) );
OA211x2_ASAP7_75t_L g768 ( .A1(n_685), .A2(n_611), .B(n_542), .C(n_593), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_737), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_676), .Y(n_770) );
INVx3_ASAP7_75t_L g771 ( .A(n_710), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_705), .B(n_614), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_654), .B(n_597), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_716), .B(n_538), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_705), .B(n_600), .Y(n_775) );
OR2x2_ASAP7_75t_L g776 ( .A(n_708), .B(n_539), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_731), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_746), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_708), .B(n_539), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_698), .B(n_605), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_644), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_744), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_658), .B(n_597), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_744), .Y(n_784) );
AND2x4_ASAP7_75t_SL g785 ( .A(n_693), .B(n_540), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_642), .Y(n_786) );
INVx1_ASAP7_75t_SL g787 ( .A(n_725), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_748), .B(n_597), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_698), .B(n_605), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_733), .B(n_540), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_646), .B(n_597), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_748), .B(n_579), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_643), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_688), .Y(n_794) );
NOR2x1p5_ASAP7_75t_SL g795 ( .A(n_703), .B(n_637), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_739), .B(n_545), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_680), .B(n_604), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_645), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g799 ( .A1(n_693), .A2(n_579), .B(n_603), .C(n_604), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_647), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_649), .Y(n_801) );
AOI32xp33_ASAP7_75t_L g802 ( .A1(n_726), .A2(n_579), .A3(n_603), .B1(n_608), .B2(n_635), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_653), .B(n_545), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_687), .B(n_547), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_652), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_730), .B(n_608), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_660), .B(n_547), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_675), .B(n_636), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_697), .B(n_553), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_659), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_697), .B(n_635), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_662), .Y(n_812) );
OAI21xp33_ASAP7_75t_SL g813 ( .A1(n_710), .A2(n_553), .B(n_571), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_671), .B(n_571), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_686), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_656), .Y(n_816) );
OR2x2_ASAP7_75t_L g817 ( .A(n_641), .B(n_574), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_641), .B(n_574), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_656), .Y(n_819) );
OR2x2_ASAP7_75t_L g820 ( .A(n_661), .B(n_580), .Y(n_820) );
OAI21xp5_ASAP7_75t_L g821 ( .A1(n_701), .A2(n_637), .B(n_631), .Y(n_821) );
INVx2_ASAP7_75t_SL g822 ( .A(n_664), .Y(n_822) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_678), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_701), .B(n_631), .C(n_581), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_661), .B(n_580), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_667), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_689), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_670), .B(n_581), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_729), .B(n_678), .Y(n_829) );
OR2x2_ASAP7_75t_L g830 ( .A(n_675), .B(n_582), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_821), .B(n_666), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_758), .Y(n_832) );
INVx1_ASAP7_75t_SL g833 ( .A(n_794), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_815), .B(n_787), .Y(n_834) );
AND2x4_ASAP7_75t_L g835 ( .A(n_771), .B(n_714), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_829), .A2(n_673), .B1(n_670), .B2(n_738), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_821), .B(n_747), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_759), .Y(n_838) );
AOI21xp33_ASAP7_75t_L g839 ( .A1(n_824), .A2(n_721), .B(n_706), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_765), .B(n_663), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_764), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_830), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_761), .B(n_672), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_766), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_768), .A2(n_682), .B1(n_690), .B2(n_706), .Y(n_845) );
NAND2x1p5_ASAP7_75t_L g846 ( .A(n_787), .B(n_735), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_750), .B(n_655), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_769), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_768), .A2(n_677), .B1(n_679), .B2(n_682), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_782), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_770), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_784), .Y(n_852) );
AND2x4_ASAP7_75t_L g853 ( .A(n_771), .B(n_718), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_824), .B(n_717), .Y(n_854) );
OAI32xp33_ASAP7_75t_L g855 ( .A1(n_813), .A2(n_777), .A3(n_823), .B1(n_819), .B2(n_816), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_753), .B(n_696), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_776), .Y(n_857) );
NAND2xp5_ASAP7_75t_SL g858 ( .A(n_813), .B(n_718), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_778), .B(n_674), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_751), .A2(n_679), .B1(n_677), .B2(n_683), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_756), .B(n_665), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_779), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_775), .B(n_704), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_811), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_811), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_753), .B(n_691), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_763), .Y(n_867) );
BUFx3_ASAP7_75t_L g868 ( .A(n_785), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_828), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_755), .B(n_704), .Y(n_870) );
AO32x1_ASAP7_75t_L g871 ( .A1(n_749), .A2(n_681), .A3(n_743), .B1(n_741), .B2(n_740), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_828), .Y(n_872) );
NAND4xp75_ASAP7_75t_L g873 ( .A(n_795), .B(n_709), .C(n_736), .D(n_734), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_767), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_780), .B(n_707), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_760), .B(n_712), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_786), .Y(n_877) );
OAI22x1_ASAP7_75t_L g878 ( .A1(n_788), .A2(n_723), .B1(n_722), .B2(n_721), .Y(n_878) );
OAI321xp33_ASAP7_75t_L g879 ( .A1(n_846), .A2(n_802), .A3(n_754), .B1(n_757), .B2(n_799), .C(n_723), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_846), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_869), .Y(n_881) );
OAI31xp33_ASAP7_75t_L g882 ( .A1(n_833), .A2(n_757), .A3(n_792), .B(n_788), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_835), .A2(n_754), .B1(n_792), .B2(n_822), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_858), .A2(n_754), .B1(n_789), .B2(n_797), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_835), .B(n_752), .Y(n_885) );
AOI21xp33_ASAP7_75t_L g886 ( .A1(n_833), .A2(n_827), .B(n_826), .Y(n_886) );
O2A1O1Ixp33_ASAP7_75t_SL g887 ( .A1(n_855), .A2(n_834), .B(n_839), .C(n_845), .Y(n_887) );
XOR2x2_ASAP7_75t_L g888 ( .A(n_868), .B(n_773), .Y(n_888) );
AOI222xp33_ASAP7_75t_L g889 ( .A1(n_878), .A2(n_812), .B1(n_810), .B2(n_793), .C1(n_805), .C2(n_800), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_839), .B(n_808), .C(n_801), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_870), .A2(n_853), .B1(n_831), .B2(n_857), .Y(n_891) );
OAI22xp33_ASAP7_75t_SL g892 ( .A1(n_836), .A2(n_774), .B1(n_772), .B2(n_797), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_844), .Y(n_893) );
OR2x2_ASAP7_75t_L g894 ( .A(n_862), .B(n_809), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_856), .B(n_762), .Y(n_895) );
AND2x4_ASAP7_75t_L g896 ( .A(n_853), .B(n_783), .Y(n_896) );
OR2x2_ASAP7_75t_L g897 ( .A(n_856), .B(n_804), .Y(n_897) );
AOI221x1_ASAP7_75t_L g898 ( .A1(n_851), .A2(n_825), .B1(n_724), .B2(n_798), .C(n_781), .Y(n_898) );
NAND3xp33_ASAP7_75t_L g899 ( .A(n_854), .B(n_825), .C(n_724), .Y(n_899) );
OAI33xp33_ASAP7_75t_L g900 ( .A1(n_872), .A2(n_820), .A3(n_818), .B1(n_817), .B2(n_796), .B3(n_790), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_876), .B(n_861), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_863), .A2(n_791), .B1(n_807), .B2(n_803), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_843), .B(n_814), .Y(n_903) );
OAI32xp33_ASAP7_75t_L g904 ( .A1(n_849), .A2(n_806), .A3(n_700), .B1(n_694), .B2(n_695), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_900), .A2(n_864), .B1(n_865), .B2(n_838), .C(n_852), .Y(n_905) );
OA22x2_ASAP7_75t_L g906 ( .A1(n_898), .A2(n_860), .B1(n_842), .B2(n_875), .Y(n_906) );
NAND2x1_ASAP7_75t_L g907 ( .A(n_879), .B(n_871), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_892), .B(n_848), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_900), .A2(n_850), .B1(n_841), .B2(n_832), .Y(n_909) );
OAI221xp5_ASAP7_75t_L g910 ( .A1(n_882), .A2(n_837), .B1(n_854), .B2(n_866), .C(n_859), .Y(n_910) );
NAND4xp25_ASAP7_75t_L g911 ( .A(n_887), .B(n_837), .C(n_866), .D(n_877), .Y(n_911) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_884), .Y(n_912) );
AOI222xp33_ASAP7_75t_L g913 ( .A1(n_879), .A2(n_867), .B1(n_874), .B2(n_847), .C1(n_732), .C2(n_727), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_902), .A2(n_883), .B1(n_891), .B2(n_896), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g915 ( .A(n_889), .B(n_840), .C(n_871), .D(n_711), .Y(n_915) );
AOI211x1_ASAP7_75t_L g916 ( .A1(n_904), .A2(n_871), .B(n_873), .C(n_684), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_889), .A2(n_728), .B1(n_702), .B2(n_699), .C(n_692), .Y(n_917) );
NOR3xp33_ASAP7_75t_L g918 ( .A(n_890), .B(n_745), .C(n_584), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_913), .B(n_899), .C(n_886), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_912), .A2(n_880), .B1(n_888), .B2(n_885), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_914), .B(n_896), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_911), .B(n_886), .Y(n_922) );
INVxp67_ASAP7_75t_SL g923 ( .A(n_918), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_909), .B(n_881), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_906), .A2(n_902), .B1(n_893), .B2(n_901), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_910), .A2(n_894), .B1(n_897), .B2(n_895), .Y(n_926) );
NOR3xp33_ASAP7_75t_L g927 ( .A(n_919), .B(n_907), .C(n_915), .Y(n_927) );
NAND4xp25_ASAP7_75t_L g928 ( .A(n_920), .B(n_916), .C(n_908), .D(n_917), .Y(n_928) );
NOR3xp33_ASAP7_75t_L g929 ( .A(n_922), .B(n_905), .C(n_903), .Y(n_929) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_923), .Y(n_930) );
AND2x4_ASAP7_75t_L g931 ( .A(n_930), .B(n_921), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_927), .Y(n_932) );
NOR2xp67_ASAP7_75t_L g933 ( .A(n_928), .B(n_925), .Y(n_933) );
NOR3xp33_ASAP7_75t_L g934 ( .A(n_932), .B(n_929), .C(n_924), .Y(n_934) );
OR2x2_ASAP7_75t_L g935 ( .A(n_931), .B(n_926), .Y(n_935) );
OAI22x1_ASAP7_75t_L g936 ( .A1(n_935), .A2(n_931), .B1(n_933), .B2(n_586), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_934), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_936), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_937), .A2(n_627), .B1(n_584), .B2(n_586), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_938), .A2(n_627), .B1(n_589), .B2(n_592), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_940), .Y(n_941) );
OR2x2_ASAP7_75t_L g942 ( .A(n_941), .B(n_939), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g943 ( .A1(n_942), .A2(n_627), .B1(n_589), .B2(n_592), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_943), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_944), .A2(n_627), .B1(n_602), .B2(n_607), .C(n_582), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_945), .A2(n_627), .B1(n_602), .B2(n_607), .Y(n_946) );
endmodule