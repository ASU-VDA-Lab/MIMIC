module fake_jpeg_3696_n_117 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_39),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_41),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_34),
.B(n_37),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_44),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_33),
.B1(n_32),
.B2(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_33),
.B1(n_32),
.B2(n_43),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_64),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_68),
.B1(n_1),
.B2(n_3),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_49),
.B(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_50),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_33),
.B1(n_42),
.B2(n_2),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_76),
.C(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_0),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_1),
.B(n_3),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_4),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_74),
.C(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_5),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_87),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_30),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_9),
.B(n_11),
.C(n_13),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_19),
.B(n_20),
.C(n_24),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_14),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_101),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_88),
.C(n_83),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_97),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_91),
.B(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_110),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_105),
.C(n_104),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_102),
.C(n_26),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_107),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_111),
.B(n_28),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_25),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_29),
.Y(n_117)
);


endmodule