module real_aes_7616_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_725;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_1), .A2(n_154), .B(n_159), .C(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_2), .A2(n_149), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g468 ( .A(n_3), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_4), .B(n_173), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_5), .A2(n_105), .B1(n_119), .B2(n_743), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_6), .A2(n_17), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_6), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g485 ( .A1(n_7), .A2(n_149), .B(n_486), .Y(n_485) );
AND2x6_ASAP7_75t_L g154 ( .A(n_8), .B(n_155), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_9), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_9), .Y(n_730) );
INVx1_ASAP7_75t_L g183 ( .A(n_10), .Y(n_183) );
INVx1_ASAP7_75t_L g111 ( .A(n_11), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_11), .B(n_45), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_12), .A2(n_261), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_13), .B(n_164), .Y(n_200) );
INVx1_ASAP7_75t_L g490 ( .A(n_14), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_15), .B(n_163), .Y(n_538) );
INVx1_ASAP7_75t_L g147 ( .A(n_16), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_17), .Y(n_735) );
INVx1_ASAP7_75t_L g550 ( .A(n_18), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_19), .A2(n_184), .B(n_209), .C(n_211), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_20), .B(n_173), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_21), .B(n_479), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_22), .B(n_149), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_23), .B(n_269), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_24), .A2(n_163), .B(n_165), .C(n_169), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_25), .A2(n_49), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_25), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_25), .B(n_173), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_26), .B(n_164), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_27), .A2(n_167), .B(n_211), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_28), .B(n_164), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_29), .Y(n_229) );
INVx1_ASAP7_75t_L g243 ( .A(n_30), .Y(n_243) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_31), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_32), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_33), .B(n_164), .Y(n_469) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_34), .A2(n_454), .B1(n_728), .B2(n_729), .C1(n_738), .C2(n_739), .Y(n_453) );
INVx1_ASAP7_75t_L g266 ( .A(n_35), .Y(n_266) );
INVx1_ASAP7_75t_L g503 ( .A(n_36), .Y(n_503) );
INVx2_ASAP7_75t_L g152 ( .A(n_37), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_38), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_39), .A2(n_163), .B(n_222), .C(n_224), .Y(n_221) );
INVxp67_ASAP7_75t_L g267 ( .A(n_40), .Y(n_267) );
CKINVDCx14_ASAP7_75t_R g220 ( .A(n_41), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_42), .A2(n_159), .B(n_242), .C(n_248), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_43), .A2(n_154), .B(n_159), .C(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_44), .A2(n_93), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_44), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_45), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g502 ( .A(n_46), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_47), .A2(n_181), .B(n_182), .C(n_185), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_48), .B(n_164), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_49), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_50), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_51), .Y(n_263) );
INVx1_ASAP7_75t_L g157 ( .A(n_52), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_53), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_54), .B(n_149), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_55), .A2(n_159), .B1(n_169), .B2(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_56), .B(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_57), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_58), .Y(n_465) );
CKINVDCx14_ASAP7_75t_R g179 ( .A(n_59), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_60), .A2(n_181), .B(n_224), .C(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_61), .Y(n_531) );
INVx1_ASAP7_75t_L g487 ( .A(n_62), .Y(n_487) );
INVx1_ASAP7_75t_L g155 ( .A(n_63), .Y(n_155) );
INVx1_ASAP7_75t_L g146 ( .A(n_64), .Y(n_146) );
INVx1_ASAP7_75t_SL g223 ( .A(n_65), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_66), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_67), .B(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g232 ( .A(n_68), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_SL g478 ( .A1(n_69), .A2(n_224), .B(n_479), .C(n_480), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_70), .Y(n_481) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_72), .A2(n_149), .B(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_73), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_74), .A2(n_149), .B(n_206), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_75), .Y(n_506) );
INVx1_ASAP7_75t_L g525 ( .A(n_76), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_77), .A2(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g207 ( .A(n_78), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_79), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_80), .A2(n_154), .B(n_159), .C(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_81), .A2(n_149), .B(n_156), .Y(n_148) );
INVx1_ASAP7_75t_L g210 ( .A(n_82), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_83), .B(n_244), .Y(n_519) );
INVx2_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
INVx1_ASAP7_75t_L g197 ( .A(n_85), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_86), .B(n_479), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_87), .A2(n_154), .B(n_159), .C(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g115 ( .A(n_88), .Y(n_115) );
OR2x2_ASAP7_75t_L g446 ( .A(n_88), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g727 ( .A(n_88), .B(n_448), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_89), .A2(n_159), .B(n_231), .C(n_234), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_90), .A2(n_733), .B1(n_734), .B2(n_737), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_90), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_91), .B(n_176), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_92), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_93), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_94), .A2(n_154), .B(n_159), .C(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_95), .Y(n_542) );
INVx1_ASAP7_75t_L g477 ( .A(n_96), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_97), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_98), .B(n_244), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_99), .B(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_100), .B(n_142), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_101), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g166 ( .A(n_102), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_103), .A2(n_149), .B(n_476), .Y(n_475) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g745 ( .A(n_108), .Y(n_745) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .C(n_116), .Y(n_113) );
AND2x2_ASAP7_75t_L g448 ( .A(n_114), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g455 ( .A(n_115), .B(n_448), .Y(n_455) );
NOR2x2_ASAP7_75t_L g741 ( .A(n_115), .B(n_447), .Y(n_741) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
AO21x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_125), .B(n_452), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g742 ( .A(n_122), .Y(n_742) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI21xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_444), .B(n_450), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_442), .B2(n_443), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_127), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_130), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_134), .B1(n_440), .B2(n_441), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_131), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_134), .A2(n_455), .B1(n_456), .B2(n_725), .Y(n_454) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g441 ( .A(n_135), .Y(n_441) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_366), .Y(n_135) );
NOR4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_308), .C(n_338), .D(n_348), .Y(n_136) );
OAI211xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_213), .B(n_271), .C(n_298), .Y(n_137) );
OAI222xp33_ASAP7_75t_L g393 ( .A1(n_138), .A2(n_313), .B1(n_394), .B2(n_395), .C1(n_396), .C2(n_397), .Y(n_393) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_188), .Y(n_138) );
AOI33xp33_ASAP7_75t_L g319 ( .A1(n_139), .A2(n_306), .A3(n_307), .B1(n_320), .B2(n_325), .B3(n_327), .Y(n_319) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_139), .A2(n_377), .B(n_379), .C(n_381), .Y(n_376) );
OR2x2_ASAP7_75t_L g392 ( .A(n_139), .B(n_378), .Y(n_392) );
INVx1_ASAP7_75t_L g425 ( .A(n_139), .Y(n_425) );
OR2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_175), .Y(n_139) );
INVx2_ASAP7_75t_L g302 ( .A(n_140), .Y(n_302) );
AND2x2_ASAP7_75t_L g318 ( .A(n_140), .B(n_204), .Y(n_318) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_140), .Y(n_353) );
AND2x2_ASAP7_75t_L g382 ( .A(n_140), .B(n_175), .Y(n_382) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_148), .B(n_172), .Y(n_140) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_141), .A2(n_205), .B(n_212), .Y(n_204) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_141), .A2(n_218), .B(n_226), .Y(n_217) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_142), .A2(n_475), .B(n_482), .Y(n_474) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g259 ( .A(n_143), .Y(n_259) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_144), .B(n_145), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx2_ASAP7_75t_L g261 ( .A(n_149), .Y(n_261) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_150), .B(n_154), .Y(n_194) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g247 ( .A(n_151), .Y(n_247) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
INVx1_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
INVx1_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
INVx3_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx1_ASAP7_75t_L g479 ( .A(n_153), .Y(n_479) );
INVx4_ASAP7_75t_SL g171 ( .A(n_154), .Y(n_171) );
BUFx3_ASAP7_75t_L g248 ( .A(n_154), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_158), .B(n_162), .C(n_171), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g178 ( .A1(n_158), .A2(n_171), .B(n_179), .C(n_180), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g206 ( .A1(n_158), .A2(n_171), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_158), .A2(n_171), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_SL g262 ( .A1(n_158), .A2(n_171), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_158), .A2(n_171), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_158), .A2(n_171), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_158), .A2(n_171), .B(n_547), .C(n_548), .Y(n_546) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx3_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_163), .B(n_223), .Y(n_222) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_167), .B(n_210), .Y(n_209) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_167), .A2(n_244), .B1(n_266), .B2(n_267), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_167), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g501 ( .A1(n_168), .A2(n_199), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g470 ( .A(n_169), .Y(n_470) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g234 ( .A(n_171), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_171), .A2(n_194), .B1(n_500), .B2(n_504), .Y(n_499) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_173), .A2(n_485), .B(n_491), .Y(n_484) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_174), .B(n_203), .Y(n_202) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_174), .A2(n_228), .B(n_235), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_174), .B(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g521 ( .A(n_174), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g282 ( .A(n_175), .Y(n_282) );
BUFx3_ASAP7_75t_L g290 ( .A(n_175), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_175), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g301 ( .A(n_175), .B(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_175), .B(n_189), .Y(n_330) );
AND2x2_ASAP7_75t_L g399 ( .A(n_175), .B(n_333), .Y(n_399) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_187), .Y(n_175) );
INVx1_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
INVx2_ASAP7_75t_L g237 ( .A(n_176), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_176), .A2(n_194), .B(n_240), .C(n_241), .Y(n_239) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_176), .A2(n_545), .B(n_551), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
INVx5_ASAP7_75t_L g244 ( .A(n_184), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_184), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_184), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g201 ( .A(n_185), .Y(n_201) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g211 ( .A(n_186), .Y(n_211) );
INVx2_ASAP7_75t_SL g293 ( .A(n_188), .Y(n_293) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_189), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g335 ( .A(n_189), .Y(n_335) );
AND2x2_ASAP7_75t_L g346 ( .A(n_189), .B(n_302), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_189), .B(n_331), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_189), .B(n_333), .Y(n_378) );
AND2x2_ASAP7_75t_L g437 ( .A(n_189), .B(n_382), .Y(n_437) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g307 ( .A(n_190), .B(n_204), .Y(n_307) );
AND2x2_ASAP7_75t_L g317 ( .A(n_190), .B(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g339 ( .A(n_190), .Y(n_339) );
AND3x2_ASAP7_75t_L g398 ( .A(n_190), .B(n_399), .C(n_400), .Y(n_398) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_202), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_191), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_191), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_191), .B(n_542), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_194), .A2(n_229), .B(n_230), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_194), .A2(n_465), .B(n_466), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_194), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_200), .C(n_201), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_201), .B(n_232), .C(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_201), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_201), .A2(n_528), .B(n_529), .Y(n_527) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_204), .Y(n_289) );
INVx1_ASAP7_75t_SL g333 ( .A(n_204), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_204), .B(n_282), .C(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_251), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_214), .A2(n_317), .B(n_369), .C(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_216), .B(n_238), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_216), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g385 ( .A(n_216), .Y(n_385) );
AND2x2_ASAP7_75t_L g406 ( .A(n_216), .B(n_253), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_216), .B(n_315), .Y(n_434) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
AND2x2_ASAP7_75t_L g279 ( .A(n_217), .B(n_270), .Y(n_279) );
INVx2_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
AND2x2_ASAP7_75t_L g306 ( .A(n_217), .B(n_253), .Y(n_306) );
AND2x2_ASAP7_75t_L g356 ( .A(n_217), .B(n_238), .Y(n_356) );
INVx1_ASAP7_75t_L g360 ( .A(n_217), .Y(n_360) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_225), .Y(n_539) );
INVx2_ASAP7_75t_SL g270 ( .A(n_227), .Y(n_270) );
BUFx2_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
AND2x2_ASAP7_75t_L g423 ( .A(n_227), .B(n_238), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g269 ( .A(n_237), .Y(n_269) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_237), .A2(n_534), .B(n_541), .Y(n_533) );
INVx3_ASAP7_75t_SL g253 ( .A(n_238), .Y(n_253) );
AND2x2_ASAP7_75t_L g278 ( .A(n_238), .B(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g285 ( .A(n_238), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g315 ( .A(n_238), .B(n_275), .Y(n_315) );
OR2x2_ASAP7_75t_L g324 ( .A(n_238), .B(n_270), .Y(n_324) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_238), .Y(n_342) );
AND2x2_ASAP7_75t_L g347 ( .A(n_238), .B(n_300), .Y(n_347) );
AND2x2_ASAP7_75t_L g375 ( .A(n_238), .B(n_255), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_238), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g413 ( .A(n_238), .B(n_254), .Y(n_413) );
OR2x6_ASAP7_75t_L g238 ( .A(n_239), .B(n_249), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_245), .C(n_246), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_244), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_247), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g337 ( .A(n_253), .B(n_286), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_253), .B(n_279), .Y(n_365) );
AND2x2_ASAP7_75t_L g383 ( .A(n_253), .B(n_300), .Y(n_383) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_270), .Y(n_254) );
AND2x2_ASAP7_75t_L g284 ( .A(n_255), .B(n_270), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_255), .B(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
OR2x2_ASAP7_75t_L g370 ( .A(n_255), .B(n_290), .Y(n_370) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_260), .B(n_268), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_257), .A2(n_276), .B(n_277), .Y(n_275) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_257), .A2(n_524), .B(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AOI21xp5_ASAP7_75t_SL g515 ( .A1(n_258), .A2(n_516), .B(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_259), .A2(n_464), .B(n_471), .Y(n_463) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_259), .A2(n_499), .B(n_505), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_259), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g276 ( .A(n_260), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_268), .Y(n_277) );
AND2x2_ASAP7_75t_L g305 ( .A(n_270), .B(n_275), .Y(n_305) );
INVx1_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
AND2x2_ASAP7_75t_L g408 ( .A(n_270), .B(n_286), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_280), .B1(n_283), .B2(n_287), .C1(n_291), .C2(n_294), .Y(n_271) );
INVx1_ASAP7_75t_L g403 ( .A(n_272), .Y(n_403) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
AND2x2_ASAP7_75t_L g299 ( .A(n_273), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g310 ( .A(n_273), .B(n_279), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_273), .B(n_301), .Y(n_326) );
OAI222xp33_ASAP7_75t_L g348 ( .A1(n_273), .A2(n_349), .B1(n_354), .B2(n_355), .C1(n_363), .C2(n_365), .Y(n_348) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g336 ( .A(n_275), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_275), .B(n_356), .Y(n_396) );
AND2x2_ASAP7_75t_L g407 ( .A(n_275), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g415 ( .A(n_278), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_280), .B(n_331), .Y(n_394) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_282), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g352 ( .A(n_282), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx3_ASAP7_75t_L g297 ( .A(n_285), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_285), .A2(n_388), .B(n_391), .C(n_393), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_285), .B(n_322), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_285), .B(n_305), .Y(n_427) );
AND2x2_ASAP7_75t_L g300 ( .A(n_286), .B(n_296), .Y(n_300) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g327 ( .A(n_289), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_290), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g379 ( .A(n_290), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_318), .Y(n_418) );
INVx1_ASAP7_75t_L g430 ( .A(n_290), .Y(n_430) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_293), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g411 ( .A(n_296), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_301), .B(n_303), .C(n_307), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_299), .A2(n_329), .B1(n_344), .B2(n_347), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_300), .B(n_314), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_300), .B(n_322), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_301), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g364 ( .A(n_301), .Y(n_364) );
AND2x2_ASAP7_75t_L g371 ( .A(n_301), .B(n_351), .Y(n_371) );
INVx2_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NOR4xp25_ASAP7_75t_L g309 ( .A(n_306), .B(n_310), .C(n_311), .D(n_314), .Y(n_309) );
INVx1_ASAP7_75t_SL g380 ( .A(n_307), .Y(n_380) );
AND2x2_ASAP7_75t_L g424 ( .A(n_307), .B(n_425), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_316), .B(n_319), .C(n_328), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_315), .B(n_385), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_317), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_435) );
INVx1_ASAP7_75t_SL g390 ( .A(n_318), .Y(n_390) );
AND2x2_ASAP7_75t_L g429 ( .A(n_318), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_322), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_326), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_327), .B(n_352), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_334), .B(n_336), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g404 ( .A(n_331), .Y(n_404) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g432 ( .A(n_332), .Y(n_432) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B(n_343), .Y(n_338) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_339), .Y(n_351) );
OR2x2_ASAP7_75t_L g389 ( .A(n_339), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI21xp33_ASAP7_75t_SL g384 ( .A1(n_342), .A2(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_346), .A2(n_373), .B1(n_376), .B2(n_383), .C(n_384), .Y(n_372) );
INVx1_ASAP7_75t_SL g416 ( .A(n_347), .Y(n_416) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OR2x2_ASAP7_75t_L g363 ( .A(n_351), .B(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g400 ( .A(n_353), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_360), .B2(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_359), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_401), .C(n_414), .D(n_426), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_372), .C(n_387), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_370), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_377), .B(n_382), .Y(n_386) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_389), .A2(n_415), .B1(n_416), .B2(n_417), .C(n_419), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_391), .A2(n_406), .B(n_407), .C(n_409), .Y(n_405) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_392), .A2(n_410), .B1(n_412), .B2(n_413), .Y(n_409) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_404), .C(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g420 ( .A(n_413), .Y(n_420) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI221xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_428), .B1(n_431), .B2(n_433), .C(n_435), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_441), .A2(n_455), .B1(n_457), .B2(n_727), .Y(n_738) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g451 ( .A(n_445), .Y(n_451) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI21xp33_ASAP7_75t_SL g452 ( .A1(n_450), .A2(n_453), .B(n_742), .Y(n_452) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_641), .Y(n_457) );
NOR5xp2_ASAP7_75t_L g458 ( .A(n_459), .B(n_564), .C(n_596), .D(n_611), .E(n_628), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_492), .B(n_511), .C(n_552), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_473), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_461), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_461), .B(n_616), .Y(n_679) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_462), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_462), .B(n_508), .Y(n_565) );
AND2x2_ASAP7_75t_L g606 ( .A(n_462), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_462), .B(n_575), .Y(n_610) );
OR2x2_ASAP7_75t_L g647 ( .A(n_462), .B(n_498), .Y(n_647) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g497 ( .A(n_463), .B(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g555 ( .A(n_463), .Y(n_555) );
OR2x2_ASAP7_75t_L g718 ( .A(n_463), .B(n_558), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_473), .A2(n_621), .B1(n_622), .B2(n_625), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_473), .B(n_555), .Y(n_704) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
AND2x2_ASAP7_75t_L g510 ( .A(n_474), .B(n_498), .Y(n_510) );
AND2x2_ASAP7_75t_L g557 ( .A(n_474), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g562 ( .A(n_474), .Y(n_562) );
INVx3_ASAP7_75t_L g575 ( .A(n_474), .Y(n_575) );
OR2x2_ASAP7_75t_L g595 ( .A(n_474), .B(n_558), .Y(n_595) );
AND2x2_ASAP7_75t_L g614 ( .A(n_474), .B(n_484), .Y(n_614) );
BUFx2_ASAP7_75t_L g646 ( .A(n_474), .Y(n_646) );
AND2x4_ASAP7_75t_L g561 ( .A(n_483), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g496 ( .A(n_484), .Y(n_496) );
INVx2_ASAP7_75t_L g509 ( .A(n_484), .Y(n_509) );
OR2x2_ASAP7_75t_L g577 ( .A(n_484), .B(n_558), .Y(n_577) );
AND2x2_ASAP7_75t_L g607 ( .A(n_484), .B(n_498), .Y(n_607) );
AND2x2_ASAP7_75t_L g624 ( .A(n_484), .B(n_555), .Y(n_624) );
AND2x2_ASAP7_75t_L g664 ( .A(n_484), .B(n_575), .Y(n_664) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_484), .B(n_510), .Y(n_700) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp33_ASAP7_75t_SL g493 ( .A(n_494), .B(n_507), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_495), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_496), .A2(n_510), .B(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_496), .B(n_498), .Y(n_694) );
AND2x2_ASAP7_75t_L g630 ( .A(n_497), .B(n_631), .Y(n_630) );
INVx3_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_498), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_507), .B(n_555), .Y(n_723) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_508), .A2(n_666), .B1(n_667), .B2(n_672), .Y(n_665) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_L g556 ( .A(n_509), .B(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g594 ( .A(n_509), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g631 ( .A(n_509), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_510), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g685 ( .A(n_510), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_532), .Y(n_512) );
INVx4_ASAP7_75t_L g571 ( .A(n_513), .Y(n_571) );
AND2x2_ASAP7_75t_L g649 ( .A(n_513), .B(n_616), .Y(n_649) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
INVx3_ASAP7_75t_L g568 ( .A(n_514), .Y(n_568) );
AND2x2_ASAP7_75t_L g582 ( .A(n_514), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_514), .Y(n_586) );
INVx2_ASAP7_75t_L g600 ( .A(n_514), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_514), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g657 ( .A(n_514), .B(n_652), .Y(n_657) );
AND2x2_ASAP7_75t_L g722 ( .A(n_514), .B(n_692), .Y(n_722) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_521), .Y(n_514) );
AND2x2_ASAP7_75t_L g563 ( .A(n_523), .B(n_544), .Y(n_563) );
INVx2_ASAP7_75t_L g583 ( .A(n_523), .Y(n_583) );
INVx1_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
AND2x2_ASAP7_75t_L g634 ( .A(n_532), .B(n_582), .Y(n_634) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_543), .Y(n_532) );
INVx2_ASAP7_75t_L g573 ( .A(n_533), .Y(n_573) );
INVx1_ASAP7_75t_L g581 ( .A(n_533), .Y(n_581) );
AND2x2_ASAP7_75t_L g599 ( .A(n_533), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_533), .B(n_583), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .Y(n_536) );
AND2x2_ASAP7_75t_L g616 ( .A(n_543), .B(n_573), .Y(n_616) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g569 ( .A(n_544), .Y(n_569) );
AND2x2_ASAP7_75t_L g652 ( .A(n_544), .B(n_583), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_559), .B(n_563), .Y(n_552) );
INVx1_ASAP7_75t_SL g597 ( .A(n_553), .Y(n_597) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_554), .B(n_561), .Y(n_654) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g603 ( .A(n_555), .B(n_558), .Y(n_603) );
AND2x2_ASAP7_75t_L g632 ( .A(n_555), .B(n_576), .Y(n_632) );
OR2x2_ASAP7_75t_L g635 ( .A(n_555), .B(n_595), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_556), .A2(n_648), .B1(n_700), .B2(n_701), .C1(n_703), .C2(n_705), .Y(n_699) );
BUFx2_ASAP7_75t_L g613 ( .A(n_558), .Y(n_613) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g602 ( .A(n_561), .B(n_603), .Y(n_602) );
INVx3_ASAP7_75t_SL g619 ( .A(n_561), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_561), .B(n_613), .Y(n_673) );
AND2x2_ASAP7_75t_L g608 ( .A(n_563), .B(n_568), .Y(n_608) );
INVx1_ASAP7_75t_L g627 ( .A(n_563), .Y(n_627) );
OAI221xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_566), .B1(n_570), .B2(n_574), .C(n_578), .Y(n_564) );
OR2x2_ASAP7_75t_L g636 ( .A(n_566), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g621 ( .A(n_568), .B(n_591), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_568), .B(n_581), .Y(n_661) );
AND2x2_ASAP7_75t_L g666 ( .A(n_568), .B(n_616), .Y(n_666) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_568), .Y(n_676) );
NAND2x1_ASAP7_75t_SL g687 ( .A(n_568), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g572 ( .A(n_569), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g592 ( .A(n_569), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_569), .B(n_587), .Y(n_618) );
INVx1_ASAP7_75t_L g684 ( .A(n_569), .Y(n_684) );
INVx1_ASAP7_75t_L g659 ( .A(n_570), .Y(n_659) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g671 ( .A(n_571), .Y(n_671) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_571), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g688 ( .A(n_572), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_572), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g591 ( .A(n_573), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_573), .B(n_583), .Y(n_604) );
INVx1_ASAP7_75t_L g670 ( .A(n_573), .Y(n_670) );
INVx1_ASAP7_75t_L g691 ( .A(n_574), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_584), .B(n_593), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g724 ( .A(n_580), .B(n_657), .Y(n_724) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g692 ( .A(n_581), .B(n_652), .Y(n_692) );
AOI32xp33_ASAP7_75t_L g605 ( .A1(n_582), .A2(n_588), .A3(n_606), .B1(n_608), .B2(n_609), .Y(n_605) );
AOI322xp5_ASAP7_75t_L g707 ( .A1(n_582), .A2(n_614), .A3(n_697), .B1(n_708), .B2(n_709), .C1(n_710), .C2(n_712), .Y(n_707) );
INVx2_ASAP7_75t_L g587 ( .A(n_583), .Y(n_587) );
INVx1_ASAP7_75t_L g697 ( .A(n_583), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_585), .B(n_591), .Y(n_640) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_586), .B(n_652), .Y(n_702) );
INVx1_ASAP7_75t_L g589 ( .A(n_587), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_587), .B(n_616), .Y(n_706) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_595), .B(n_690), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B1(n_601), .B2(n_604), .C(n_605), .Y(n_596) );
OR2x2_ASAP7_75t_L g617 ( .A(n_598), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g626 ( .A(n_598), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g651 ( .A(n_599), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g655 ( .A(n_609), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B1(n_617), .B2(n_619), .C(n_620), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_613), .A2(n_644), .B1(n_648), .B2(n_649), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_614), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_614), .Y(n_719) );
INVx1_ASAP7_75t_L g713 ( .A(n_616), .Y(n_713) );
INVx1_ASAP7_75t_SL g648 ( .A(n_617), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_619), .B(n_647), .Y(n_709) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_624), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g690 ( .A(n_624), .Y(n_690) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
OAI221xp5_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_633), .B1(n_635), .B2(n_636), .C(n_638), .Y(n_628) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_630), .A2(n_648), .B1(n_694), .B2(n_695), .Y(n_693) );
CKINVDCx14_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g712 ( .A1(n_635), .A2(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR3xp33_ASAP7_75t_SL g641 ( .A(n_642), .B(n_674), .C(n_698), .Y(n_641) );
NAND4xp25_ASAP7_75t_L g642 ( .A(n_643), .B(n_650), .C(n_658), .D(n_665), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g721 ( .A(n_646), .Y(n_721) );
INVx3_ASAP7_75t_SL g715 ( .A(n_647), .Y(n_715) );
OR2x2_ASAP7_75t_L g720 ( .A(n_647), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_655), .B2(n_657), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_652), .B(n_670), .Y(n_711) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_660), .B(n_662), .Y(n_658) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_677), .B(n_680), .C(n_693), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g708 ( .A(n_679), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B1(n_686), .B2(n_689), .C1(n_691), .C2(n_692), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND4xp25_ASAP7_75t_SL g717 ( .A(n_690), .B(n_718), .C(n_719), .D(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g698 ( .A(n_699), .B(n_707), .C(n_716), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_716) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
endmodule