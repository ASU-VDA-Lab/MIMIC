module fake_jpeg_14583_n_364 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_364);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_364;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_58),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_64),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_14),
.Y(n_62)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_35),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_24),
.B1(n_21),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_34),
.C(n_32),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_99),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_24),
.B1(n_21),
.B2(n_30),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_24),
.B1(n_14),
.B2(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_14),
.B1(n_36),
.B2(n_26),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_36),
.B1(n_18),
.B2(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_82),
.A2(n_89),
.B1(n_97),
.B2(n_87),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_83),
.B(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_18),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_39),
.A2(n_25),
.B1(n_33),
.B2(n_17),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_96),
.B(n_106),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_17),
.B1(n_19),
.B2(n_33),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_34),
.C(n_32),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_34),
.B(n_32),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_0),
.B(n_6),
.Y(n_152)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_48),
.A2(n_23),
.B1(n_19),
.B2(n_31),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_38),
.A2(n_31),
.B1(n_29),
.B2(n_35),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_56),
.A2(n_31),
.B1(n_35),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_31),
.B1(n_1),
.B2(n_3),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_8),
.C(n_1),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_11),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_41),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_153)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_65),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_118),
.B(n_141),
.Y(n_181)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_60),
.B1(n_63),
.B2(n_43),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_12),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_123),
.B(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_131),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_55),
.B1(n_46),
.B2(n_45),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_126),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_69),
.Y(n_127)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_11),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_66),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_139),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_73),
.B(n_10),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_134),
.B(n_150),
.Y(n_195)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_54),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_147),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_163),
.B(n_130),
.Y(n_182)
);

INVx2_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_144),
.A2(n_152),
.B(n_168),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_54),
.B1(n_3),
.B2(n_5),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_153),
.B1(n_155),
.B2(n_72),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_5),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_90),
.B(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_6),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_163),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_72),
.Y(n_154)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_13),
.B1(n_12),
.B2(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_90),
.B(n_12),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_162),
.B(n_86),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g211 ( 
.A(n_158),
.Y(n_211)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_84),
.A2(n_0),
.B1(n_13),
.B2(n_115),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_98),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_78),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_0),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_84),
.A2(n_115),
.B1(n_107),
.B2(n_88),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_109),
.A2(n_107),
.B1(n_88),
.B2(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_126),
.Y(n_196)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_204),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_78),
.C(n_91),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_100),
.B1(n_94),
.B2(n_108),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_174),
.A2(n_179),
.B1(n_191),
.B2(n_192),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_104),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_175),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_108),
.B1(n_135),
.B2(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_176),
.A2(n_188),
.B1(n_203),
.B2(n_206),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_124),
.B1(n_151),
.B2(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_131),
.C(n_125),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_190),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_140),
.A2(n_148),
.B(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_193),
.B(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_167),
.B1(n_149),
.B2(n_129),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_120),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_164),
.B1(n_149),
.B2(n_129),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_127),
.B1(n_154),
.B2(n_122),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_166),
.B(n_133),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_119),
.A2(n_121),
.B1(n_159),
.B2(n_136),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_178),
.B1(n_194),
.B2(n_198),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_185),
.B(n_200),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_122),
.A2(n_127),
.B1(n_154),
.B2(n_138),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_133),
.C(n_138),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_142),
.A2(n_139),
.B1(n_145),
.B2(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_124),
.B(n_130),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_205),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_141),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_139),
.A2(n_145),
.B1(n_118),
.B2(n_144),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_209),
.A2(n_202),
.B1(n_176),
.B2(n_178),
.Y(n_238)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_222),
.Y(n_274)
);

NAND2x1p5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_181),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_216),
.A2(n_219),
.B(n_230),
.Y(n_268)
);

AO21x2_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_196),
.B(n_184),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_217),
.A2(n_240),
.B1(n_242),
.B2(n_247),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_220),
.B(n_238),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_183),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_228),
.B(n_239),
.Y(n_279)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_246),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_208),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_251),
.B(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_180),
.B(n_200),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_175),
.A2(n_209),
.B1(n_206),
.B2(n_184),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_188),
.B(n_182),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_198),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_186),
.A2(n_175),
.B1(n_204),
.B2(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_172),
.B(n_192),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_192),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_189),
.A2(n_176),
.B1(n_130),
.B2(n_178),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_217),
.B1(n_225),
.B2(n_242),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_215),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_236),
.C(n_220),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_257),
.A2(n_258),
.B(n_265),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_248),
.B(n_251),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_217),
.A2(n_250),
.B1(n_234),
.B2(n_219),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_264),
.B1(n_266),
.B2(n_270),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_236),
.C(n_216),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_217),
.B1(n_251),
.B2(n_230),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_216),
.B(n_218),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_234),
.A2(n_238),
.B1(n_221),
.B2(n_244),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_221),
.B(n_223),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_267),
.A2(n_271),
.B(n_272),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_218),
.A2(n_230),
.B1(n_247),
.B2(n_231),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_232),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_222),
.B(n_226),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_229),
.C(n_233),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_252),
.A2(n_242),
.B1(n_217),
.B2(n_176),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_236),
.C(n_139),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_218),
.A2(n_217),
.B1(n_246),
.B2(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_264),
.B(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_290),
.B(n_271),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_253),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_279),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_270),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_254),
.Y(n_298)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_302),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_305),
.B1(n_276),
.B2(n_274),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_257),
.C(n_265),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_267),
.C(n_260),
.Y(n_320)
);

BUFx4f_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_294),
.A2(n_280),
.B1(n_269),
.B2(n_259),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_315),
.B1(n_287),
.B2(n_301),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_269),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_304),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_267),
.B1(n_277),
.B2(n_263),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_297),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_287),
.B1(n_285),
.B2(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_327),
.B1(n_329),
.B2(n_335),
.Y(n_337)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_299),
.B(n_297),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_320),
.C(n_314),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_285),
.B1(n_300),
.B2(n_293),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_300),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_298),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_334),
.B(n_308),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_295),
.B(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_341),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_313),
.B1(n_318),
.B2(n_319),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_342),
.A2(n_345),
.B1(n_305),
.B2(n_327),
.Y(n_346)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_346),
.A2(n_345),
.B1(n_335),
.B2(n_334),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_340),
.A2(n_330),
.B1(n_324),
.B2(n_326),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_348),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_325),
.Y(n_348)
);

NOR2x1_ASAP7_75t_SL g351 ( 
.A(n_349),
.B(n_305),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_352),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_325),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_353),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_358),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_353),
.B(n_354),
.Y(n_358)
);

AOI321xp33_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_318),
.A3(n_319),
.B1(n_350),
.B2(n_324),
.C(n_330),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_289),
.B1(n_332),
.B2(n_331),
.Y(n_361)
);

AO221x1_ASAP7_75t_L g362 ( 
.A1(n_361),
.A2(n_271),
.B1(n_336),
.B2(n_343),
.C(n_344),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_310),
.B(n_290),
.C(n_338),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_337),
.Y(n_364)
);


endmodule