module fake_jpeg_3643_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_17),
.B(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_48),
.B1(n_62),
.B2(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_82),
.B1(n_72),
.B2(n_71),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_48),
.B1(n_62),
.B2(n_60),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_51),
.B1(n_58),
.B2(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_48),
.B1(n_62),
.B2(n_61),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_66),
.B1(n_65),
.B2(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_60),
.B1(n_50),
.B2(n_49),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_68),
.B1(n_6),
.B2(n_8),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_99),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_24),
.B(n_42),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_72),
.C(n_71),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_104),
.B1(n_100),
.B2(n_95),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_1),
.C(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_4),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_23),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_81),
.B1(n_79),
.B2(n_55),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_25),
.C(n_41),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_22),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_144),
.C(n_13),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_10),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_142),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_43),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_12),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_28),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_114),
.B(n_121),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_30),
.C(n_39),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_158),
.C(n_34),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_21),
.C(n_36),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_16),
.B(n_17),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_165),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_141),
.B(n_132),
.C(n_144),
.D(n_134),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_150),
.Y(n_182)
);

OA21x2_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_31),
.B(n_33),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_174),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_35),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_179),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_161),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_156),
.B1(n_148),
.B2(n_153),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_172),
.B1(n_168),
.B2(n_167),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_154),
.C(n_151),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_178),
.B(n_184),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_192),
.B(n_185),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_185),
.B(n_177),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_40),
.C(n_152),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_170),
.Y(n_198)
);


endmodule