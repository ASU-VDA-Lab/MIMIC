module real_aes_8909_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_385;
wire n_275;
wire n_649;
wire n_358;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_691;
wire n_498;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_623;
wire n_249;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_698;
wire n_371;
wire n_541;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_0), .A2(n_209), .B1(n_316), .B2(n_320), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g322 ( .A1(n_1), .A2(n_93), .B1(n_323), .B2(n_329), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_2), .A2(n_219), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_3), .A2(n_216), .B1(n_390), .B2(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_4), .A2(n_226), .B1(n_374), .B2(n_465), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_5), .A2(n_28), .B1(n_664), .B2(n_677), .C(n_678), .Y(n_676) );
AOI22xp5_ASAP7_75t_SL g391 ( .A1(n_6), .A2(n_49), .B1(n_392), .B2(n_394), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_7), .A2(n_148), .B1(n_424), .B2(n_509), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_8), .B(n_415), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_9), .A2(n_236), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_10), .A2(n_108), .B1(n_370), .B2(n_416), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_11), .A2(n_196), .B1(n_335), .B2(n_339), .Y(n_334) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_12), .A2(n_125), .B1(n_295), .B2(n_359), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_13), .A2(n_123), .B1(n_420), .B2(n_564), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_14), .A2(n_198), .B1(n_369), .B2(n_521), .C(n_693), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_15), .A2(n_97), .B1(n_114), .B2(n_468), .C1(n_529), .C2(n_531), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_16), .A2(n_23), .B1(n_362), .B2(n_462), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_17), .A2(n_231), .B1(n_296), .B2(n_462), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_18), .A2(n_156), .B1(n_316), .B2(n_343), .Y(n_667) );
AOI22xp5_ASAP7_75t_SL g388 ( .A1(n_19), .A2(n_232), .B1(n_389), .B2(n_390), .Y(n_388) );
AO22x2_ASAP7_75t_L g262 ( .A1(n_20), .A2(n_70), .B1(n_263), .B2(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g717 ( .A(n_20), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_21), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_22), .A2(n_53), .B1(n_508), .B2(n_509), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_24), .B(n_365), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_25), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_26), .A2(n_140), .B1(n_317), .B2(n_335), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_27), .A2(n_173), .B1(n_654), .B2(n_691), .Y(n_743) );
AOI22xp5_ASAP7_75t_SL g380 ( .A1(n_29), .A2(n_120), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_30), .A2(n_224), .B1(n_423), .B2(n_424), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_31), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_32), .A2(n_199), .B1(n_449), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_33), .A2(n_230), .B1(n_375), .B2(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g758 ( .A(n_34), .Y(n_758) );
AO22x1_ASAP7_75t_L g760 ( .A1(n_34), .A2(n_722), .B1(n_758), .B2(n_761), .Y(n_760) );
AO22x2_ASAP7_75t_L g266 ( .A1(n_35), .A2(n_73), .B1(n_263), .B2(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g718 ( .A(n_35), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_36), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_37), .A2(n_169), .B1(n_347), .B2(n_392), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_38), .A2(n_180), .B1(n_378), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_39), .A2(n_86), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_40), .A2(n_55), .B1(n_412), .B2(n_462), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_41), .A2(n_144), .B1(n_348), .B2(n_517), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_42), .A2(n_142), .B1(n_190), .B2(n_407), .C1(n_614), .C2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_43), .A2(n_238), .B1(n_348), .B2(n_566), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_44), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_45), .A2(n_67), .B1(n_495), .B2(n_496), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_46), .Y(n_456) );
XOR2xp5_ASAP7_75t_L g513 ( .A(n_47), .B(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_48), .A2(n_483), .B1(n_484), .B2(n_511), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_48), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_50), .A2(n_221), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_51), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_52), .A2(n_176), .B1(n_316), .B2(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_54), .A2(n_111), .B1(n_382), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_56), .A2(n_168), .B1(n_317), .B2(n_599), .Y(n_598) );
AOI222xp33_ASAP7_75t_L g697 ( .A1(n_57), .A2(n_77), .B1(n_134), .B2(n_359), .C1(n_408), .C2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_58), .A2(n_131), .B1(n_461), .B2(n_465), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_59), .B(n_370), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_60), .A2(n_102), .B1(n_385), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_61), .A2(n_110), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_62), .A2(n_109), .B1(n_566), .B2(n_684), .C(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_63), .A2(n_217), .B1(n_374), .B2(n_377), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_64), .A2(n_721), .B1(n_748), .B2(n_749), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_64), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_65), .A2(n_71), .B1(n_520), .B2(n_521), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_66), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_68), .A2(n_189), .B1(n_347), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_69), .A2(n_130), .B1(n_329), .B2(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_72), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_74), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_75), .B(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_76), .A2(n_159), .B1(n_421), .B2(n_427), .Y(n_652) );
AND2x2_ASAP7_75t_L g246 ( .A(n_78), .B(n_247), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_79), .Y(n_441) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_80), .A2(n_138), .B1(n_389), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_81), .A2(n_99), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_82), .A2(n_126), .B1(n_361), .B2(n_362), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_83), .A2(n_166), .B1(n_502), .B2(n_564), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_84), .Y(n_642) );
INVx1_ASAP7_75t_L g243 ( .A(n_85), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_87), .A2(n_100), .B1(n_385), .B2(n_451), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_88), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_89), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_90), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_91), .A2(n_106), .B1(n_343), .B2(n_526), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_92), .Y(n_312) );
OA22x2_ASAP7_75t_L g602 ( .A1(n_94), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_94), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_95), .A2(n_127), .B1(n_430), .B2(n_655), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_96), .A2(n_98), .B1(n_329), .B2(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_101), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_103), .A2(n_107), .B1(n_526), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_104), .A2(n_152), .B1(n_359), .B2(n_362), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_105), .A2(n_194), .B1(n_321), .B2(n_325), .Y(n_586) );
XOR2x2_ASAP7_75t_L g632 ( .A(n_112), .B(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_113), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_115), .A2(n_193), .B1(n_343), .B2(n_347), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_116), .Y(n_304) );
XNOR2x2_ASAP7_75t_L g660 ( .A(n_117), .B(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_118), .A2(n_139), .B1(n_394), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_119), .Y(n_357) );
INVx2_ASAP7_75t_L g247 ( .A(n_121), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_122), .A2(n_155), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_124), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_128), .Y(n_736) );
OA22x2_ASAP7_75t_L g537 ( .A1(n_129), .A2(n_538), .B1(n_539), .B2(n_558), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_129), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_132), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_133), .B(n_367), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_135), .B(n_520), .Y(n_572) );
AND2x6_ASAP7_75t_L g242 ( .A(n_136), .B(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_136), .Y(n_711) );
AO22x2_ASAP7_75t_L g272 ( .A1(n_137), .A2(n_201), .B1(n_263), .B2(n_267), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_141), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_143), .A2(n_220), .B1(n_296), .B2(n_462), .Y(n_570) );
AOI22xp5_ASAP7_75t_SL g383 ( .A1(n_145), .A2(n_200), .B1(n_384), .B2(n_385), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_146), .A2(n_210), .B1(n_389), .B2(n_566), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_147), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_149), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_150), .A2(n_188), .B1(n_282), .B2(n_375), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_151), .B(n_369), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_153), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_154), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_157), .A2(n_163), .B1(n_423), .B2(n_453), .Y(n_626) );
AO22x2_ASAP7_75t_L g270 ( .A1(n_158), .A2(n_212), .B1(n_263), .B2(n_264), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_160), .A2(n_235), .B1(n_317), .B2(n_430), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_161), .A2(n_435), .B1(n_473), .B2(n_474), .Y(n_434) );
INVx1_ASAP7_75t_L g473 ( .A(n_161), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_162), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_164), .B(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_165), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_167), .A2(n_181), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_170), .A2(n_191), .B1(n_381), .B2(n_390), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_171), .A2(n_195), .B1(n_394), .B2(n_552), .Y(n_668) );
INVx1_ASAP7_75t_L g396 ( .A(n_172), .Y(n_396) );
AO22x1_ASAP7_75t_L g674 ( .A1(n_174), .A2(n_675), .B1(n_699), .B2(n_700), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_174), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_175), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_177), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_178), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_179), .A2(n_227), .B1(n_329), .B2(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_182), .A2(n_183), .B1(n_394), .B2(n_423), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_184), .A2(n_234), .B1(n_424), .B2(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_185), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_186), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_187), .B(n_367), .Y(n_573) );
OA22x2_ASAP7_75t_L g399 ( .A1(n_192), .A2(n_400), .B1(n_401), .B2(n_431), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_192), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g239 ( .A1(n_197), .A2(n_240), .B(n_248), .C(n_719), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_201), .B(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_202), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_203), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_204), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_205), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_206), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_207), .A2(n_237), .B1(n_337), .B2(n_345), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_208), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_211), .Y(n_590) );
INVx1_ASAP7_75t_L g714 ( .A(n_212), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_213), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_214), .B(n_361), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_215), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_218), .Y(n_273) );
INVx1_ASAP7_75t_L g263 ( .A(n_222), .Y(n_263) );
INVx1_ASAP7_75t_L g265 ( .A(n_222), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_223), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_225), .A2(n_229), .B1(n_430), .B2(n_453), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_228), .B(n_365), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_233), .Y(n_735) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_243), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_244), .A2(n_709), .B(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_534), .B1(n_704), .B2(n_705), .C(n_706), .Y(n_248) );
INVx1_ASAP7_75t_L g705 ( .A(n_249), .Y(n_705) );
AOI22xp5_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_477), .B1(n_478), .B2(n_533), .Y(n_249) );
INVx1_ASAP7_75t_L g533 ( .A(n_250), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B1(n_398), .B2(n_476), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_350), .B1(n_351), .B2(n_397), .Y(n_252) );
INVx2_ASAP7_75t_L g397 ( .A(n_253), .Y(n_397) );
XNOR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_313), .Y(n_255) );
NOR3xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_278), .C(n_300), .Y(n_256) );
OAI22xp5_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_273), .B1(n_274), .B2(n_277), .Y(n_257) );
OAI221xp5_ASAP7_75t_SL g455 ( .A1(n_258), .A2(n_456), .B1(n_457), .B2(n_459), .C(n_460), .Y(n_455) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx3_ASAP7_75t_L g609 ( .A(n_259), .Y(n_609) );
INVx2_ASAP7_75t_L g638 ( .A(n_259), .Y(n_638) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
INVx2_ASAP7_75t_L g338 ( .A(n_260), .Y(n_338) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_266), .Y(n_260) );
AND2x2_ASAP7_75t_L g276 ( .A(n_261), .B(n_266), .Y(n_276) );
AND2x2_ASAP7_75t_L g319 ( .A(n_261), .B(n_285), .Y(n_319) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g286 ( .A(n_262), .B(n_272), .Y(n_286) );
AND2x2_ASAP7_75t_L g290 ( .A(n_262), .B(n_266), .Y(n_290) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g267 ( .A(n_265), .Y(n_267) );
INVx2_ASAP7_75t_L g285 ( .A(n_266), .Y(n_285) );
INVx1_ASAP7_75t_L g331 ( .A(n_266), .Y(n_331) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g349 ( .A(n_269), .B(n_319), .Y(n_349) );
AND2x6_ASAP7_75t_L g367 ( .A(n_269), .B(n_276), .Y(n_367) );
AND2x4_ASAP7_75t_L g372 ( .A(n_269), .B(n_338), .Y(n_372) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g284 ( .A(n_270), .Y(n_284) );
INVx1_ASAP7_75t_L g292 ( .A(n_270), .Y(n_292) );
INVx1_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_270), .B(n_272), .Y(n_332) );
AND2x2_ASAP7_75t_L g291 ( .A(n_271), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g328 ( .A(n_272), .B(n_311), .Y(n_328) );
INVx2_ASAP7_75t_L g458 ( .A(n_274), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_274), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
BUFx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g728 ( .A(n_275), .Y(n_728) );
AND2x4_ASAP7_75t_L g321 ( .A(n_276), .B(n_291), .Y(n_321) );
AND2x2_ASAP7_75t_L g327 ( .A(n_276), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_276), .B(n_328), .Y(n_688) );
OAI222xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_287), .B1(n_288), .B2(n_293), .C1(n_294), .C2(n_299), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_282), .Y(n_361) );
BUFx2_ASAP7_75t_L g407 ( .A(n_282), .Y(n_407) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_282), .Y(n_465) );
BUFx4f_ASAP7_75t_SL g575 ( .A(n_282), .Y(n_575) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g298 ( .A(n_284), .Y(n_298) );
INVx1_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
AND2x4_ASAP7_75t_L g297 ( .A(n_286), .B(n_298), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_286), .B(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g375 ( .A(n_286), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx4_ASAP7_75t_L g356 ( .A(n_289), .Y(n_356) );
INVx2_ASAP7_75t_L g404 ( .A(n_289), .Y(n_404) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_289), .Y(n_468) );
BUFx3_ASAP7_75t_L g614 ( .A(n_289), .Y(n_614) );
INVx2_ASAP7_75t_L g641 ( .A(n_289), .Y(n_641) );
AND2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g308 ( .A(n_290), .Y(n_308) );
AND2x4_ASAP7_75t_L g378 ( .A(n_290), .B(n_310), .Y(n_378) );
AND2x2_ASAP7_75t_L g318 ( .A(n_291), .B(n_319), .Y(n_318) );
AND2x6_ASAP7_75t_L g337 ( .A(n_291), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx4f_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_297), .Y(n_362) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_297), .Y(n_409) );
OAI22xp5_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_304), .B1(n_305), .B2(n_312), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_301), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_301), .A2(n_305), .B1(n_735), .B2(n_736), .Y(n_734) );
BUFx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_302), .A2(n_307), .B1(n_616), .B2(n_617), .Y(n_615) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_302), .Y(n_648) );
AND2x2_ASAP7_75t_L g564 ( .A(n_303), .B(n_341), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_305), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_646) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g696 ( .A(n_306), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_307), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_333), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_322), .Y(n_314) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx3_ASAP7_75t_L g428 ( .A(n_317), .Y(n_428) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_317), .Y(n_508) );
BUFx3_ASAP7_75t_L g740 ( .A(n_317), .Y(n_740) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_SL g381 ( .A(n_318), .Y(n_381) );
INVx2_ASAP7_75t_L g621 ( .A(n_318), .Y(n_621) );
BUFx2_ASAP7_75t_SL g677 ( .A(n_318), .Y(n_677) );
AND2x4_ASAP7_75t_L g340 ( .A(n_319), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g346 ( .A(n_319), .B(n_328), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_319), .B(n_328), .Y(n_440) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx6_ASAP7_75t_L g395 ( .A(n_321), .Y(n_395) );
BUFx3_ASAP7_75t_L g424 ( .A(n_321), .Y(n_424) );
BUFx3_ASAP7_75t_L g453 ( .A(n_321), .Y(n_453) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g384 ( .A(n_325), .Y(n_384) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_325), .Y(n_654) );
INVx4_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g430 ( .A(n_326), .Y(n_430) );
INVx2_ASAP7_75t_L g446 ( .A(n_326), .Y(n_446) );
BUFx3_ASAP7_75t_L g505 ( .A(n_326), .Y(n_505) );
INVx1_ASAP7_75t_L g556 ( .A(n_326), .Y(n_556) );
INVx5_ASAP7_75t_L g623 ( .A(n_326), .Y(n_623) );
INVx8_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx6_ASAP7_75t_SL g386 ( .A(n_330), .Y(n_386) );
INVx1_ASAP7_75t_L g655 ( .A(n_330), .Y(n_655) );
OR2x6_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g376 ( .A(n_331), .Y(n_376) );
INVx1_ASAP7_75t_L g341 ( .A(n_332), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_342), .Y(n_333) );
INVx5_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g449 ( .A(n_336), .Y(n_449) );
INVx4_ASAP7_75t_L g552 ( .A(n_336), .Y(n_552) );
INVx2_ASAP7_75t_SL g578 ( .A(n_336), .Y(n_578) );
INVx11_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx11_ASAP7_75t_L g393 ( .A(n_337), .Y(n_393) );
INVx1_ASAP7_75t_L g442 ( .A(n_339), .Y(n_442) );
BUFx2_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g390 ( .A(n_340), .Y(n_390) );
BUFx2_ASAP7_75t_SL g421 ( .A(n_340), .Y(n_421) );
BUFx3_ASAP7_75t_L g526 ( .A(n_340), .Y(n_526) );
BUFx3_ASAP7_75t_L g566 ( .A(n_340), .Y(n_566) );
BUFx3_ASAP7_75t_L g599 ( .A(n_340), .Y(n_599) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx4f_ASAP7_75t_SL g509 ( .A(n_345), .Y(n_509) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g389 ( .A(n_346), .Y(n_389) );
BUFx3_ASAP7_75t_L g420 ( .A(n_346), .Y(n_420) );
BUFx3_ASAP7_75t_L g525 ( .A(n_346), .Y(n_525) );
BUFx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g382 ( .A(n_349), .Y(n_382) );
BUFx3_ASAP7_75t_L g451 ( .A(n_349), .Y(n_451) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_349), .Y(n_502) );
INVx2_ASAP7_75t_L g742 ( .A(n_349), .Y(n_742) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
XOR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_396), .Y(n_352) );
NAND3x1_ASAP7_75t_L g353 ( .A(n_354), .B(n_379), .C(n_387), .Y(n_353) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_363), .Y(n_354) );
OAI21xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_357), .B(n_358), .Y(n_355) );
BUFx2_ASAP7_75t_L g546 ( .A(n_356), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_356), .A2(n_569), .B(n_570), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_356), .A2(n_590), .B(n_591), .Y(n_589) );
INVx4_ASAP7_75t_L g698 ( .A(n_356), .Y(n_698) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx4_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g530 ( .A(n_362), .Y(n_530) );
BUFx4f_ASAP7_75t_SL g673 ( .A(n_362), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_368), .C(n_373), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g416 ( .A(n_366), .Y(n_416) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g492 ( .A(n_367), .Y(n_492) );
BUFx4f_ASAP7_75t_L g521 ( .A(n_367), .Y(n_521) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx5_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
INVx2_ASAP7_75t_L g520 ( .A(n_371), .Y(n_520) );
INVx4_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
BUFx2_ASAP7_75t_L g461 ( .A(n_375), .Y(n_461) );
BUFx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_378), .Y(n_462) );
BUFx3_ASAP7_75t_L g531 ( .A(n_378), .Y(n_531) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g517 ( .A(n_386), .Y(n_517) );
BUFx4f_ASAP7_75t_SL g691 ( .A(n_386), .Y(n_691) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_391), .Y(n_387) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx4_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
INVx3_ASAP7_75t_L g684 ( .A(n_393), .Y(n_684) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g681 ( .A(n_395), .Y(n_681) );
INVx2_ASAP7_75t_L g746 ( .A(n_395), .Y(n_746) );
INVx1_ASAP7_75t_L g476 ( .A(n_398), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_432), .B1(n_433), .B2(n_475), .Y(n_398) );
INVx1_ASAP7_75t_L g475 ( .A(n_399), .Y(n_475) );
INVx2_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
NAND2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_417), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_410), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g730 ( .A(n_407), .Y(n_730) );
INVx2_ASAP7_75t_L g643 ( .A(n_408), .Y(n_643) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g471 ( .A(n_409), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g495 ( .A(n_413), .Y(n_495) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_425), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_436), .B(n_454), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_447), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_441), .B1(n_442), .B2(n_443), .C(n_444), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_438), .A2(n_679), .B1(n_680), .B2(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_463), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_457), .A2(n_636), .B1(n_637), .B2(n_639), .Y(n_635) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g497 ( .A(n_462), .Y(n_497) );
OAI222xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B1(n_467), .B2(n_469), .C1(n_470), .C2(n_472), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
OAI222xp33_ASAP7_75t_L g729 ( .A1(n_467), .A2(n_643), .B1(n_730), .B2(n_731), .C1(n_732), .C2(n_733), .Y(n_729) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g487 ( .A(n_468), .Y(n_487) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B1(n_512), .B2(n_532), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g511 ( .A(n_484), .Y(n_511) );
NAND3x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_498), .C(n_506), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_486), .B(n_490), .Y(n_485) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_488), .B(n_489), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .C(n_494), .Y(n_490) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g664 ( .A(n_501), .Y(n_664) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_510), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_512), .Y(n_532) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND5xp2_ASAP7_75t_SL g514 ( .A(n_515), .B(n_516), .C(n_518), .D(n_523), .E(n_528), .Y(n_514) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_519), .B(n_522), .Y(n_518) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g704 ( .A(n_534), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_581), .B1(n_702), .B2(n_703), .Y(n_534) );
INVx1_ASAP7_75t_L g702 ( .A(n_535), .Y(n_702) );
OAI22xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_537), .B1(n_559), .B2(n_560), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g558 ( .A(n_539), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
NOR2xp67_ASAP7_75t_SL g540 ( .A(n_541), .B(n_545), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .C(n_544), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
XOR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_580), .Y(n_560) );
NAND3x1_ASAP7_75t_L g561 ( .A(n_562), .B(n_567), .C(n_576), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .C(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g703 ( .A(n_581), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_628), .B1(n_629), .B2(n_701), .Y(n_581) );
CKINVDCx14_ASAP7_75t_R g701 ( .A(n_582), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_601), .B1(n_602), .B2(n_627), .Y(n_582) );
INVx3_ASAP7_75t_L g627 ( .A(n_583), .Y(n_627) );
XOR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_600), .Y(n_583) );
NAND3x1_ASAP7_75t_SL g584 ( .A(n_585), .B(n_588), .C(n_596), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .C(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND3x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_618), .C(n_624), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .C(n_615), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
XOR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_674), .Y(n_629) );
OAI22xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_632), .B1(n_659), .B2(n_660), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_650), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_640), .C(n_646), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_637), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND4xp75_ASAP7_75t_L g661 ( .A(n_662), .B(n_666), .C(n_669), .D(n_672), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AND2x2_ASAP7_75t_SL g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g700 ( .A(n_675), .Y(n_700) );
AND4x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_683), .C(n_692), .D(n_697), .Y(n_675) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_689), .B2(n_690), .Y(n_685) );
BUFx2_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .Y(n_707) );
OR2x2_ASAP7_75t_SL g764 ( .A(n_708), .B(n_713), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_710), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_710), .B(n_754), .Y(n_757) );
CKINVDCx16_ASAP7_75t_R g754 ( .A(n_711), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OAI322xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_750), .A3(n_751), .B1(n_755), .B2(n_758), .C1(n_759), .C2(n_762), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_721), .Y(n_749) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g761 ( .A(n_722), .Y(n_761) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_737), .Y(n_722) );
NOR3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_729), .C(n_734), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_744), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_745), .B(n_747), .Y(n_744) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
endmodule