module fake_netlist_1_8090_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_0), .B(n_6), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_14), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_13), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_18), .B(n_13), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_17), .B1(n_20), .B2(n_19), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_17), .B(n_15), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_21), .B(n_22), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_23), .B(n_11), .Y(n_27) );
OAI33xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_0), .A3(n_1), .B1(n_2), .B2(n_16), .B3(n_4), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_23), .Y(n_29) );
NOR2xp33_ASAP7_75t_L g30 ( .A(n_29), .B(n_24), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_26), .B1(n_25), .B2(n_1), .C(n_2), .Y(n_31) );
AOI21xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_27), .B(n_25), .Y(n_32) );
AOI221xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_28), .B1(n_25), .B2(n_1), .C(n_5), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_32), .Y(n_34) );
INVxp67_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
OAI22xp5_ASAP7_75t_SL g36 ( .A1(n_34), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_36) );
AND2x4_ASAP7_75t_L g37 ( .A(n_35), .B(n_7), .Y(n_37) );
AOI222xp33_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_7), .B1(n_8), .B2(n_9), .C1(n_10), .C2(n_37), .Y(n_38) );
endmodule