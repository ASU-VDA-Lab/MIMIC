module fake_jpeg_20021_n_213 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_26),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_14),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_16),
.B1(n_22),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_16),
.B1(n_22),
.B2(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_31),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_98),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_92),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_29),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_88),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_91),
.B1(n_97),
.B2(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_21),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_13),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_12),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_67),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_6),
.B(n_8),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_111),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_63),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_63),
.B1(n_48),
.B2(n_54),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_122),
.B1(n_92),
.B2(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_84),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_67),
.B1(n_8),
.B2(n_9),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_11),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_12),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_72),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_142),
.B(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_145),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_74),
.C(n_73),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_125),
.C(n_107),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_141),
.B1(n_115),
.B2(n_105),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_80),
.B1(n_70),
.B2(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_74),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_143),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_98),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_121),
.C(n_114),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_69),
.B1(n_88),
.B2(n_82),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_92),
.B(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_144),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_11),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_144),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_152),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_110),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_158),
.C(n_129),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_110),
.B(n_114),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_159),
.B(n_142),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_136),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_116),
.C(n_106),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_138),
.B(n_126),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.C(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_168),
.C(n_175),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_169),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_133),
.B1(n_122),
.B2(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_134),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_130),
.C(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_176),
.B(n_155),
.C(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_130),
.C(n_117),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_113),
.B1(n_146),
.B2(n_117),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_161),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_154),
.C(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_165),
.C(n_176),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_186),
.B(n_166),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_149),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_189),
.C(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_187),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_166),
.B1(n_149),
.B2(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_182),
.B(n_131),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_184),
.B1(n_183),
.B2(n_179),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_178),
.C(n_180),
.Y(n_196)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_194),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_179),
.B1(n_177),
.B2(n_109),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_196),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_189),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_193),
.B1(n_197),
.B2(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_103),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_204),
.B1(n_102),
.B2(n_104),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_102),
.B(n_9),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_209),
.C(n_103),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_119),
.Y(n_213)
);


endmodule