module fake_jpeg_1755_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_5),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_15),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_12),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_33),
.B1(n_21),
.B2(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_26),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_16),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_23),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_33),
.C(n_31),
.Y(n_40)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.C(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_42),
.C(n_32),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_33),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_32),
.B(n_39),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_49),
.B(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_25),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_22),
.C(n_27),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_27),
.B(n_29),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_51),
.B(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_27),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_48),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_25),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_11),
.A3(n_15),
.B1(n_9),
.B2(n_7),
.C1(n_3),
.C2(n_6),
.Y(n_56)
);

AOI31xp33_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_7),
.A3(n_10),
.B(n_14),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_24),
.B(n_10),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.C(n_14),
.Y(n_60)
);


endmodule