module real_jpeg_13177_n_12 (n_5, n_4, n_8, n_0, n_310, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_310;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_3),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_3),
.A2(n_37),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_37),
.B1(n_148),
.B2(n_160),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_7),
.A2(n_43),
.B1(n_46),
.B2(n_152),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_7),
.A2(n_100),
.B1(n_101),
.B2(n_152),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_7),
.A2(n_148),
.B1(n_152),
.B2(n_160),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_9),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_9),
.A2(n_45),
.B1(n_148),
.B2(n_160),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_10),
.B(n_29),
.C(n_48),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_30),
.B1(n_43),
.B2(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_10),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_10),
.B(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_30),
.B1(n_100),
.B2(n_101),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_10),
.A2(n_57),
.B(n_101),
.C(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_30),
.B1(n_148),
.B2(n_160),
.Y(n_165)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_302),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_294),
.B(n_301),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_256),
.B(n_291),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_237),
.B(n_255),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_216),
.B(n_236),
.Y(n_16)
);

AOI321xp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_176),
.A3(n_209),
.B1(n_214),
.B2(n_215),
.C(n_310),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_139),
.B(n_175),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_116),
.B(n_138),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_93),
.B(n_115),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_71),
.B(n_92),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_25),
.B(n_89),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_35),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_27),
.A2(n_32),
.B(n_35),
.Y(n_111)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_75),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_30),
.A2(n_46),
.B(n_58),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_30),
.B(n_101),
.C(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_32),
.A2(n_89),
.B(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_34),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_35),
.A2(n_151),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_41),
.B(n_68),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_41),
.A2(n_173),
.B(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_42),
.B(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_51),
.Y(n_173)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_59),
.C(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_55),
.B(n_106),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_55),
.A2(n_103),
.B(n_106),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_55),
.A2(n_169),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_56),
.B(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_70),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_85),
.B(n_91),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_79),
.B(n_84),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_107),
.C(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_101),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_102),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_104),
.B(n_133),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_104),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_108),
.A2(n_174),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_108),
.B(n_120),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_110),
.A2(n_111),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_110),
.A2(n_111),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_111),
.B(n_233),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_111),
.A2(n_244),
.B(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_137),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_137),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_124),
.B1(n_125),
.B2(n_136),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_125),
.B(n_144),
.C(n_154),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_127),
.CI(n_131),
.CON(n_125),
.SN(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_128),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_130),
.B1(n_148),
.B2(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_132),
.B(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_132),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_141),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_154),
.B2(n_155),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_153),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_166),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_168),
.C(n_171),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_163),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_162),
.A2(n_165),
.B(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_162),
.A2(n_180),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_181),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_169),
.B(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_171),
.A2(n_172),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_171),
.A2(n_172),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_172),
.B(n_264),
.C(n_269),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_172),
.B(n_288),
.C(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_203),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_203),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_187),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_188),
.C(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_186),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_184),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_199),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_196),
.C(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_195),
.A2(n_248),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_195),
.B(n_226),
.Y(n_304)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_196),
.A2(n_198),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_196),
.B(n_299),
.C(n_300),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_201),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_205),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_213),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_235),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_231),
.B2(n_232),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_232),
.C(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.C(n_229),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_239),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_242),
.C(n_250),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_249),
.B2(n_250),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_262),
.B1(n_263),
.B2(n_273),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_260),
.C(n_262),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_274),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_265),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_277),
.C(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_269),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_276),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_285),
.B1(n_286),
.B2(n_290),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_296),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_304),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);


endmodule