module fake_aes_6853_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_30;
wire n_26;
wire n_13;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_10), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_4), .B(n_7), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_6), .A2(n_9), .B1(n_7), .B2(n_5), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
AOI21xp33_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B(n_1), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_17), .B(n_11), .Y(n_19) );
OAI21xp33_ASAP7_75t_L g20 ( .A1(n_14), .A2(n_0), .B(n_2), .Y(n_20) );
INVxp67_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
AOI33xp33_ASAP7_75t_L g22 ( .A1(n_13), .A2(n_0), .A3(n_2), .B1(n_3), .B2(n_4), .B3(n_5), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_19), .B(n_15), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
AO31x2_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_15), .A3(n_13), .B(n_5), .Y(n_25) );
NOR2xp33_ASAP7_75t_SL g26 ( .A(n_23), .B(n_20), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
OR2x6_ASAP7_75t_L g28 ( .A(n_25), .B(n_20), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_18), .B(n_12), .Y(n_30) );
OAI22xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_26), .B1(n_12), .B2(n_16), .Y(n_31) );
NAND3xp33_ASAP7_75t_SL g32 ( .A(n_29), .B(n_25), .C(n_18), .Y(n_32) );
OAI22xp5_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_28), .B1(n_4), .B2(n_6), .Y(n_33) );
CKINVDCx16_ASAP7_75t_R g34 ( .A(n_32), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_32), .Y(n_35) );
OAI22xp5_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_28), .B1(n_3), .B2(n_10), .Y(n_36) );
AOI22xp33_ASAP7_75t_SL g37 ( .A1(n_36), .A2(n_34), .B1(n_35), .B2(n_28), .Y(n_37) );
endmodule