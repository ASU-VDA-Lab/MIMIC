module real_jpeg_21595_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_0),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_0),
.A2(n_26),
.B1(n_32),
.B2(n_50),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_1),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_133),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_133),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_133),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_3),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_126),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_126),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_4),
.B(n_28),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_4),
.A2(n_14),
.B(n_63),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_131),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_4),
.A2(n_105),
.B1(n_110),
.B2(n_190),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_87),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_30),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_4),
.A2(n_30),
.B(n_217),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_257)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_7),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_8),
.B(n_62),
.Y(n_106)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_8),
.B(n_209),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_128),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_128),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_45),
.B(n_60),
.C(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_14),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_319),
.Y(n_325)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_23),
.A2(n_36),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_23),
.A2(n_36),
.B1(n_144),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_23),
.A2(n_265),
.B(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_23),
.A2(n_84),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_24),
.A2(n_28),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_25),
.B(n_30),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_26),
.B(n_131),
.CON(n_130),
.SN(n_130)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_29),
.B1(n_130),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_28),
.B(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_29),
.A2(n_44),
.A3(n_45),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_42),
.B(n_43),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_43),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_31),
.A2(n_36),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_51),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_41),
.A2(n_52),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_49),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_42),
.A2(n_53),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_42),
.A2(n_53),
.B1(n_163),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_42),
.A2(n_51),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_42),
.A2(n_53),
.B1(n_76),
.B2(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g218 ( 
.A(n_43),
.B(n_46),
.Y(n_218)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_46),
.A2(n_64),
.B(n_131),
.C(n_181),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_52),
.A2(n_87),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_52),
.A2(n_77),
.B(n_88),
.Y(n_267)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_68),
.C(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_58),
.A2(n_67),
.B1(n_74),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_65),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_59),
.A2(n_65),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_59),
.A2(n_61),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_59),
.A2(n_61),
.B1(n_185),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_59),
.A2(n_61),
.B1(n_206),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_59),
.A2(n_224),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_59),
.A2(n_61),
.B1(n_113),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_59),
.A2(n_121),
.B(n_257),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_61),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_61),
.B(n_131),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_62),
.B(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_66),
.B(n_122),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_70),
.C(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_70),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_70),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_73),
.B(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_74),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_316),
.A3(n_326),
.B1(n_329),
.B2(n_330),
.C(n_333),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_296),
.B(n_315),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_272),
.B(n_295),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_165),
.B(n_248),
.C(n_271),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_149),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_99),
.B(n_149),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_134),
.B2(n_148),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_118),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_102),
.B(n_118),
.C(n_148),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_112),
.B2(n_117),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_103),
.B(n_117),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_105),
.A2(n_174),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_105),
.A2(n_177),
.B(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_105),
.A2(n_191),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_106),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_106),
.A2(n_109),
.B(n_209),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_139),
.B(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_110),
.B(n_131),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_114),
.B(n_239),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_129),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_135),
.B(n_141),
.C(n_146),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_158),
.B(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_161),
.B(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_247),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_242),
.B(n_246),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_229),
.B(n_241),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_211),
.B(n_228),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_198),
.B(n_210),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_186),
.B(n_197),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_182),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_192),
.B(n_196),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_200),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_209),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_213),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_219),
.B1(n_226),
.B2(n_227),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_238),
.C(n_240),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_269),
.B2(n_270),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_258),
.B2(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_259),
.C(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_268),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_267),
.C(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_294),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_287),
.B2(n_288),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_288),
.C(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_282),
.C(n_286),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_282),
.B1(n_283),
.B2(n_286),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_280),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_285),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_290),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_306),
.B(n_310),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_298),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_313),
.B2(n_314),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_305),
.C(n_314),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_318),
.C(n_323),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_304),
.B(n_318),
.CI(n_323),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_328),
.Y(n_331)
);


endmodule