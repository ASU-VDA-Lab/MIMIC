module fake_jpeg_23996_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_SL g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_39),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_1),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_3),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_26),
.B1(n_25),
.B2(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_50),
.B1(n_62),
.B2(n_13),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_23),
.B1(n_21),
.B2(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_5),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_30),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_61),
.B1(n_42),
.B2(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_49),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_24),
.B(n_18),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_35),
.B(n_11),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_18),
.B1(n_15),
.B2(n_10),
.Y(n_62)
);

XNOR2x1_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_31),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_35),
.B1(n_9),
.B2(n_11),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_67),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_59),
.B(n_48),
.C(n_53),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_55),
.B1(n_51),
.B2(n_60),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_61),
.B1(n_42),
.B2(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_9),
.B(n_12),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_81),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_13),
.B1(n_61),
.B2(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_80),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_88),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_95),
.B1(n_64),
.B2(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_52),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_68),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_68),
.CON(n_100),
.SN(n_100)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_101),
.B(n_92),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_77),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.C(n_106),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_68),
.B(n_66),
.C(n_76),
.D(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_111),
.B(n_94),
.Y(n_119)
);

BUFx12f_ASAP7_75t_SL g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_90),
.C(n_96),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_110),
.B(n_108),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_84),
.C(n_95),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_84),
.B(n_96),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_114),
.B1(n_91),
.B2(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_103),
.B1(n_106),
.B2(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_124),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_126),
.B2(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_126),
.Y(n_132)
);


endmodule