module real_aes_7002_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_358;
wire n_214;
wire n_275;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g472 ( .A1(n_0), .A2(n_155), .B(n_473), .C(n_476), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_1), .B(n_467), .Y(n_478) );
INVx1_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
INVx1_ASAP7_75t_L g193 ( .A(n_3), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_4), .B(n_156), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_5), .A2(n_134), .B1(n_135), .B2(n_441), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_5), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_5), .A2(n_97), .B1(n_441), .B2(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_6), .A2(n_452), .B(n_499), .Y(n_498) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_7), .A2(n_162), .B(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_8), .A2(n_38), .B1(n_159), .B2(n_211), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_9), .B(n_162), .Y(n_179) );
AND2x6_ASAP7_75t_L g164 ( .A(n_10), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_11), .A2(n_164), .B(n_455), .C(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_12), .B(n_39), .Y(n_118) );
INVx1_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
INVx1_ASAP7_75t_L g185 ( .A(n_14), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_15), .B(n_152), .Y(n_205) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_16), .A2(n_41), .B1(n_527), .B2(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_16), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_17), .B(n_156), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_18), .B(n_142), .Y(n_141) );
AO32x2_ASAP7_75t_L g222 ( .A1(n_19), .A2(n_162), .A3(n_163), .B1(n_182), .B2(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_20), .B(n_159), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_21), .B(n_142), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_22), .A2(n_54), .B1(n_159), .B2(n_211), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g219 ( .A1(n_23), .A2(n_82), .B1(n_152), .B2(n_159), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_24), .B(n_159), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_25), .A2(n_163), .B(n_455), .C(n_457), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_26), .A2(n_163), .B(n_455), .C(n_533), .Y(n_532) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_28), .A2(n_98), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_28), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_29), .B(n_201), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_30), .A2(n_452), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_31), .B(n_201), .Y(n_238) );
INVx2_ASAP7_75t_L g154 ( .A(n_32), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_33), .A2(n_487), .B(n_488), .C(n_492), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_34), .B(n_159), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_35), .B(n_201), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_36), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_36), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_37), .B(n_207), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_40), .B(n_451), .Y(n_450) );
AOI222xp33_ASAP7_75t_SL g104 ( .A1(n_41), .A2(n_105), .B1(n_119), .B2(n_735), .C1(n_740), .C2(n_757), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_41), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_42), .B(n_156), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_43), .B(n_452), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_44), .A2(n_487), .B(n_492), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_45), .B(n_159), .Y(n_172) );
INVx1_ASAP7_75t_L g474 ( .A(n_46), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_47), .A2(n_748), .B1(n_749), .B2(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g751 ( .A(n_47), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_48), .A2(n_91), .B1(n_211), .B2(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g513 ( .A(n_49), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_50), .B(n_159), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_51), .B(n_159), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_52), .B(n_452), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_53), .B(n_177), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g158 ( .A1(n_55), .A2(n_60), .B1(n_152), .B2(n_159), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_56), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_56), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_57), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_58), .B(n_159), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_59), .B(n_159), .Y(n_258) );
INVx1_ASAP7_75t_L g165 ( .A(n_61), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_62), .B(n_452), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_63), .B(n_467), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_64), .A2(n_177), .B(n_188), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_65), .B(n_159), .Y(n_194) );
INVx1_ASAP7_75t_L g145 ( .A(n_66), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_67), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_68), .B(n_156), .Y(n_490) );
AO32x2_ASAP7_75t_L g215 ( .A1(n_69), .A2(n_162), .A3(n_163), .B1(n_216), .B2(n_220), .Y(n_215) );
AOI222xp33_ASAP7_75t_SL g120 ( .A1(n_70), .A2(n_121), .B1(n_122), .B2(n_131), .C1(n_726), .C2(n_732), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_71), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_72), .B(n_157), .Y(n_524) );
INVx1_ASAP7_75t_L g257 ( .A(n_73), .Y(n_257) );
INVx1_ASAP7_75t_L g233 ( .A(n_74), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_75), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_76), .B(n_459), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_77), .A2(n_455), .B(n_492), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_78), .B(n_152), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_79), .Y(n_500) );
INVx1_ASAP7_75t_L g110 ( .A(n_80), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_81), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_83), .B(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_84), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_85), .B(n_152), .Y(n_237) );
INVx2_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_87), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_88), .B(n_149), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_89), .B(n_152), .Y(n_173) );
OR2x2_ASAP7_75t_L g114 ( .A(n_90), .B(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g442 ( .A(n_90), .B(n_116), .Y(n_442) );
INVx2_ASAP7_75t_L g725 ( .A(n_90), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_92), .A2(n_103), .B1(n_152), .B2(n_153), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_93), .B(n_452), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_94), .Y(n_489) );
INVxp67_ASAP7_75t_L g503 ( .A(n_95), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_96), .B(n_152), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_97), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_98), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_99), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g520 ( .A(n_100), .Y(n_520) );
INVx1_ASAP7_75t_L g549 ( .A(n_101), .Y(n_549) );
AND2x2_ASAP7_75t_L g515 ( .A(n_102), .B(n_201), .Y(n_515) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_112), .Y(n_107) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g739 ( .A(n_109), .Y(n_739) );
INVx1_ASAP7_75t_L g738 ( .A(n_111), .Y(n_738) );
OA21x2_ASAP7_75t_L g758 ( .A1(n_111), .A2(n_739), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_114), .Y(n_752) );
INVx1_ASAP7_75t_SL g755 ( .A(n_114), .Y(n_755) );
BUFx2_ASAP7_75t_L g759 ( .A(n_114), .Y(n_759) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_115), .B(n_725), .Y(n_734) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g724 ( .A(n_116), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g129 ( .A(n_126), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_442), .B1(n_443), .B2(n_724), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_133), .A2(n_727), .B1(n_729), .B2(n_730), .Y(n_726) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
XNOR2xp5_ASAP7_75t_L g744 ( .A(n_135), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_375), .Y(n_135) );
NOR5xp2_ASAP7_75t_L g136 ( .A(n_137), .B(n_288), .C(n_334), .D(n_347), .E(n_359), .Y(n_136) );
OAI211xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_196), .B(n_242), .C(n_269), .Y(n_137) );
INVx1_ASAP7_75t_SL g370 ( .A(n_138), .Y(n_370) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_166), .Y(n_138) );
AND2x2_ASAP7_75t_L g294 ( .A(n_139), .B(n_167), .Y(n_294) );
AND2x2_ASAP7_75t_L g322 ( .A(n_139), .B(n_268), .Y(n_322) );
AND2x2_ASAP7_75t_L g330 ( .A(n_139), .B(n_273), .Y(n_330) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g260 ( .A(n_140), .B(n_168), .Y(n_260) );
INVx2_ASAP7_75t_L g272 ( .A(n_140), .Y(n_272) );
AND2x2_ASAP7_75t_L g397 ( .A(n_140), .B(n_339), .Y(n_397) );
OR2x2_ASAP7_75t_L g399 ( .A(n_140), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_147), .Y(n_140) );
INVx1_ASAP7_75t_L g266 ( .A(n_141), .Y(n_266) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx1_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_143), .B(n_144), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
NAND3xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_161), .C(n_163), .Y(n_147) );
AO21x1_ASAP7_75t_L g265 ( .A1(n_148), .A2(n_161), .B(n_266), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B1(n_155), .B2(n_158), .Y(n_148) );
INVx2_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
OAI22xp5_ASAP7_75t_SL g216 ( .A1(n_149), .A2(n_157), .B1(n_217), .B2(n_219), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_149), .A2(n_155), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g475 ( .A(n_149), .Y(n_475) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
INVx1_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
AND2x2_ASAP7_75t_L g453 ( .A(n_150), .B(n_178), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_150), .Y(n_456) );
INVx2_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
INVx1_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_175), .B(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_156), .A2(n_172), .B(n_173), .Y(n_171) );
O2A1O1Ixp5_ASAP7_75t_SL g231 ( .A1(n_156), .A2(n_232), .B(n_233), .C(n_234), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_156), .A2(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_156), .B(n_503), .Y(n_502) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g232 ( .A(n_159), .Y(n_232) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_159), .Y(n_551) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
BUFx3_ASAP7_75t_L g218 ( .A(n_160), .Y(n_218) );
AND2x6_ASAP7_75t_L g455 ( .A(n_160), .B(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g467 ( .A(n_161), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_161), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_161), .A2(n_519), .B(n_526), .Y(n_518) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_161), .A2(n_546), .B(n_553), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_161), .B(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_162), .A2(n_170), .B(n_179), .Y(n_169) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_162), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_162), .A2(n_531), .B(n_532), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_163), .A2(n_253), .B(n_256), .Y(n_252) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_164), .A2(n_171), .B(n_174), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_164), .A2(n_184), .B(n_191), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_164), .A2(n_203), .B(n_208), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_164), .A2(n_231), .B(n_235), .Y(n_230) );
AND2x4_ASAP7_75t_L g452 ( .A(n_164), .B(n_453), .Y(n_452) );
INVx4_ASAP7_75t_SL g477 ( .A(n_164), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_164), .B(n_453), .Y(n_521) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g310 ( .A(n_167), .B(n_282), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_167), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g424 ( .A(n_167), .B(n_264), .Y(n_424) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
AND2x2_ASAP7_75t_L g267 ( .A(n_168), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g314 ( .A(n_168), .Y(n_314) );
AND2x2_ASAP7_75t_L g339 ( .A(n_168), .B(n_251), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_168), .B(n_372), .Y(n_409) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g273 ( .A(n_169), .B(n_251), .Y(n_273) );
AND2x2_ASAP7_75t_L g287 ( .A(n_169), .B(n_250), .Y(n_287) );
AND2x2_ASAP7_75t_L g304 ( .A(n_169), .B(n_180), .Y(n_304) );
AND2x2_ASAP7_75t_L g361 ( .A(n_169), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_169), .B(n_268), .Y(n_374) );
AND2x2_ASAP7_75t_L g426 ( .A(n_169), .B(n_351), .Y(n_426) );
INVx2_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g249 ( .A(n_180), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_180), .B(n_251), .Y(n_345) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B(n_195), .Y(n_180) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_181), .A2(n_252), .B(n_259), .Y(n_251) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_182), .B(n_527), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_188), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_186), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_186), .A2(n_534), .B(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_188), .A2(n_549), .B(n_550), .C(n_551), .Y(n_548) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_189), .A2(n_236), .B(n_237), .Y(n_235) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g459 ( .A(n_190), .Y(n_459) );
O2A1O1Ixp5_ASAP7_75t_L g256 ( .A1(n_192), .A2(n_212), .B(n_257), .C(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_192), .A2(n_458), .B(n_460), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_226), .B(n_239), .Y(n_196) );
INVx1_ASAP7_75t_SL g358 ( .A(n_197), .Y(n_358) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_214), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_199), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g241 ( .A(n_200), .Y(n_241) );
INVx1_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
AND2x2_ASAP7_75t_L g299 ( .A(n_200), .B(n_221), .Y(n_299) );
AND2x2_ASAP7_75t_L g333 ( .A(n_200), .B(n_222), .Y(n_333) );
OR2x2_ASAP7_75t_L g352 ( .A(n_200), .B(n_228), .Y(n_352) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_200), .Y(n_366) );
AND2x2_ASAP7_75t_L g379 ( .A(n_200), .B(n_380), .Y(n_379) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_213), .Y(n_200) );
INVx2_ASAP7_75t_L g220 ( .A(n_201), .Y(n_220) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_201), .A2(n_230), .B(n_238), .Y(n_229) );
INVx1_ASAP7_75t_L g465 ( .A(n_201), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_201), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_201), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_203) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_212), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_214), .A2(n_301), .B1(n_302), .B2(n_311), .Y(n_300) );
AND2x2_ASAP7_75t_L g384 ( .A(n_214), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .Y(n_214) );
INVx1_ASAP7_75t_L g245 ( .A(n_215), .Y(n_245) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_215), .Y(n_282) );
INVx1_ASAP7_75t_L g293 ( .A(n_215), .Y(n_293) );
AND2x2_ASAP7_75t_L g308 ( .A(n_215), .B(n_222), .Y(n_308) );
INVx2_ASAP7_75t_L g476 ( .A(n_218), .Y(n_476) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_218), .Y(n_491) );
INVx1_ASAP7_75t_L g462 ( .A(n_220), .Y(n_462) );
OR2x2_ASAP7_75t_L g262 ( .A(n_221), .B(n_247), .Y(n_262) );
AND2x2_ASAP7_75t_L g292 ( .A(n_221), .B(n_293), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_221), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g240 ( .A(n_222), .B(n_241), .Y(n_240) );
BUFx2_ASAP7_75t_L g349 ( .A(n_222), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_226), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g327 ( .A(n_227), .B(n_293), .Y(n_327) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g239 ( .A(n_228), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g298 ( .A(n_228), .Y(n_298) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g247 ( .A(n_229), .Y(n_247) );
OR2x2_ASAP7_75t_L g277 ( .A(n_229), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_229), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g369 ( .A1(n_239), .A2(n_299), .A3(n_370), .B1(n_371), .B2(n_373), .Y(n_369) );
AND2x2_ASAP7_75t_L g295 ( .A(n_240), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_240), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_240), .B(n_327), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_240), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B1(n_261), .B2(n_263), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
AND2x2_ASAP7_75t_L g348 ( .A(n_244), .B(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_245), .B(n_247), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_246), .A2(n_270), .B1(n_274), .B2(n_284), .Y(n_269) );
AND2x2_ASAP7_75t_L g291 ( .A(n_246), .B(n_292), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_246), .A2(n_260), .B(n_308), .C(n_343), .Y(n_342) );
OAI332xp33_ASAP7_75t_L g347 ( .A1(n_246), .A2(n_348), .A3(n_350), .B1(n_352), .B2(n_353), .B3(n_355), .C1(n_356), .C2(n_358), .Y(n_347) );
INVx2_ASAP7_75t_L g388 ( .A(n_246), .Y(n_388) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_247), .Y(n_306) );
INVx1_ASAP7_75t_L g381 ( .A(n_247), .Y(n_381) );
AND2x2_ASAP7_75t_L g435 ( .A(n_247), .B(n_299), .Y(n_435) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_260), .Y(n_248) );
AND2x2_ASAP7_75t_L g315 ( .A(n_250), .B(n_265), .Y(n_315) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g363 ( .A(n_251), .B(n_265), .Y(n_363) );
INVx1_ASAP7_75t_L g372 ( .A(n_251), .Y(n_372) );
INVx1_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g430 ( .A(n_262), .B(n_282), .Y(n_430) );
INVx1_ASAP7_75t_SL g341 ( .A(n_263), .Y(n_341) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
AND2x2_ASAP7_75t_L g368 ( .A(n_264), .B(n_326), .Y(n_368) );
INVx1_ASAP7_75t_L g387 ( .A(n_264), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_264), .B(n_354), .Y(n_389) );
INVx1_ASAP7_75t_L g286 ( .A(n_265), .Y(n_286) );
AND2x2_ASAP7_75t_L g290 ( .A(n_267), .B(n_271), .Y(n_290) );
AND2x2_ASAP7_75t_L g357 ( .A(n_267), .B(n_315), .Y(n_357) );
INVx2_ASAP7_75t_L g400 ( .A(n_267), .Y(n_400) );
INVx2_ASAP7_75t_L g283 ( .A(n_268), .Y(n_283) );
AND2x2_ASAP7_75t_L g285 ( .A(n_268), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g301 ( .A(n_271), .Y(n_301) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_272), .B(n_345), .Y(n_351) );
OR2x2_ASAP7_75t_L g415 ( .A(n_272), .B(n_374), .Y(n_415) );
INVx1_ASAP7_75t_L g439 ( .A(n_272), .Y(n_439) );
INVx1_ASAP7_75t_L g395 ( .A(n_273), .Y(n_395) );
AND2x2_ASAP7_75t_L g440 ( .A(n_273), .B(n_283), .Y(n_440) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_277), .A2(n_303), .B1(n_305), .B2(n_309), .Y(n_302) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI322xp33_ASAP7_75t_SL g386 ( .A1(n_280), .A2(n_387), .A3(n_388), .B1(n_389), .B2(n_390), .C1(n_393), .C2(n_395), .Y(n_386) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
AND2x2_ASAP7_75t_L g383 ( .A(n_281), .B(n_299), .Y(n_383) );
OR2x2_ASAP7_75t_L g417 ( .A(n_281), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g420 ( .A(n_281), .B(n_352), .Y(n_420) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g365 ( .A(n_282), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g421 ( .A(n_282), .B(n_352), .Y(n_421) );
INVx3_ASAP7_75t_L g354 ( .A(n_283), .Y(n_354) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g410 ( .A(n_285), .Y(n_410) );
AOI222xp33_ASAP7_75t_L g289 ( .A1(n_287), .A2(n_290), .B1(n_291), .B2(n_294), .C1(n_295), .C2(n_297), .Y(n_289) );
INVx1_ASAP7_75t_L g320 ( .A(n_287), .Y(n_320) );
NAND3xp33_ASAP7_75t_SL g288 ( .A(n_289), .B(n_300), .C(n_317), .Y(n_288) );
AND2x2_ASAP7_75t_L g405 ( .A(n_292), .B(n_306), .Y(n_405) );
BUFx2_ASAP7_75t_L g296 ( .A(n_293), .Y(n_296) );
INVx1_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_294), .A2(n_330), .B1(n_383), .B2(n_384), .C(n_386), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_296), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
AND2x2_ASAP7_75t_L g336 ( .A(n_299), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_304), .B(n_315), .Y(n_316) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OAI21xp33_ASAP7_75t_L g311 ( .A1(n_306), .A2(n_312), .B(n_316), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_306), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g403 ( .A(n_308), .B(n_385), .Y(n_403) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g326 ( .A(n_314), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_315), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g432 ( .A(n_315), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_323), .B1(n_324), .B2(n_327), .C(n_328), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_319), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g428 ( .A(n_327), .B(n_333), .Y(n_428) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
OAI31xp33_ASAP7_75t_SL g396 ( .A1(n_331), .A2(n_370), .A3(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g385 ( .A(n_332), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_333), .B(n_337), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_338), .B1(n_340), .B2(n_341), .C(n_342), .Y(n_334) );
INVx1_ASAP7_75t_L g340 ( .A(n_336), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_339), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g355 ( .A(n_348), .Y(n_355) );
INVx2_ASAP7_75t_L g391 ( .A(n_349), .Y(n_391) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g377 ( .A(n_354), .B(n_363), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_354), .A2(n_371), .B(n_428), .C(n_429), .Y(n_427) );
OAI221xp5_ASAP7_75t_SL g359 ( .A1(n_355), .A2(n_360), .B1(n_364), .B2(n_367), .C(n_369), .Y(n_359) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_358), .A2(n_423), .B(n_425), .C(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_361), .A2(n_412), .B1(n_414), .B2(n_416), .C(n_419), .Y(n_411) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_401), .C(n_422), .D(n_433), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_378), .B(n_382), .C(n_396), .Y(n_376) );
INVx1_ASAP7_75t_SL g431 ( .A(n_383), .Y(n_431) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g394 ( .A(n_392), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_399), .A2(n_408), .B1(n_420), .B2(n_421), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_406), .C(n_411), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI31xp33_ASAP7_75t_L g433 ( .A1(n_404), .A2(n_434), .A3(n_436), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g728 ( .A(n_442), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_443), .Y(n_729) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_660), .Y(n_443) );
NOR5xp2_ASAP7_75t_L g444 ( .A(n_445), .B(n_591), .C(n_620), .D(n_640), .E(n_647), .Y(n_444) );
OAI211xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_479), .B(n_536), .C(n_578), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_447), .A2(n_663), .B1(n_665), .B2(n_666), .Y(n_662) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_466), .Y(n_447) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_448), .Y(n_539) );
AND2x4_ASAP7_75t_L g571 ( .A(n_448), .B(n_572), .Y(n_571) );
INVx5_ASAP7_75t_L g589 ( .A(n_448), .Y(n_589) );
AND2x2_ASAP7_75t_L g598 ( .A(n_448), .B(n_590), .Y(n_598) );
AND2x2_ASAP7_75t_L g610 ( .A(n_448), .B(n_483), .Y(n_610) );
AND2x2_ASAP7_75t_L g706 ( .A(n_448), .B(n_574), .Y(n_706) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_463), .Y(n_448) );
AOI21xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_454), .B(n_462), .Y(n_449) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx5_ASAP7_75t_L g471 ( .A(n_455), .Y(n_471) );
INVx2_ASAP7_75t_L g461 ( .A(n_459), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_461), .A2(n_489), .B(n_490), .C(n_491), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_461), .A2(n_491), .B(n_513), .C(n_514), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_L g572 ( .A(n_466), .Y(n_572) );
AND2x2_ASAP7_75t_L g590 ( .A(n_466), .B(n_545), .Y(n_590) );
AND2x2_ASAP7_75t_L g609 ( .A(n_466), .B(n_544), .Y(n_609) );
AND2x2_ASAP7_75t_L g649 ( .A(n_466), .B(n_589), .Y(n_649) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_478), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_471), .B(n_472), .C(n_477), .Y(n_469) );
INVx2_ASAP7_75t_L g487 ( .A(n_471), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_471), .A2(n_477), .B(n_500), .C(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g492 ( .A(n_477), .Y(n_492) );
INVxp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_505), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI322xp5_ASAP7_75t_L g708 ( .A1(n_482), .A2(n_516), .A3(n_563), .B1(n_571), .B2(n_625), .C1(n_709), .C2(n_712), .Y(n_708) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
INVx5_ASAP7_75t_L g541 ( .A(n_483), .Y(n_541) );
AND2x2_ASAP7_75t_L g557 ( .A(n_483), .B(n_543), .Y(n_557) );
BUFx2_ASAP7_75t_L g635 ( .A(n_483), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_483), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g712 ( .A(n_483), .B(n_619), .Y(n_712) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_495), .B(n_507), .Y(n_566) );
INVx1_ASAP7_75t_L g593 ( .A(n_495), .Y(n_593) );
AND2x2_ASAP7_75t_L g606 ( .A(n_495), .B(n_528), .Y(n_606) );
AND2x2_ASAP7_75t_L g707 ( .A(n_495), .B(n_625), .Y(n_707) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g561 ( .A(n_496), .B(n_507), .Y(n_561) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_496), .Y(n_569) );
OR2x2_ASAP7_75t_L g576 ( .A(n_496), .B(n_528), .Y(n_576) );
AND2x2_ASAP7_75t_L g586 ( .A(n_496), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_496), .B(n_518), .Y(n_615) );
INVxp67_ASAP7_75t_L g639 ( .A(n_496), .Y(n_639) );
AND2x2_ASAP7_75t_L g646 ( .A(n_496), .B(n_516), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_496), .B(n_528), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_496), .B(n_517), .Y(n_672) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_504), .Y(n_496) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_507), .B(n_529), .Y(n_616) );
OR2x2_ASAP7_75t_L g638 ( .A(n_507), .B(n_517), .Y(n_638) );
AND2x2_ASAP7_75t_L g651 ( .A(n_507), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_507), .B(n_606), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_507), .A2(n_662), .B(n_667), .C(n_676), .Y(n_661) );
AND2x2_ASAP7_75t_L g722 ( .A(n_507), .B(n_528), .Y(n_722) );
INVx5_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g575 ( .A(n_508), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_508), .B(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_508), .B(n_570), .Y(n_582) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_508), .Y(n_584) );
OR2x2_ASAP7_75t_L g595 ( .A(n_508), .B(n_517), .Y(n_595) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_508), .B(n_586), .Y(n_600) );
AND2x2_ASAP7_75t_L g625 ( .A(n_508), .B(n_517), .Y(n_625) );
AND2x2_ASAP7_75t_L g645 ( .A(n_508), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g683 ( .A(n_508), .B(n_516), .Y(n_683) );
OR2x2_ASAP7_75t_L g686 ( .A(n_508), .B(n_672), .Y(n_686) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_517), .A2(n_630), .B(n_633), .C(n_639), .Y(n_629) );
INVx5_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_518), .B(n_528), .Y(n_560) );
AND2x2_ASAP7_75t_L g564 ( .A(n_518), .B(n_529), .Y(n_564) );
OR2x2_ASAP7_75t_L g570 ( .A(n_518), .B(n_528), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_SL g587 ( .A(n_528), .Y(n_587) );
OR2x2_ASAP7_75t_L g715 ( .A(n_528), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_555), .B(n_558), .C(n_567), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI31xp33_ASAP7_75t_L g640 ( .A1(n_538), .A2(n_641), .A3(n_643), .B(n_644), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_539), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_540), .B(n_571), .Y(n_577) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_541), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g597 ( .A(n_541), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g602 ( .A(n_541), .B(n_572), .Y(n_602) );
AND2x2_ASAP7_75t_L g612 ( .A(n_541), .B(n_571), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_541), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g632 ( .A(n_541), .B(n_589), .Y(n_632) );
AND2x2_ASAP7_75t_L g637 ( .A(n_541), .B(n_609), .Y(n_637) );
OR2x2_ASAP7_75t_L g656 ( .A(n_541), .B(n_543), .Y(n_656) );
OR2x2_ASAP7_75t_L g658 ( .A(n_541), .B(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_541), .Y(n_705) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g605 ( .A(n_543), .B(n_572), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_543), .B(n_589), .Y(n_628) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g574 ( .A(n_545), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .Y(n_546) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g665 ( .A(n_557), .B(n_589), .Y(n_665) );
AOI322xp5_ASAP7_75t_L g667 ( .A1(n_557), .A2(n_571), .A3(n_609), .B1(n_668), .B2(n_669), .C1(n_670), .C2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g675 ( .A(n_557), .Y(n_675) );
NAND2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVx1_ASAP7_75t_SL g669 ( .A(n_559), .Y(n_669) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
OR2x2_ASAP7_75t_L g621 ( .A(n_560), .B(n_566), .Y(n_621) );
INVx1_ASAP7_75t_L g652 ( .A(n_560), .Y(n_652) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI32xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .A3(n_573), .B1(n_575), .B2(n_577), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AOI21xp33_ASAP7_75t_SL g607 ( .A1(n_570), .A2(n_585), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g622 ( .A(n_571), .Y(n_622) );
AND2x4_ASAP7_75t_L g619 ( .A(n_572), .B(n_589), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_572), .B(n_655), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g684 ( .A1(n_573), .A2(n_600), .A3(n_619), .B1(n_652), .B2(n_685), .C1(n_687), .C2(n_688), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_573), .A2(n_650), .B1(n_714), .B2(n_715), .C(n_717), .Y(n_713) );
AND2x2_ASAP7_75t_L g601 ( .A(n_574), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g581 ( .A(n_576), .Y(n_581) );
OR2x2_ASAP7_75t_L g653 ( .A(n_576), .B(n_638), .Y(n_653) );
OAI31xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .A3(n_583), .B(n_588), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_579), .A2(n_612), .B1(n_613), .B2(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g624 ( .A(n_581), .B(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_583), .A2(n_624), .B1(n_677), .B2(n_680), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g666 ( .A(n_586), .B(n_635), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_586), .B(n_625), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_587), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g700 ( .A(n_587), .B(n_638), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_588), .A2(n_683), .B1(n_696), .B2(n_699), .Y(n_695) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g604 ( .A(n_589), .Y(n_604) );
AND2x2_ASAP7_75t_L g687 ( .A(n_589), .B(n_609), .Y(n_687) );
OR2x2_ASAP7_75t_L g689 ( .A(n_589), .B(n_656), .Y(n_689) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_589), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_590), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_590), .B(n_635), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B(n_599), .C(n_611), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B1(n_603), .B2(n_606), .C(n_607), .Y(n_599) );
INVxp67_ASAP7_75t_L g711 ( .A(n_602), .Y(n_711) );
INVx1_ASAP7_75t_L g678 ( .A(n_603), .Y(n_678) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g642 ( .A(n_604), .B(n_609), .Y(n_642) );
INVx1_ASAP7_75t_L g659 ( .A(n_605), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_605), .B(n_632), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g674 ( .A(n_609), .Y(n_674) );
AND2x2_ASAP7_75t_L g680 ( .A(n_609), .B(n_635), .Y(n_680) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_SL g668 ( .A(n_616), .Y(n_668) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_619), .B(n_655), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_623), .B2(n_626), .C(n_629), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g716 ( .A(n_625), .Y(n_716) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g634 ( .A(n_628), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_632), .B(n_691), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_638), .Y(n_633) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_636), .A2(n_682), .B(n_684), .C(n_690), .Y(n_681) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g693 ( .A(n_638), .Y(n_693) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI222xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B1(n_653), .B2(n_654), .C1(n_657), .C2(n_658), .Y(n_647) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g723 ( .A(n_654), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_655), .B(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_655), .A2(n_702), .B1(n_704), .B2(n_707), .Y(n_701) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
NOR4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_681), .C(n_694), .D(n_713), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_663), .B(n_693), .Y(n_703) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g670 ( .A(n_668), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_671), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_701), .C(n_708), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx2_ASAP7_75t_L g710 ( .A(n_706), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
OAI21xp5_ASAP7_75t_SL g717 ( .A1(n_718), .A2(n_720), .B(n_723), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g731 ( .A(n_724), .Y(n_731) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_752), .B(n_753), .Y(n_741) );
XOR2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule