module fake_netlist_1_5095_n_483 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_483);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_483;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g69 ( .A(n_56), .Y(n_69) );
INVxp33_ASAP7_75t_SL g70 ( .A(n_55), .Y(n_70) );
CKINVDCx20_ASAP7_75t_R g71 ( .A(n_3), .Y(n_71) );
BUFx2_ASAP7_75t_L g72 ( .A(n_51), .Y(n_72) );
INVx1_ASAP7_75t_SL g73 ( .A(n_26), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_17), .Y(n_74) );
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_11), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_11), .Y(n_76) );
INVxp67_ASAP7_75t_L g77 ( .A(n_5), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_36), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_0), .Y(n_79) );
INVx1_ASAP7_75t_SL g80 ( .A(n_14), .Y(n_80) );
BUFx2_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_58), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_53), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_5), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_57), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_10), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_14), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_33), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_52), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_31), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_28), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_3), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_45), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_64), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_44), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_20), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_34), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_72), .B(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_69), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_72), .B(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_81), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_81), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_74), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_75), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_78), .B(n_98), .Y(n_110) );
INVx6_ASAP7_75t_L g111 ( .A(n_100), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_76), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_70), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_98), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_84), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_92), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_91), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_95), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_102), .B(n_99), .Y(n_124) );
INVx8_ASAP7_75t_L g125 ( .A(n_101), .Y(n_125) );
INVx5_ASAP7_75t_L g126 ( .A(n_113), .Y(n_126) );
AND3x4_ASAP7_75t_L g127 ( .A(n_118), .B(n_91), .C(n_71), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_113), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_101), .B(n_99), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_108), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_113), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_115), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_104), .B(n_87), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_107), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_111), .B(n_87), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_103), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_111), .B(n_88), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_117), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_128), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_135), .B(n_111), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_138), .A2(n_122), .B(n_110), .C(n_121), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
INVxp67_ASAP7_75t_SL g159 ( .A(n_146), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_130), .B(n_111), .Y(n_161) );
INVx1_ASAP7_75t_SL g162 ( .A(n_125), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_137), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_146), .B(n_111), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_130), .B(n_105), .Y(n_165) );
NOR2xp33_ASAP7_75t_R g166 ( .A(n_141), .B(n_109), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_146), .B(n_106), .Y(n_167) );
NOR3xp33_ASAP7_75t_SL g168 ( .A(n_124), .B(n_114), .C(n_123), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_129), .B(n_120), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_136), .B(n_121), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_140), .B(n_122), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_140), .B(n_96), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_141), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_138), .B(n_97), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_125), .Y(n_178) );
NOR2xp33_ASAP7_75t_R g179 ( .A(n_125), .B(n_97), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_136), .B(n_79), .Y(n_181) );
OR2x6_ASAP7_75t_L g182 ( .A(n_125), .B(n_94), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_129), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_165), .B(n_129), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_182), .A2(n_127), .B1(n_136), .B2(n_149), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_182), .A2(n_127), .B1(n_136), .B2(n_139), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_182), .A2(n_127), .B1(n_149), .B2(n_148), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_172), .B(n_139), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_165), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_176), .B(n_144), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_150), .A2(n_148), .B(n_142), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_158), .B(n_144), .Y(n_194) );
INVxp67_ASAP7_75t_L g195 ( .A(n_161), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_182), .A2(n_145), .B1(n_143), .B2(n_142), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_172), .B(n_147), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_166), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_180), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_172), .B(n_147), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_170), .B(n_143), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_178), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
BUFx8_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_155), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_205), .B(n_183), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_205), .A2(n_183), .B1(n_162), .B2(n_178), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_190), .B(n_162), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_212), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_184), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_200), .B(n_172), .Y(n_220) );
OAI211xp5_ASAP7_75t_L g221 ( .A1(n_189), .A2(n_154), .B(n_168), .C(n_167), .Y(n_221) );
CKINVDCx11_ASAP7_75t_R g222 ( .A(n_201), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_200), .B(n_181), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_191), .A2(n_161), .B1(n_167), .B2(n_173), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_184), .Y(n_226) );
BUFx12f_ASAP7_75t_L g227 ( .A(n_212), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_186), .A2(n_181), .B1(n_159), .B2(n_175), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_196), .Y(n_229) );
AOI222xp33_ASAP7_75t_L g230 ( .A1(n_188), .A2(n_181), .B1(n_80), .B2(n_88), .C1(n_79), .C2(n_85), .Y(n_230) );
NOR2x1_ASAP7_75t_SL g231 ( .A(n_196), .B(n_153), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_189), .B(n_164), .C(n_153), .Y(n_234) );
BUFx12f_ASAP7_75t_L g235 ( .A(n_212), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_186), .A2(n_181), .B1(n_179), .B2(n_160), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_212), .A2(n_124), .B1(n_164), .B2(n_177), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_211), .A2(n_145), .B1(n_160), .B2(n_147), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_227), .A2(n_211), .B1(n_209), .B2(n_206), .Y(n_239) );
INVx5_ASAP7_75t_SL g240 ( .A(n_215), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_219), .B(n_192), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_229), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_218), .B(n_197), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_226), .A2(n_195), .B1(n_190), .B2(n_192), .C(n_207), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_232), .A2(n_194), .B1(n_177), .B2(n_185), .C(n_187), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_235), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_236), .A2(n_235), .B1(n_218), .B2(n_230), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_220), .Y(n_249) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_233), .A2(n_194), .B1(n_185), .B2(n_187), .C(n_202), .Y(n_250) );
OAI22xp5_ASAP7_75t_SL g251 ( .A1(n_237), .A2(n_199), .B1(n_206), .B2(n_209), .Y(n_251) );
OAI21xp33_ASAP7_75t_SL g252 ( .A1(n_238), .A2(n_202), .B(n_204), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_220), .B(n_197), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_211), .B1(n_194), .B2(n_204), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_217), .A2(n_194), .B1(n_210), .B2(n_198), .Y(n_255) );
NAND2x1_ASAP7_75t_L g256 ( .A(n_224), .B(n_198), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_221), .A2(n_193), .B(n_213), .C(n_208), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
OAI221xp5_ASAP7_75t_SL g259 ( .A1(n_225), .A2(n_85), .B1(n_94), .B2(n_83), .C(n_89), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_248), .A2(n_217), .B1(n_223), .B2(n_215), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_244), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_253), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_244), .B(n_215), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_258), .Y(n_264) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_257), .A2(n_234), .B(n_231), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_242), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_253), .Y(n_268) );
OAI211xp5_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_222), .B(n_228), .C(n_89), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_247), .Y(n_270) );
AOI33xp33_ASAP7_75t_L g271 ( .A1(n_249), .A2(n_86), .A3(n_90), .B1(n_93), .B2(n_223), .B3(n_73), .Y(n_271) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_257), .B(n_86), .C(n_90), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_258), .Y(n_273) );
OAI211xp5_ASAP7_75t_L g274 ( .A1(n_239), .A2(n_222), .B(n_93), .C(n_132), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_241), .B(n_224), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_247), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_259), .B(n_224), .C(n_229), .Y(n_277) );
AOI222xp33_ASAP7_75t_L g278 ( .A1(n_246), .A2(n_213), .B1(n_216), .B2(n_131), .C1(n_132), .C2(n_208), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_243), .B(n_229), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_251), .A2(n_196), .B1(n_210), .B2(n_133), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_240), .A2(n_196), .B1(n_210), .B2(n_214), .Y(n_281) );
OAI22xp5_ASAP7_75t_SL g282 ( .A1(n_242), .A2(n_229), .B1(n_214), .B2(n_131), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_247), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_262), .B(n_240), .Y(n_284) );
OAI31xp33_ASAP7_75t_L g285 ( .A1(n_269), .A2(n_254), .A3(n_255), .B(n_134), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_262), .B(n_240), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_261), .B(n_240), .Y(n_288) );
OAI31xp33_ASAP7_75t_SL g289 ( .A1(n_274), .A2(n_250), .A3(n_252), .B(n_4), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_273), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_260), .A2(n_133), .B1(n_256), .B2(n_128), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_268), .B(n_243), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_264), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_266), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_268), .B(n_243), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_265), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_263), .B(n_243), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_280), .A2(n_133), .B1(n_243), .B2(n_134), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_126), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_275), .B(n_126), .Y(n_303) );
AOI221x1_ASAP7_75t_L g304 ( .A1(n_272), .A2(n_133), .B1(n_171), .B2(n_157), .C(n_156), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_263), .B(n_134), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_265), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_267), .A2(n_126), .B1(n_171), .B2(n_157), .C(n_156), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_270), .B(n_1), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_283), .Y(n_310) );
OAI21xp33_ASAP7_75t_L g311 ( .A1(n_271), .A2(n_174), .B(n_171), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_265), .B(n_126), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_272), .B(n_126), .C(n_157), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_265), .Y(n_314) );
OAI21xp5_ASAP7_75t_SL g315 ( .A1(n_278), .A2(n_2), .B(n_6), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
NAND4xp25_ASAP7_75t_L g317 ( .A(n_278), .B(n_6), .C(n_7), .D(n_8), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_290), .B(n_276), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_293), .B(n_279), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_293), .B(n_279), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_297), .B(n_270), .Y(n_322) );
OAI211xp5_ASAP7_75t_SL g323 ( .A1(n_289), .A2(n_277), .B(n_281), .C(n_276), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_291), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_310), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_315), .A2(n_276), .B1(n_270), .B2(n_277), .C(n_126), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_286), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_291), .B(n_7), .Y(n_329) );
INVx4_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_295), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_296), .B(n_8), .Y(n_332) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_296), .B(n_174), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_294), .B(n_9), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g337 ( .A(n_299), .B(n_9), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_297), .B(n_10), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_300), .B(n_12), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_298), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_284), .B(n_12), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_284), .B(n_287), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_317), .B(n_13), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_305), .B(n_13), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_300), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_15), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_299), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_307), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_302), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_307), .B(n_15), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_287), .B(n_16), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_302), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_316), .B(n_16), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_312), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_316), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_126), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_318), .B(n_18), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_303), .B(n_19), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_288), .B(n_21), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_288), .B(n_22), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_344), .A2(n_327), .B1(n_359), .B2(n_323), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_335), .A2(n_313), .B(n_304), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_359), .B(n_306), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_357), .B(n_306), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_326), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_351), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_319), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_331), .B(n_292), .Y(n_374) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_352), .A2(n_313), .B1(n_311), .B2(n_301), .C1(n_308), .C2(n_285), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_351), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_330), .A2(n_311), .B1(n_174), .B2(n_156), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_342), .A2(n_152), .B1(n_304), .B2(n_25), .C(n_27), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g379 ( .A1(n_350), .A2(n_23), .B(n_24), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_346), .B(n_29), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_335), .A2(n_152), .B(n_32), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_325), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_346), .B(n_30), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_335), .B(n_152), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_352), .B(n_35), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_320), .B(n_37), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_340), .A2(n_38), .B(n_39), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_338), .B(n_40), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_338), .B(n_361), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
OAI22xp33_ASAP7_75t_SL g394 ( .A1(n_329), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_332), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_337), .A2(n_46), .B(n_48), .C(n_49), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_336), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_355), .B(n_50), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_340), .B(n_54), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_329), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g402 ( .A1(n_337), .A2(n_59), .B(n_60), .C(n_61), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_353), .B(n_68), .C(n_63), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_339), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_358), .B(n_66), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_324), .Y(n_406) );
OAI21xp33_ASAP7_75t_SL g407 ( .A1(n_330), .A2(n_62), .B(n_65), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_354), .B(n_362), .C(n_347), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_330), .A2(n_364), .B1(n_343), .B2(n_363), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_376), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_367), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_385), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_371), .B(n_320), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_408), .B(n_330), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_401), .B(n_341), .Y(n_418) );
NOR3xp33_ASAP7_75t_SL g419 ( .A(n_407), .B(n_365), .C(n_341), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_372), .Y(n_420) );
XNOR2x1_ASAP7_75t_L g421 ( .A(n_409), .B(n_321), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_366), .A2(n_362), .B1(n_360), .B2(n_347), .C(n_345), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_404), .Y(n_424) );
NOR3xp33_ASAP7_75t_SL g425 ( .A(n_379), .B(n_334), .C(n_364), .Y(n_425) );
NOR3xp33_ASAP7_75t_SL g426 ( .A(n_390), .B(n_334), .C(n_364), .Y(n_426) );
XNOR2xp5_ASAP7_75t_L g427 ( .A(n_392), .B(n_322), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_386), .B(n_322), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_373), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_395), .B(n_345), .Y(n_430) );
NAND2xp33_ASAP7_75t_SL g431 ( .A(n_387), .B(n_366), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_397), .A2(n_364), .B(n_363), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_393), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_398), .B(n_349), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_367), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_370), .B(n_360), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_369), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_370), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_431), .A2(n_374), .B1(n_389), .B2(n_375), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_414), .B(n_394), .C(n_378), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_439), .B(n_349), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_423), .B(n_356), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_438), .B(n_356), .Y(n_445) );
NAND2xp33_ASAP7_75t_SL g446 ( .A(n_426), .B(n_387), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_414), .B(n_432), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_410), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_SL g450 ( .A1(n_412), .A2(n_381), .B(n_384), .C(n_399), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_435), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_421), .B(n_400), .Y(n_452) );
AOI31xp33_ASAP7_75t_L g453 ( .A1(n_420), .A2(n_382), .A3(n_368), .B(n_402), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_415), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
OAI221xp5_ASAP7_75t_SL g457 ( .A1(n_422), .A2(n_391), .B1(n_377), .B2(n_402), .C(n_397), .Y(n_457) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_447), .A2(n_437), .B1(n_433), .B2(n_430), .C1(n_428), .C2(n_429), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_448), .B(n_427), .Y(n_459) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_440), .B(n_413), .Y(n_460) );
AOI21xp33_ASAP7_75t_L g461 ( .A1(n_450), .A2(n_437), .B(n_388), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_441), .A2(n_426), .B1(n_419), .B2(n_425), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_442), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_445), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_441), .A2(n_425), .B(n_419), .C(n_433), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_444), .Y(n_466) );
NOR4xp25_ASAP7_75t_L g467 ( .A(n_457), .B(n_405), .C(n_418), .D(n_434), .Y(n_467) );
OAI311xp33_ASAP7_75t_L g468 ( .A1(n_453), .A2(n_403), .A3(n_436), .B1(n_333), .C1(n_328), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_452), .A2(n_328), .B1(n_333), .B2(n_446), .C(n_455), .Y(n_469) );
OAI22x1_ASAP7_75t_L g470 ( .A1(n_452), .A2(n_454), .B1(n_456), .B2(n_451), .Y(n_470) );
OA22x2_ASAP7_75t_L g471 ( .A1(n_449), .A2(n_440), .B1(n_448), .B2(n_410), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_447), .B(n_443), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_471), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_459), .Y(n_474) );
OR2x6_ASAP7_75t_L g475 ( .A(n_465), .B(n_470), .Y(n_475) );
AND3x2_ASAP7_75t_L g476 ( .A(n_467), .B(n_469), .C(n_472), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_474), .Y(n_477) );
NAND4xp75_ASAP7_75t_L g478 ( .A(n_473), .B(n_462), .C(n_461), .D(n_467), .Y(n_478) );
XNOR2xp5_ASAP7_75t_L g479 ( .A(n_478), .B(n_460), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_477), .Y(n_480) );
OR3x2_ASAP7_75t_L g481 ( .A(n_479), .B(n_475), .C(n_476), .Y(n_481) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_481), .A2(n_480), .B(n_458), .C(n_475), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_482), .A2(n_468), .B1(n_464), .B2(n_466), .C(n_463), .Y(n_483) );
endmodule