module fake_jpeg_13075_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_0),
.B(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_43),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_16),
.C(n_15),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_5),
.C(n_6),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_24),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_57),
.Y(n_82)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_61),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_64),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_67),
.Y(n_91)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_4),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_73),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_25),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_37),
.B1(n_38),
.B2(n_21),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_86),
.A2(n_88),
.B1(n_108),
.B2(n_119),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_17),
.B1(n_38),
.B2(n_31),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_11),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_41),
.A2(n_16),
.B1(n_31),
.B2(n_21),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_103),
.B1(n_110),
.B2(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_44),
.A2(n_47),
.B1(n_68),
.B2(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_91),
.B1(n_111),
.B2(n_109),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_15),
.B1(n_17),
.B2(n_40),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_112),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_59),
.A2(n_36),
.B1(n_25),
.B2(n_28),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_65),
.B1(n_70),
.B2(n_56),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_58),
.A2(n_36),
.B1(n_28),
.B2(n_7),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_82),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_55),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_132),
.Y(n_169)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_116),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_80),
.B(n_85),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_93),
.B(n_81),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_113),
.Y(n_156)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_110),
.B1(n_103),
.B2(n_97),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_153),
.B(n_127),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_139),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_94),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_90),
.B(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_85),
.B1(n_105),
.B2(n_111),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_150),
.B1(n_151),
.B2(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_80),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_152),
.Y(n_159)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_98),
.A2(n_87),
.B1(n_94),
.B2(n_96),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_89),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_113),
.B1(n_95),
.B2(n_105),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_113),
.B(n_134),
.C(n_130),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_163),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_173),
.B1(n_154),
.B2(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_129),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_132),
.A3(n_131),
.B1(n_143),
.B2(n_140),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_176),
.B(n_165),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_121),
.B(n_143),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_136),
.B1(n_144),
.B2(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_177),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_148),
.B(n_141),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_160),
.C(n_162),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_193),
.C(n_194),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_181),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_165),
.B(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_182),
.B1(n_184),
.B2(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_165),
.B(n_174),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_158),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_180),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_156),
.C(n_168),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_206),
.C(n_208),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_185),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_170),
.B(n_169),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_180),
.B(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_178),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_157),
.B1(n_173),
.B2(n_169),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_187),
.B1(n_190),
.B2(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_216),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_199),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_215),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_207),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_218),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_167),
.B1(n_195),
.B2(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_226),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_196),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_203),
.C(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_217),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_232),
.B(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_201),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_198),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_213),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_212),
.B(n_214),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_232),
.Y(n_233)
);

OAI221xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_197),
.C(n_217),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_213),
.B1(n_228),
.B2(n_222),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_204),
.B(n_200),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_225),
.B1(n_219),
.B2(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_222),
.C(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_200),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_242),
.B(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_243),
.B(n_202),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_244),
.Y(n_246)
);


endmodule