module fake_jpeg_17987_n_359 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_42),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_49),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_10),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_20),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_23),
.Y(n_101)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_75),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_38),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_46),
.B1(n_40),
.B2(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_84),
.A2(n_85),
.B1(n_111),
.B2(n_118),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_40),
.B1(n_54),
.B2(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_119),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_101),
.Y(n_123)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_94),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_40),
.B1(n_23),
.B2(n_39),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_105),
.B1(n_29),
.B2(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_33),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_28),
.B1(n_20),
.B2(n_37),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_102),
.Y(n_149)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_55),
.B1(n_49),
.B2(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_25),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_113),
.Y(n_124)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_55),
.B1(n_30),
.B2(n_29),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_28),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g115 ( 
.A(n_69),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_29),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_25),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_132),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_76),
.B1(n_68),
.B2(n_78),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_100),
.B1(n_99),
.B2(n_103),
.Y(n_160)
);

OR2x4_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_95),
.Y(n_145)
);

NOR2x1_ASAP7_75t_R g159 ( 
.A(n_145),
.B(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_105),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_88),
.B(n_31),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_59),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_27),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_83),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_152),
.B(n_154),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_86),
.B1(n_81),
.B2(n_87),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_167),
.B1(n_98),
.B2(n_82),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_89),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_155),
.B(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_108),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_172),
.B1(n_174),
.B2(n_27),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_124),
.B(n_142),
.Y(n_186)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_114),
.B1(n_99),
.B2(n_91),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_112),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_122),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_169),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_36),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_149),
.B(n_125),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_110),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_173),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_82),
.B1(n_97),
.B2(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_21),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_26),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_178),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_16),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

XOR2x2_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_144),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_187),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_132),
.B1(n_148),
.B2(n_126),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_190),
.B1(n_175),
.B2(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_121),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_156),
.C(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_197),
.C(n_201),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_142),
.B1(n_125),
.B2(n_139),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_191),
.B(n_185),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_142),
.B(n_36),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_193),
.A2(n_194),
.B(n_195),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_141),
.C(n_128),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_141),
.C(n_78),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_1),
.B(n_2),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_3),
.B(n_4),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_190),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_162),
.B1(n_157),
.B2(n_136),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_211),
.A2(n_220),
.B1(n_222),
.B2(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_223),
.Y(n_261)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_164),
.B1(n_179),
.B2(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g223 ( 
.A(n_180),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_226),
.B(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_177),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_157),
.C(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_201),
.C(n_204),
.Y(n_246)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_229),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_1),
.B(n_2),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_2),
.B(n_135),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_238),
.B(n_239),
.Y(n_242)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_233),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_241),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_133),
.B1(n_178),
.B2(n_135),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_231),
.B1(n_217),
.B2(n_229),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_194),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_208),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_250),
.C(n_218),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_182),
.C(n_183),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_206),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_35),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_195),
.B(n_193),
.C(n_196),
.D(n_203),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_255),
.B(n_38),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_133),
.Y(n_257)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_237),
.B1(n_230),
.B2(n_222),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_212),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_263),
.B(n_266),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_36),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_68),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_264),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_3),
.B(n_4),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_274),
.C(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_235),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_264),
.C(n_261),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_275),
.A2(n_277),
.B1(n_265),
.B2(n_7),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_226),
.C(n_235),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_238),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_6),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_35),
.C(n_24),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_35),
.C(n_38),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_258),
.C(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_245),
.B1(n_251),
.B2(n_252),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_285),
.A2(n_262),
.B1(n_254),
.B2(n_263),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_291),
.A2(n_293),
.B1(n_294),
.B2(n_300),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_259),
.B1(n_254),
.B2(n_245),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_272),
.A2(n_252),
.B(n_265),
.C(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_267),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_251),
.B1(n_265),
.B2(n_248),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_288),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_306),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_306)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_316),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_314),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_277),
.B(n_276),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_322),
.B(n_294),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_273),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_284),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_320),
.Y(n_323)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_294),
.B1(n_305),
.B2(n_304),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_286),
.C(n_280),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_282),
.B1(n_14),
.B2(n_15),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_304),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_310),
.A2(n_293),
.B(n_294),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_324),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_308),
.A2(n_315),
.B(n_318),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_325),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_309),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_333),
.B1(n_322),
.B2(n_319),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_316),
.C(n_330),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.C(n_338),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_309),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_339),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_320),
.C(n_305),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_312),
.C(n_31),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_31),
.C(n_38),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_31),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_329),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_347),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_337),
.A2(n_324),
.B(n_326),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_346),
.A2(n_348),
.B(n_338),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_16),
.Y(n_348)
);

OAI21x1_ASAP7_75t_L g350 ( 
.A1(n_343),
.A2(n_334),
.B(n_340),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_350),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_349),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_345),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_353),
.B(n_344),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_16),
.B1(n_17),
.B2(n_31),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_357),
.B(n_17),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_38),
.Y(n_359)
);


endmodule