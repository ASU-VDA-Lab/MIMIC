module fake_netlist_1_2448_n_604 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_604);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_604;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_73;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g70 ( .A(n_49), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_14), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_20), .Y(n_72) );
INVxp67_ASAP7_75t_SL g73 ( .A(n_60), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_51), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_33), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_27), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_4), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_1), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_30), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_58), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_52), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_2), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_31), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_26), .Y(n_88) );
NOR2xp67_ASAP7_75t_L g89 ( .A(n_23), .B(n_59), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_21), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_6), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_29), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_22), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_47), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_42), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_8), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_12), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_16), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_21), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_15), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_87), .B(n_0), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_102), .B(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_102), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_90), .Y(n_116) );
AND2x6_ASAP7_75t_L g117 ( .A(n_75), .B(n_36), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_107), .B(n_2), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_107), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_91), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_81), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_93), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_70), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_92), .Y(n_129) );
CKINVDCx6p67_ASAP7_75t_R g130 ( .A(n_91), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_95), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_71), .Y(n_141) );
NOR2xp33_ASAP7_75t_R g142 ( .A(n_96), .B(n_37), .Y(n_142) );
INVx2_ASAP7_75t_SL g143 ( .A(n_85), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_99), .B(n_3), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_91), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_117), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_119), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_121), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_130), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_145), .B(n_71), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_145), .B(n_109), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_110), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_145), .B(n_72), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_143), .B(n_113), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_141), .B(n_72), .Y(n_165) );
AO22x2_ASAP7_75t_L g166 ( .A1(n_115), .A2(n_100), .B1(n_101), .B2(n_105), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_117), .A2(n_77), .B1(n_78), .B2(n_105), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_122), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_128), .B(n_106), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_116), .B(n_77), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_129), .B(n_73), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_117), .A2(n_135), .B1(n_144), .B2(n_134), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_115), .B(n_78), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_120), .B(n_97), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_147), .B(n_104), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
NOR3xp33_ASAP7_75t_L g180 ( .A(n_112), .B(n_84), .C(n_108), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_120), .B(n_99), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_121), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_135), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_117), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_117), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_118), .B(n_104), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_139), .Y(n_190) );
CKINVDCx11_ASAP7_75t_R g191 ( .A(n_146), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_121), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_126), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_126), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_123), .B(n_103), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_123), .B(n_94), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_121), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_124), .B(n_94), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_124), .B(n_94), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_117), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_127), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_131), .B(n_94), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_137), .B(n_98), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_147), .B(n_94), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_187), .B(n_111), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_186), .Y(n_207) );
NOR2x1p5_ASAP7_75t_L g208 ( .A(n_151), .B(n_134), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_199), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_199), .Y(n_210) );
HB1xp67_ASAP7_75t_SL g211 ( .A(n_151), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_191), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_148), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_165), .B(n_133), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_165), .B(n_176), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_172), .B(n_140), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_183), .A2(n_138), .B(n_133), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_187), .B(n_131), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_150), .B(n_138), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_171), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_202), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
INVxp33_ASAP7_75t_L g225 ( .A(n_149), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_165), .B(n_132), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_202), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_203), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_150), .B(n_132), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_176), .B(n_136), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_203), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_187), .B(n_136), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_189), .Y(n_233) );
NOR2x1p5_ASAP7_75t_L g234 ( .A(n_173), .B(n_3), .Y(n_234) );
BUFx8_ASAP7_75t_L g235 ( .A(n_157), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_187), .B(n_89), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_157), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_189), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_157), .A2(n_142), .B1(n_5), .B2(n_6), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_186), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_150), .B(n_41), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_205), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_205), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_156), .B(n_4), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_156), .B(n_5), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_189), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_159), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_176), .B(n_7), .Y(n_249) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_157), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_180), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_178), .B(n_14), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_156), .B(n_16), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_205), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_153), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_153), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_157), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_257) );
INVx4_ASAP7_75t_L g258 ( .A(n_157), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_157), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_158), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_174), .B(n_53), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_166), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_158), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_258), .B(n_201), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_260), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_258), .B(n_259), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_258), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_219), .B(n_196), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_260), .Y(n_270) );
OAI21x1_ASAP7_75t_SL g271 ( .A1(n_259), .A2(n_175), .B(n_167), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_259), .B(n_160), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_238), .B(n_154), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g274 ( .A1(n_213), .A2(n_204), .B1(n_170), .B2(n_160), .Y(n_274) );
NAND2xp33_ASAP7_75t_L g275 ( .A(n_207), .B(n_184), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_219), .B(n_181), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_263), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_224), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_263), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_238), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_245), .Y(n_283) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_245), .B(n_201), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_219), .B(n_181), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_245), .B(n_201), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_225), .B(n_164), .Y(n_288) );
INVx5_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_255), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_256), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_213), .B(n_177), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_246), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_220), .A2(n_184), .B(n_183), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_246), .A2(n_163), .B1(n_161), .B2(n_193), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_206), .B(n_215), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_253), .A2(n_163), .B1(n_161), .B2(n_194), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_253), .B(n_155), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_253), .B(n_206), .Y(n_300) );
BUFx10_ASAP7_75t_L g301 ( .A(n_232), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_207), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
BUFx12f_ASAP7_75t_L g304 ( .A(n_212), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_225), .B(n_194), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_217), .B(n_193), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_240), .B(n_195), .C(n_184), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_207), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_220), .A2(n_184), .B(n_155), .Y(n_310) );
INVx6_ASAP7_75t_L g311 ( .A(n_241), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_269), .A2(n_262), .B1(n_232), .B2(n_234), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_269), .A2(n_209), .B1(n_210), .B2(n_214), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_296), .A2(n_226), .B1(n_243), .B2(n_231), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_274), .A2(n_248), .B1(n_212), .B2(n_237), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_229), .B(n_218), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_304), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_295), .A2(n_230), .B1(n_249), .B2(n_252), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_300), .A2(n_208), .B1(n_237), .B2(n_211), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_293), .A2(n_229), .B(n_184), .Y(n_320) );
BUFx2_ASAP7_75t_R g321 ( .A(n_266), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_292), .B(n_237), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_305), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_295), .A2(n_227), .B1(n_223), .B2(n_257), .Y(n_324) );
OAI21x1_ASAP7_75t_L g325 ( .A1(n_294), .A2(n_242), .B(n_221), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_284), .A2(n_239), .B(n_233), .Y(n_327) );
OR2x6_ASAP7_75t_L g328 ( .A(n_298), .B(n_250), .Y(n_328) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_283), .B(n_243), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_297), .A2(n_251), .B1(n_254), .B2(n_228), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_296), .A2(n_231), .B1(n_243), .B2(n_244), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_288), .A2(n_236), .B1(n_231), .B2(n_261), .C(n_222), .Y(n_332) );
NAND2xp33_ASAP7_75t_R g333 ( .A(n_298), .B(n_300), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_277), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
INVx4_ASAP7_75t_SL g337 ( .A(n_298), .Y(n_337) );
AO31x2_ASAP7_75t_L g338 ( .A1(n_265), .A2(n_247), .A3(n_216), .B(n_239), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_276), .B(n_247), .Y(n_340) );
AOI21x1_ASAP7_75t_L g341 ( .A1(n_328), .A2(n_242), .B(n_308), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_323), .B(n_276), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_329), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_336), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_329), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_328), .A2(n_284), .B1(n_283), .B2(n_300), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_313), .B(n_285), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_315), .A2(n_330), .B1(n_312), .B2(n_322), .Y(n_348) );
AOI21xp33_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_306), .B(n_308), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_306), .B1(n_265), .B2(n_287), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_324), .A2(n_287), .B1(n_307), .B2(n_279), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_326), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
AO21x2_ASAP7_75t_L g354 ( .A1(n_327), .A2(n_271), .B(n_277), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_319), .A2(n_307), .B1(n_287), .B2(n_272), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_334), .Y(n_356) );
BUFx10_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_314), .A2(n_331), .B1(n_332), .B2(n_333), .C(n_340), .Y(n_358) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_337), .A2(n_304), .B1(n_287), .B2(n_272), .C1(n_279), .C2(n_271), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_335), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_316), .A2(n_310), .B(n_272), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_356), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_352), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_353), .B(n_338), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_358), .A2(n_333), .B1(n_321), .B2(n_282), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_350), .B(n_349), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_356), .B(n_337), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_360), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_348), .A2(n_331), .B1(n_290), .B2(n_303), .C(n_299), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_360), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_346), .B(n_338), .Y(n_373) );
NOR2x1p5_ASAP7_75t_L g374 ( .A(n_345), .B(n_268), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_353), .B(n_338), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g376 ( .A(n_359), .B(n_289), .C(n_309), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_352), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_351), .A2(n_325), .B(n_286), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_355), .A2(n_281), .B1(n_280), .B2(n_291), .C(n_320), .Y(n_380) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_341), .A2(n_291), .B(n_216), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_347), .B(n_338), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_361), .B(n_289), .C(n_309), .Y(n_384) );
AO21x2_ASAP7_75t_L g385 ( .A1(n_341), .A2(n_275), .B(n_192), .Y(n_385) );
AO21x1_ASAP7_75t_SL g386 ( .A1(n_343), .A2(n_289), .B(n_301), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_343), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
AOI222xp33_ASAP7_75t_L g390 ( .A1(n_342), .A2(n_357), .B1(n_345), .B2(n_343), .C1(n_267), .C2(n_289), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_364), .B(n_354), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_376), .B(n_345), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_390), .B(n_289), .C(n_286), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_354), .B1(n_357), .B2(n_309), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_383), .B(n_354), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_383), .B(n_19), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_368), .B(n_20), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_368), .B(n_25), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_366), .B(n_286), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_286), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_373), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_389), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_366), .B(n_379), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_387), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_371), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_367), .B(n_286), .Y(n_419) );
AO21x2_ASAP7_75t_L g420 ( .A1(n_378), .A2(n_152), .B(n_168), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_371), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_379), .B(n_302), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_376), .A2(n_273), .B1(n_267), .B2(n_311), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_369), .B(n_302), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_387), .B(n_302), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_367), .B(n_28), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_370), .A2(n_357), .B1(n_309), .B2(n_302), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_382), .B(n_34), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_382), .B(n_309), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_389), .B(n_302), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_384), .Y(n_432) );
INVx4_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_377), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_388), .B(n_35), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_377), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_411), .B(n_381), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_393), .B(n_390), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_406), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_411), .B(n_381), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_397), .B(n_381), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_397), .B(n_381), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_413), .B(n_385), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_398), .B(n_374), .Y(n_446) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_395), .A2(n_380), .B(n_190), .C(n_169), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_409), .B(n_385), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_433), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_398), .B(n_38), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_402), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_410), .B(n_386), .Y(n_453) );
OR2x6_ASAP7_75t_L g454 ( .A(n_393), .B(n_374), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_410), .B(n_44), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_391), .B(n_386), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_391), .B(n_45), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_402), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_412), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_396), .B(n_46), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_399), .B(n_48), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_416), .B(n_54), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_399), .B(n_404), .Y(n_464) );
NOR4xp25_ASAP7_75t_SL g465 ( .A(n_412), .B(n_55), .C(n_56), .D(n_57), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_437), .B(n_415), .Y(n_466) );
NAND4xp25_ASAP7_75t_L g467 ( .A(n_395), .B(n_179), .C(n_188), .D(n_185), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_424), .B(n_62), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_415), .B(n_63), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_407), .B(n_426), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_400), .B(n_64), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_426), .B(n_67), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_405), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_414), .B(n_68), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_433), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_414), .B(n_152), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_401), .Y(n_478) );
INVxp33_ASAP7_75t_L g479 ( .A(n_392), .Y(n_479) );
XNOR2x1_ASAP7_75t_L g480 ( .A(n_392), .B(n_267), .Y(n_480) );
NAND2xp33_ASAP7_75t_SL g481 ( .A(n_423), .B(n_264), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_433), .B(n_162), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_422), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_432), .B(n_182), .C(n_192), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_400), .B(n_182), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_419), .B(n_197), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_450), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_454), .A2(n_427), .B1(n_423), .B2(n_433), .Y(n_489) );
OAI322xp33_ASAP7_75t_L g490 ( .A1(n_440), .A2(n_432), .A3(n_436), .B1(n_419), .B2(n_421), .C1(n_434), .C2(n_400), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_446), .B(n_435), .Y(n_491) );
AO22x1_ASAP7_75t_L g492 ( .A1(n_476), .A2(n_436), .B1(n_435), .B2(n_429), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_463), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_466), .B(n_421), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_456), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_466), .B(n_421), .Y(n_498) );
OAI21xp33_ASAP7_75t_L g499 ( .A1(n_479), .A2(n_430), .B(n_434), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_464), .B(n_417), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_452), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_454), .A2(n_480), .B1(n_476), .B2(n_451), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_449), .Y(n_503) );
AOI21xp33_ASAP7_75t_SL g504 ( .A1(n_480), .A2(n_431), .B(n_425), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_483), .Y(n_505) );
NAND2x1p5_ASAP7_75t_L g506 ( .A(n_449), .B(n_469), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_453), .B(n_403), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_R g508 ( .A1(n_475), .A2(n_403), .B(n_418), .C(n_417), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_449), .B(n_403), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_456), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_471), .B(n_428), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_474), .B(n_418), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_443), .B(n_408), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_458), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_441), .B(n_420), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_479), .A2(n_273), .A3(n_198), .B(n_420), .Y(n_517) );
AOI21xp33_ASAP7_75t_SL g518 ( .A1(n_473), .A2(n_420), .B(n_273), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_482), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_438), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_444), .A2(n_198), .B(n_420), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_447), .A2(n_241), .B(n_197), .Y(n_522) );
OAI22xp33_ASAP7_75t_L g523 ( .A1(n_467), .A2(n_241), .B1(n_197), .B2(n_200), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_448), .B(n_197), .Y(n_524) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_445), .A2(n_241), .B(n_197), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_448), .B(n_197), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_478), .B(n_197), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_487), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_502), .A2(n_461), .B(n_455), .C(n_460), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_505), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_496), .B(n_470), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_497), .Y(n_532) );
NOR2xp33_ASAP7_75t_R g533 ( .A(n_503), .B(n_481), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_488), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_519), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_501), .Y(n_536) );
XOR2x2_ASAP7_75t_L g537 ( .A(n_502), .B(n_469), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_520), .B(n_438), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g539 ( .A1(n_504), .A2(n_457), .B(n_481), .C(n_465), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_493), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_513), .B(n_442), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_514), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_500), .B(n_442), .Y(n_543) );
XOR2xp5_ASAP7_75t_L g544 ( .A(n_506), .B(n_468), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_507), .B(n_472), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_515), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_494), .B(n_472), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_498), .Y(n_548) );
XNOR2xp5_ASAP7_75t_L g549 ( .A(n_510), .B(n_462), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_511), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_495), .B(n_477), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_512), .B(n_485), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_503), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_509), .Y(n_554) );
AOI22x1_ASAP7_75t_L g555 ( .A1(n_544), .A2(n_506), .B1(n_519), .B2(n_516), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_533), .B(n_518), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_550), .Y(n_557) );
OA22x2_ASAP7_75t_L g558 ( .A1(n_549), .A2(n_489), .B1(n_492), .B2(n_499), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_541), .B(n_516), .Y(n_559) );
AOI21xp33_ASAP7_75t_SL g560 ( .A1(n_549), .A2(n_517), .B(n_523), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_528), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_529), .A2(n_491), .B(n_521), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_544), .A2(n_525), .B1(n_526), .B2(n_524), .Y(n_563) );
XNOR2x1_ASAP7_75t_L g564 ( .A(n_537), .B(n_482), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_533), .B(n_508), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_537), .A2(n_527), .B1(n_482), .B2(n_486), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_530), .B(n_490), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_531), .A2(n_484), .B1(n_522), .B2(n_200), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_539), .A2(n_200), .B(n_241), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_538), .B(n_200), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_534), .Y(n_571) );
OA21x2_ASAP7_75t_L g572 ( .A1(n_554), .A2(n_200), .B(n_553), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_548), .B(n_547), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_540), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_567), .B(n_543), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_564), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_567), .B(n_565), .C(n_569), .Y(n_577) );
AO22x2_ASAP7_75t_L g578 ( .A1(n_556), .A2(n_535), .B1(n_532), .B2(n_536), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_561), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_557), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_558), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_558), .Y(n_582) );
NAND3xp33_ASAP7_75t_SL g583 ( .A(n_556), .B(n_545), .C(n_551), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_562), .A2(n_552), .B(n_532), .Y(n_584) );
OA22x2_ASAP7_75t_L g585 ( .A1(n_566), .A2(n_542), .B1(n_546), .B2(n_559), .Y(n_585) );
AOI221x1_ASAP7_75t_L g586 ( .A1(n_560), .A2(n_542), .B1(n_571), .B2(n_574), .C(n_563), .Y(n_586) );
OA22x2_ASAP7_75t_L g587 ( .A1(n_573), .A2(n_555), .B1(n_568), .B2(n_570), .Y(n_587) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_572), .A2(n_569), .B(n_556), .C(n_562), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_572), .A2(n_558), .B1(n_537), .B2(n_567), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_565), .A2(n_567), .B(n_569), .C(n_556), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_576), .Y(n_591) );
OR3x2_ASAP7_75t_L g592 ( .A(n_582), .B(n_581), .C(n_590), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_582), .B(n_575), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_580), .B(n_577), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_579), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_594), .A2(n_589), .B(n_586), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_594), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_592), .A2(n_588), .B(n_583), .C(n_584), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_597), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_596), .Y(n_600) );
AOI22xp5_ASAP7_75t_SL g601 ( .A1(n_599), .A2(n_591), .B1(n_593), .B2(n_587), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_600), .A2(n_598), .B1(n_593), .B2(n_578), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_602), .A2(n_578), .B1(n_585), .B2(n_595), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_603), .A2(n_601), .B(n_578), .Y(n_604) );
endmodule