module fake_jpeg_1059_n_522 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_522);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_522;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_61),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_67),
.Y(n_119)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_6),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_76),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_87),
.Y(n_117)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_35),
.B(n_6),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_34),
.B(n_6),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_42),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_46),
.A2(n_44),
.B1(n_28),
.B2(n_27),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_102),
.A2(n_145),
.B1(n_15),
.B2(n_89),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_36),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_130),
.B(n_131),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_67),
.B(n_42),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_55),
.B(n_29),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_59),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_50),
.B(n_27),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_146),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_86),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_155),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_60),
.A2(n_29),
.B1(n_23),
.B2(n_39),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_69),
.B(n_15),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_93),
.B(n_20),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_88),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_47),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_46),
.B(n_20),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_92),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_28),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_163),
.B(n_183),
.Y(n_215)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_78),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_73),
.B1(n_75),
.B2(n_72),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_176),
.B1(n_194),
.B2(n_83),
.Y(n_228)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_170),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_175),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_102),
.A2(n_81),
.B1(n_84),
.B2(n_79),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_23),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_126),
.B(n_66),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_195),
.C(n_112),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_38),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_193),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_120),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_52),
.B1(n_45),
.B2(n_58),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_133),
.B(n_68),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_132),
.B(n_38),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_198),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_111),
.B(n_112),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_203),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_114),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_49),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_124),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_161),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_156),
.B1(n_118),
.B2(n_107),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_229),
.B1(n_237),
.B2(n_243),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_242),
.B1(n_202),
.B2(n_170),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_230),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_168),
.A2(n_107),
.B1(n_118),
.B2(n_135),
.Y(n_229)
);

AOI32xp33_ASAP7_75t_L g235 ( 
.A1(n_165),
.A2(n_153),
.A3(n_158),
.B1(n_154),
.B2(n_139),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_150),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_135),
.B1(n_151),
.B2(n_100),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_151),
.B1(n_134),
.B2(n_129),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_228),
.B1(n_243),
.B2(n_237),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_201),
.A2(n_158),
.B1(n_154),
.B2(n_147),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_183),
.A2(n_129),
.B1(n_134),
.B2(n_115),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_162),
.B1(n_203),
.B2(n_199),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_221),
.Y(n_246)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_247),
.A2(n_261),
.B1(n_266),
.B2(n_177),
.Y(n_289)
);

CKINVDCx12_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_195),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_171),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_253),
.A2(n_233),
.B1(n_232),
.B2(n_211),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_196),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_226),
.B(n_196),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_216),
.A2(n_163),
.B1(n_185),
.B2(n_186),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_271),
.B1(n_273),
.B2(n_212),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_220),
.A2(n_150),
.B1(n_173),
.B2(n_201),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_179),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_186),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_265),
.B(n_268),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_229),
.A2(n_190),
.B1(n_180),
.B2(n_164),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_219),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_184),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_125),
.B1(n_139),
.B2(n_109),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_224),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_175),
.B(n_209),
.C(n_192),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_230),
.B1(n_227),
.B2(n_223),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_281),
.B1(n_290),
.B2(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_172),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_215),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_280),
.B(n_136),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_235),
.B(n_214),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_259),
.B(n_262),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_288),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_250),
.B1(n_252),
.B2(n_268),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_297),
.B1(n_300),
.B2(n_302),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_256),
.A2(n_211),
.B1(n_210),
.B2(n_217),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_250),
.A2(n_166),
.B1(n_167),
.B2(n_208),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_249),
.A2(n_258),
.B1(n_269),
.B2(n_265),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_301),
.A2(n_255),
.B1(n_270),
.B2(n_241),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_217),
.B1(n_213),
.B2(n_219),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_263),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_245),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_320),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_306),
.A2(n_312),
.B(n_334),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_329),
.Y(n_335)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_308),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_257),
.B(n_254),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_310),
.C(n_314),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_286),
.B(n_279),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_261),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_313),
.C(n_315),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_274),
.B(n_248),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_225),
.C(n_209),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_240),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_239),
.C(n_240),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_297),
.B(n_267),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_316),
.B(n_322),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_283),
.A2(n_260),
.B(n_222),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_239),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_315),
.C(n_304),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_287),
.Y(n_336)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_222),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_204),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_333),
.Y(n_341)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_330),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_299),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_275),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_275),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_272),
.B(n_246),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_342),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_321),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_338),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_334),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_318),
.A2(n_300),
.B1(n_302),
.B2(n_292),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_326),
.B1(n_312),
.B2(n_331),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_316),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_363),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_178),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_328),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_292),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_353),
.B(n_356),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_182),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_306),
.A2(n_298),
.B1(n_299),
.B2(n_284),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_357),
.A2(n_272),
.B1(n_246),
.B2(n_264),
.Y(n_382)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_362),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_284),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_364),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_365),
.B(n_298),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_313),
.C(n_319),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_372),
.C(n_380),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_341),
.Y(n_367)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_311),
.C(n_330),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_326),
.Y(n_373)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_382),
.B1(n_388),
.B2(n_390),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_345),
.A2(n_352),
.B1(n_351),
.B2(n_349),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_375),
.A2(n_379),
.B1(n_343),
.B2(n_358),
.Y(n_410)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_351),
.A2(n_317),
.B1(n_305),
.B2(n_287),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_305),
.C(n_148),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_SL g381 ( 
.A(n_359),
.B(n_349),
.C(n_355),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_381),
.B(n_385),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_144),
.C(n_109),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_384),
.C(n_364),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_101),
.C(n_270),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_335),
.B(n_236),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_264),
.B1(n_213),
.B2(n_241),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_98),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_357),
.A2(n_200),
.B1(n_125),
.B2(n_159),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_241),
.B(n_174),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_394),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_172),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_382),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_400),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_373),
.A2(n_354),
.B1(n_361),
.B2(n_340),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_408),
.B1(n_391),
.B2(n_387),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_378),
.B(n_372),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_362),
.C(n_339),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_402),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_340),
.C(n_347),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_392),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_412),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_347),
.Y(n_405)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_373),
.A2(n_343),
.B1(n_339),
.B2(n_358),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_410),
.A2(n_189),
.B1(n_96),
.B2(n_138),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_393),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_378),
.B(n_172),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_414),
.B(n_415),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_369),
.B(n_360),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_360),
.Y(n_416)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_416),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_381),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_418),
.Y(n_423)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_419),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_371),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_420),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_377),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_421),
.A2(n_33),
.B1(n_124),
.B2(n_106),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_410),
.A2(n_377),
.B(n_386),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_424),
.A2(n_397),
.B(n_405),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_396),
.A2(n_375),
.B1(n_379),
.B2(n_386),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_366),
.C(n_384),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_431),
.B(n_435),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_399),
.A2(n_390),
.B1(n_383),
.B2(n_159),
.Y(n_433)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_433),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_406),
.B(n_39),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_436),
.A2(n_437),
.B1(n_444),
.B2(n_408),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_407),
.A2(n_74),
.B1(n_90),
.B2(n_33),
.Y(n_437)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_439),
.Y(n_448)
);

BUFx24_ASAP7_75t_SL g441 ( 
.A(n_404),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_441),
.Y(n_459)
);

AOI221xp5_ASAP7_75t_L g442 ( 
.A1(n_407),
.A2(n_420),
.B1(n_409),
.B2(n_402),
.C(n_417),
.Y(n_442)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_106),
.C(n_95),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_398),
.C(n_401),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_396),
.A2(n_106),
.B1(n_62),
.B2(n_54),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_414),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_449),
.Y(n_466)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_450),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_440),
.A2(n_409),
.B(n_397),
.Y(n_451)
);

OAI21x1_ASAP7_75t_SL g476 ( 
.A1(n_451),
.A2(n_458),
.B(n_9),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_452),
.B(n_460),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_400),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_454),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_411),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_462),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_423),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_412),
.C(n_413),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_416),
.C(n_40),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_461),
.B(n_463),
.Y(n_472)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_427),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_422),
.B(n_425),
.C(n_443),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_438),
.C(n_428),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_467),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_430),
.C(n_434),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_455),
.A2(n_430),
.B1(n_433),
.B2(n_423),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_470),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_445),
.A2(n_436),
.B1(n_437),
.B2(n_444),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_446),
.B(n_463),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_473),
.B(n_474),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_448),
.B(n_9),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_477),
.B(n_8),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_451),
.A2(n_8),
.B(n_14),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_447),
.C(n_453),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_472),
.C(n_465),
.Y(n_493)
);

OAI211xp5_ASAP7_75t_L g480 ( 
.A1(n_450),
.A2(n_8),
.B(n_13),
.C(n_10),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_480),
.A2(n_40),
.B(n_5),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_478),
.A2(n_449),
.B(n_464),
.Y(n_483)
);

AOI31xp67_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_486),
.A3(n_477),
.B(n_470),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_475),
.A2(n_464),
.B1(n_461),
.B2(n_459),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_488),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_485),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_469),
.A2(n_25),
.B(n_40),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_5),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_468),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_495),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_10),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_479),
.B(n_13),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_SL g503 ( 
.A(n_492),
.B(n_494),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_41),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_41),
.C(n_1),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_13),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_482),
.C(n_471),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_496),
.A2(n_499),
.B(n_0),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_497),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_489),
.A2(n_466),
.B(n_41),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_500),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_487),
.A2(n_466),
.B1(n_41),
.B2(n_5),
.Y(n_501)
);

MAJx2_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_502),
.C(n_494),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_487),
.C(n_492),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_507),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_504),
.A2(n_0),
.B(n_1),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_509),
.A2(n_511),
.B1(n_512),
.B2(n_505),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_504),
.A2(n_0),
.B(n_1),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_513),
.Y(n_517)
);

AO21x1_ASAP7_75t_SL g514 ( 
.A1(n_510),
.A2(n_503),
.B(n_1),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_515),
.C(n_0),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_508),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_515)
);

A2O1A1O1Ixp25_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_514),
.B(n_516),
.C(n_4),
.D(n_2),
.Y(n_519)
);

OA21x2_ASAP7_75t_SL g520 ( 
.A1(n_519),
.A2(n_517),
.B(n_3),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_520),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_4),
.B1(n_517),
.B2(n_510),
.Y(n_522)
);


endmodule