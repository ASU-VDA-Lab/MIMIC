module fake_jpeg_376_n_697 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_697);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_697;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_566;
wire n_374;
wire n_417;
wire n_362;
wire n_142;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_59),
.Y(n_191)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_64),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_66),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_46),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_68),
.B(n_70),
.Y(n_227)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_19),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_71),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_77),
.Y(n_197)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_18),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

CKINVDCx6p67_ASAP7_75t_R g151 ( 
.A(n_80),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_93),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_83),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g180 ( 
.A(n_87),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_89),
.Y(n_210)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_17),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_16),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_100),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_96),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_99),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_30),
.B(n_16),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_106),
.Y(n_154)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_22),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_14),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_110),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_16),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_126),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_49),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_23),
.Y(n_118)
);

INVx5_ASAP7_75t_SL g145 ( 
.A(n_118),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_15),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_35),
.B(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_15),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

BUFx2_ASAP7_75t_R g181 ( 
.A(n_131),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_141),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_68),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_146),
.A2(n_159),
.B1(n_161),
.B2(n_165),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_95),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_150),
.A2(n_171),
.B1(n_217),
.B2(n_220),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_100),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_157),
.A2(n_187),
.B1(n_214),
.B2(n_58),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_70),
.A2(n_72),
.B1(n_81),
.B2(n_79),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_112),
.A2(n_23),
.B1(n_26),
.B2(n_56),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_26),
.B1(n_54),
.B2(n_57),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_118),
.B(n_26),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_167),
.B(n_184),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_104),
.A2(n_37),
.B1(n_57),
.B2(n_35),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_178),
.B(n_4),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_67),
.B(n_35),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_193),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_114),
.A2(n_37),
.B1(n_57),
.B2(n_42),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_80),
.A2(n_33),
.B(n_21),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_189),
.A2(n_4),
.B(n_5),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_115),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_192),
.B(n_211),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_92),
.B(n_37),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_74),
.B(n_42),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_196),
.B(n_203),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_124),
.B(n_42),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_117),
.B(n_33),
.C(n_24),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_204),
.B(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_119),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_121),
.A2(n_45),
.B1(n_21),
.B2(n_47),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_87),
.A2(n_45),
.B1(n_47),
.B2(n_44),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_123),
.A2(n_45),
.B1(n_33),
.B2(n_31),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_128),
.B(n_21),
.C(n_24),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_59),
.A2(n_24),
.B1(n_25),
.B2(n_47),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_64),
.B(n_25),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_221),
.B(n_222),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_65),
.B(n_44),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_73),
.B(n_44),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_224),
.B(n_11),
.Y(n_314)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_96),
.Y(n_226)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

AO22x1_ASAP7_75t_SL g228 ( 
.A1(n_129),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_228)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_113),
.B1(n_84),
.B2(n_82),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_131),
.A2(n_31),
.B1(n_32),
.B2(n_3),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_229),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_132),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_233),
.Y(n_364)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_234),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_235),
.B(n_272),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_75),
.B1(n_32),
.B2(n_53),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_236),
.A2(n_293),
.B1(n_294),
.B2(n_273),
.Y(n_372)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_237),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_239),
.B(n_244),
.Y(n_332)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_162),
.Y(n_240)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_240),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_148),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_241),
.Y(n_358)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_152),
.Y(n_242)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_242),
.Y(n_378)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_243),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_246),
.Y(n_330)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_248),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_137),
.B1(n_175),
.B2(n_168),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_250),
.Y(n_319)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_254),
.Y(n_380)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_155),
.Y(n_255)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_257),
.Y(n_371)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_164),
.Y(n_258)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_260),
.B(n_304),
.Y(n_353)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_169),
.Y(n_262)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_L g342 ( 
.A1(n_263),
.A2(n_173),
.B1(n_180),
.B2(n_145),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_146),
.A2(n_58),
.B1(n_53),
.B2(n_41),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_273),
.B1(n_275),
.B2(n_286),
.Y(n_329)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_265),
.Y(n_352)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_163),
.Y(n_266)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_266),
.Y(n_356)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_267),
.Y(n_357)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_271),
.Y(n_360)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_278),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_216),
.A2(n_53),
.B1(n_41),
.B2(n_58),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

CKINVDCx12_ASAP7_75t_R g379 ( 
.A(n_276),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_279),
.Y(n_325)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_285),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_153),
.A2(n_58),
.B1(n_53),
.B2(n_41),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_282),
.A2(n_294),
.B1(n_141),
.B2(n_174),
.Y(n_322)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_136),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_296),
.Y(n_346)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_186),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_284),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_159),
.B(n_13),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_287),
.B(n_300),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_176),
.A2(n_58),
.B1(n_53),
.B2(n_41),
.Y(n_288)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_290),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_226),
.A2(n_58),
.B1(n_53),
.B2(n_41),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_149),
.A2(n_41),
.B1(n_12),
.B2(n_6),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_228),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_150),
.A2(n_12),
.B1(n_5),
.B2(n_7),
.Y(n_294)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_163),
.Y(n_296)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_301),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_8),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_143),
.B(n_12),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_139),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_305),
.Y(n_345)
);

BUFx12_ASAP7_75t_L g303 ( 
.A(n_182),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_303),
.Y(n_323)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_138),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_149),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_307),
.Y(n_375)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_199),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_217),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_308),
.A2(n_316),
.B1(n_317),
.B2(n_173),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_229),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_309),
.A2(n_154),
.B1(n_218),
.B2(n_215),
.Y(n_355)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_139),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_313),
.Y(n_376)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_311),
.B(n_314),
.Y(n_381)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_199),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_133),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_315),
.Y(n_367)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_133),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_181),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_174),
.B(n_7),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_181),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_322),
.A2(n_372),
.B1(n_266),
.B2(n_298),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_331),
.B(n_350),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_333),
.B(n_9),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_250),
.B(n_205),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_366),
.C(n_288),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_180),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_349),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_295),
.B(n_145),
.CI(n_180),
.CON(n_347),
.SN(n_347)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_282),
.C(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_190),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_312),
.B(n_190),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_317),
.A2(n_143),
.B1(n_154),
.B2(n_148),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_289),
.B(n_215),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_362),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_236),
.B1(n_277),
.B2(n_321),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_263),
.A2(n_218),
.B(n_186),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_361),
.A2(n_291),
.B(n_292),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_252),
.B(n_140),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_295),
.B(n_197),
.C(n_188),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_264),
.A2(n_197),
.B1(n_188),
.B2(n_210),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_269),
.A2(n_210),
.B1(n_170),
.B2(n_225),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_373),
.A2(n_276),
.B1(n_241),
.B2(n_275),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_297),
.B(n_295),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_235),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_377),
.A2(n_269),
.B1(n_247),
.B2(n_309),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_393),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_383),
.A2(n_405),
.B1(n_416),
.B2(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_387),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_395),
.Y(n_450)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_270),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_394),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_235),
.Y(n_394)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_293),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_409),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_238),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_403),
.C(n_411),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_310),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_251),
.C(n_249),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_329),
.A2(n_209),
.B1(n_158),
.B2(n_147),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_404),
.A2(n_407),
.B1(n_339),
.B2(n_357),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_329),
.A2(n_253),
.B1(n_267),
.B2(n_290),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_334),
.Y(n_406)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_333),
.B(n_301),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_303),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_356),
.Y(n_412)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_412),
.Y(n_471)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_332),
.B(n_302),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_420),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_321),
.A2(n_144),
.B1(n_209),
.B2(n_134),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_321),
.A2(n_144),
.B1(n_158),
.B2(n_134),
.Y(n_417)
);

AOI22x1_ASAP7_75t_L g418 ( 
.A1(n_347),
.A2(n_279),
.B1(n_276),
.B2(n_303),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_419),
.Y(n_447)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_353),
.B(n_296),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_319),
.B(n_311),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_423),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_319),
.B(n_331),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_346),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_426),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_261),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_363),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_427),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_338),
.B(n_284),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_428),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_322),
.B(n_256),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_431),
.C(n_361),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_340),
.A2(n_261),
.B1(n_233),
.B2(n_156),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_430),
.A2(n_325),
.B(n_358),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_323),
.B(n_142),
.C(n_156),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_432),
.Y(n_434)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_442),
.B(n_367),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_390),
.A2(n_347),
.B1(n_342),
.B2(n_339),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_444),
.A2(n_455),
.B1(n_459),
.B2(n_408),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_382),
.A2(n_327),
.B1(n_323),
.B2(n_368),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_445),
.A2(n_451),
.B1(n_413),
.B2(n_396),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_394),
.A2(n_407),
.B1(n_398),
.B2(n_388),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_446),
.A2(n_457),
.B1(n_470),
.B2(n_401),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_352),
.C(n_359),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_449),
.B(n_475),
.C(n_360),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_429),
.A2(n_388),
.B1(n_418),
.B2(n_392),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_397),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_464),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_404),
.A2(n_363),
.B1(n_345),
.B2(n_376),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_425),
.A2(n_147),
.B1(n_140),
.B2(n_363),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_424),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_395),
.A2(n_368),
.B1(n_375),
.B2(n_346),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_393),
.A2(n_346),
.B(n_380),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_423),
.A2(n_365),
.B(n_367),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_465),
.A2(n_427),
.B(n_385),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_387),
.A2(n_368),
.B1(n_142),
.B2(n_364),
.Y(n_470)
);

AOI32xp33_ASAP7_75t_L g473 ( 
.A1(n_386),
.A2(n_409),
.A3(n_418),
.B1(n_408),
.B2(n_421),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_386),
.B(n_359),
.Y(n_475)
);

MAJx2_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_411),
.C(n_384),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_477),
.B(n_486),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_403),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_478),
.B(n_492),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_479),
.B(n_490),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_480),
.A2(n_488),
.B1(n_489),
.B2(n_499),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_431),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_481),
.B(n_509),
.C(n_442),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_483),
.A2(n_441),
.B1(n_447),
.B2(n_465),
.Y(n_524)
);

HAxp5_ASAP7_75t_SL g484 ( 
.A(n_443),
.B(n_430),
.CON(n_484),
.SN(n_484)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_487),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_446),
.A2(n_401),
.B1(n_421),
.B2(n_414),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_456),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_406),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_491),
.B(n_510),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_460),
.B(n_410),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_456),
.Y(n_494)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_494),
.Y(n_528)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_472),
.Y(n_495)
);

INVx3_ASAP7_75t_SL g531 ( 
.A(n_495),
.Y(n_531)
);

AOI322xp5_ASAP7_75t_L g496 ( 
.A1(n_461),
.A2(n_427),
.A3(n_402),
.B1(n_391),
.B2(n_419),
.C1(n_432),
.C2(n_414),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_496),
.B(n_503),
.Y(n_519)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_435),
.Y(n_497)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_379),
.C(n_397),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_514),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_451),
.A2(n_432),
.B1(n_364),
.B2(n_412),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_500),
.A2(n_502),
.B1(n_515),
.B2(n_494),
.Y(n_547)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_501),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_470),
.A2(n_426),
.B1(n_352),
.B2(n_360),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_436),
.B(n_380),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_326),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_505),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_462),
.B(n_326),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_462),
.B(n_326),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_506),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_443),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_341),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_508),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_433),
.B(n_458),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_460),
.B(n_341),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_511),
.Y(n_544)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_512),
.Y(n_521)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_439),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_436),
.B(n_371),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_371),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_482),
.A2(n_441),
.B1(n_444),
.B2(n_447),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_520),
.A2(n_533),
.B1(n_542),
.B2(n_546),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_523),
.B(n_543),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_524),
.A2(n_525),
.B1(n_536),
.B2(n_541),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_499),
.A2(n_441),
.B1(n_445),
.B2(n_447),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_526),
.B(n_545),
.C(n_549),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_477),
.B(n_459),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_532),
.B(n_530),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_482),
.A2(n_467),
.B1(n_438),
.B2(n_473),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_483),
.A2(n_464),
.B1(n_454),
.B2(n_463),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_493),
.A2(n_464),
.B1(n_457),
.B2(n_455),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_493),
.A2(n_464),
.B1(n_448),
.B2(n_466),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_466),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_481),
.B(n_448),
.C(n_439),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_480),
.A2(n_476),
.B1(n_485),
.B2(n_488),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_547),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_476),
.A2(n_452),
.B(n_453),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_548),
.A2(n_513),
.B(n_512),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_452),
.C(n_469),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_485),
.A2(n_434),
.B1(n_469),
.B2(n_474),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_550),
.A2(n_474),
.B1(n_472),
.B2(n_348),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_369),
.C(n_348),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_497),
.C(n_487),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_507),
.B(n_486),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_554),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_508),
.B(n_378),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_504),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_555),
.B(n_562),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_SL g597 ( 
.A(n_556),
.B(n_559),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_544),
.B(n_511),
.Y(n_557)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_557),
.Y(n_594)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_521),
.Y(n_558)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_558),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_530),
.B(n_532),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_521),
.Y(n_560)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_489),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_517),
.B(n_490),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_564),
.B(n_571),
.Y(n_599)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_565),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_533),
.A2(n_479),
.B1(n_500),
.B2(n_506),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_566),
.A2(n_578),
.B1(n_525),
.B2(n_550),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_568),
.A2(n_534),
.B(n_528),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_505),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_582),
.Y(n_589)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_570),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_501),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_552),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_580),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_575),
.C(n_586),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_523),
.B(n_471),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_574),
.B(n_577),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_526),
.B(n_502),
.C(n_471),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_527),
.A2(n_495),
.B(n_434),
.Y(n_577)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_531),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_579),
.Y(n_605)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_581),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_SL g582 ( 
.A(n_545),
.B(n_379),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_587),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_553),
.B(n_474),
.C(n_378),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_535),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_588),
.A2(n_590),
.B1(n_585),
.B2(n_561),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_563),
.A2(n_541),
.B1(n_536),
.B2(n_524),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_549),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_595),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_567),
.B(n_542),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_546),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_576),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_568),
.B(n_539),
.Y(n_598)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_598),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_563),
.A2(n_534),
.B(n_548),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_601),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_575),
.B(n_528),
.C(n_554),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_603),
.B(n_606),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_584),
.B(n_576),
.C(n_586),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_585),
.A2(n_538),
.B1(n_520),
.B2(n_529),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_607),
.A2(n_578),
.B1(n_531),
.B2(n_556),
.Y(n_626)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_608),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_584),
.B(n_519),
.C(n_540),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_611),
.B(n_562),
.C(n_569),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_615),
.A2(n_609),
.B1(n_604),
.B2(n_600),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_595),
.B(n_555),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_618),
.B(n_619),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_620),
.B(n_627),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_591),
.B(n_566),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_622),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_612),
.Y(n_622)
);

AO22x1_ASAP7_75t_L g623 ( 
.A1(n_590),
.A2(n_587),
.B1(n_580),
.B2(n_551),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_623),
.B(n_608),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_572),
.C(n_573),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_624),
.B(n_625),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_599),
.A2(n_535),
.B1(n_551),
.B2(n_539),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_626),
.B(n_630),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_596),
.B(n_559),
.C(n_472),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_369),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_606),
.B(n_603),
.C(n_611),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_631),
.B(n_633),
.C(n_605),
.Y(n_639)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_602),
.Y(n_632)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_632),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_592),
.B(n_328),
.C(n_330),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_634),
.Y(n_644)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_610),
.Y(n_636)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_636),
.Y(n_654)
);

FAx1_ASAP7_75t_L g638 ( 
.A(n_629),
.B(n_628),
.CI(n_601),
.CON(n_638),
.SN(n_638)
);

AOI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_638),
.A2(n_645),
.B(n_644),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_639),
.B(n_646),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_645),
.A2(n_627),
.B1(n_617),
.B2(n_619),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_624),
.B(n_607),
.C(n_588),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_616),
.A2(n_598),
.B(n_614),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_647),
.A2(n_655),
.B(n_328),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_622),
.B(n_594),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_648),
.B(n_649),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_635),
.B(n_589),
.C(n_597),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_650),
.B(n_651),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_631),
.B(n_589),
.C(n_597),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_620),
.B(n_613),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_652),
.B(n_618),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_621),
.B(n_609),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_656),
.B(n_640),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_657),
.A2(n_665),
.B(n_649),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_638),
.A2(n_623),
.B1(n_600),
.B2(n_604),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_658),
.A2(n_642),
.B1(n_641),
.B2(n_651),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_633),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_659),
.B(n_660),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_637),
.B(n_630),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_661),
.A2(n_650),
.B1(n_374),
.B2(n_337),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_617),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_662),
.B(n_663),
.Y(n_673)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_654),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_640),
.B(n_365),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_664),
.B(n_667),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_653),
.B(n_330),
.C(n_374),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_647),
.A2(n_655),
.B(n_638),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_670),
.B(n_646),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_672),
.B(n_675),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_676),
.A2(n_680),
.B(n_657),
.Y(n_681)
);

BUFx24_ASAP7_75t_SL g677 ( 
.A(n_668),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_677),
.B(n_660),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_678),
.B(n_679),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_666),
.B(n_641),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_681),
.B(n_682),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_671),
.A2(n_669),
.B(n_658),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_683),
.B(n_337),
.C(n_177),
.Y(n_690)
);

OAI321xp33_ASAP7_75t_L g686 ( 
.A1(n_673),
.A2(n_672),
.A3(n_663),
.B1(n_674),
.B2(n_680),
.C(n_667),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_686),
.B(n_687),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_679),
.B(n_661),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_685),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_689),
.A2(n_690),
.B(n_684),
.Y(n_692)
);

OAI21x1_ASAP7_75t_SL g694 ( 
.A1(n_692),
.A2(n_693),
.B(n_688),
.Y(n_694)
);

AOI321xp33_ASAP7_75t_L g693 ( 
.A1(n_691),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_677),
.C(n_682),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_694),
.B(n_9),
.C(n_10),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_695),
.B(n_9),
.Y(n_696)
);

XNOR2xp5_ASAP7_75t_L g697 ( 
.A(n_696),
.B(n_10),
.Y(n_697)
);


endmodule